
module fpregfile ( rs, rd, rData, wData, regWr, clk, fp );
  input [4:0] rs;
  input [4:0] rd;
  output [31:0] rData;
  input [31:0] wData;
  input regWr, clk, fp;
  wire   N9, N10, N11, N12, N13, \mem[31][31] , \mem[31][30] , \mem[31][29] ,
         \mem[31][28] , \mem[31][27] , \mem[31][26] , \mem[31][25] ,
         \mem[31][24] , \mem[31][23] , \mem[31][22] , \mem[31][21] ,
         \mem[31][20] , \mem[31][19] , \mem[31][18] , \mem[31][17] ,
         \mem[31][16] , \mem[31][15] , \mem[31][14] , \mem[31][13] ,
         \mem[31][12] , \mem[31][11] , \mem[31][10] , \mem[31][9] ,
         \mem[31][8] , \mem[31][7] , \mem[31][6] , \mem[31][5] , \mem[31][4] ,
         \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] , \mem[30][31] ,
         \mem[30][30] , \mem[30][29] , \mem[30][28] , \mem[30][27] ,
         \mem[30][26] , \mem[30][25] , \mem[30][24] , \mem[30][23] ,
         \mem[30][22] , \mem[30][21] , \mem[30][20] , \mem[30][19] ,
         \mem[30][18] , \mem[30][17] , \mem[30][16] , \mem[30][15] ,
         \mem[30][14] , \mem[30][13] , \mem[30][12] , \mem[30][11] ,
         \mem[30][10] , \mem[30][9] , \mem[30][8] , \mem[30][7] , \mem[30][6] ,
         \mem[30][5] , \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] ,
         \mem[30][0] , \mem[29][31] , \mem[29][30] , \mem[29][29] ,
         \mem[29][28] , \mem[29][27] , \mem[29][26] , \mem[29][25] ,
         \mem[29][24] , \mem[29][23] , \mem[29][22] , \mem[29][21] ,
         \mem[29][20] , \mem[29][19] , \mem[29][18] , \mem[29][17] ,
         \mem[29][16] , \mem[29][15] , \mem[29][14] , \mem[29][13] ,
         \mem[29][12] , \mem[29][11] , \mem[29][10] , \mem[29][9] ,
         \mem[29][8] , \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] ,
         \mem[29][3] , \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[28][31] ,
         \mem[28][30] , \mem[28][29] , \mem[28][28] , \mem[28][27] ,
         \mem[28][26] , \mem[28][25] , \mem[28][24] , \mem[28][23] ,
         \mem[28][22] , \mem[28][21] , \mem[28][20] , \mem[28][19] ,
         \mem[28][18] , \mem[28][17] , \mem[28][16] , \mem[28][15] ,
         \mem[28][14] , \mem[28][13] , \mem[28][12] , \mem[28][11] ,
         \mem[28][10] , \mem[28][9] , \mem[28][8] , \mem[28][7] , \mem[28][6] ,
         \mem[28][5] , \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] ,
         \mem[28][0] , \mem[27][31] , \mem[27][30] , \mem[27][29] ,
         \mem[27][28] , \mem[27][27] , \mem[27][26] , \mem[27][25] ,
         \mem[27][24] , \mem[27][23] , \mem[27][22] , \mem[27][21] ,
         \mem[27][20] , \mem[27][19] , \mem[27][18] , \mem[27][17] ,
         \mem[27][16] , \mem[27][15] , \mem[27][14] , \mem[27][13] ,
         \mem[27][12] , \mem[27][11] , \mem[27][10] , \mem[27][9] ,
         \mem[27][8] , \mem[27][7] , \mem[27][6] , \mem[27][5] , \mem[27][4] ,
         \mem[27][3] , \mem[27][2] , \mem[27][1] , \mem[27][0] , \mem[26][31] ,
         \mem[26][30] , \mem[26][29] , \mem[26][28] , \mem[26][27] ,
         \mem[26][26] , \mem[26][25] , \mem[26][24] , \mem[26][23] ,
         \mem[26][22] , \mem[26][21] , \mem[26][20] , \mem[26][19] ,
         \mem[26][18] , \mem[26][17] , \mem[26][16] , \mem[26][15] ,
         \mem[26][14] , \mem[26][13] , \mem[26][12] , \mem[26][11] ,
         \mem[26][10] , \mem[26][9] , \mem[26][8] , \mem[26][7] , \mem[26][6] ,
         \mem[26][5] , \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] ,
         \mem[26][0] , \mem[25][31] , \mem[25][30] , \mem[25][29] ,
         \mem[25][28] , \mem[25][27] , \mem[25][26] , \mem[25][25] ,
         \mem[25][24] , \mem[25][23] , \mem[25][22] , \mem[25][21] ,
         \mem[25][20] , \mem[25][19] , \mem[25][18] , \mem[25][17] ,
         \mem[25][16] , \mem[25][15] , \mem[25][14] , \mem[25][13] ,
         \mem[25][12] , \mem[25][11] , \mem[25][10] , \mem[25][9] ,
         \mem[25][8] , \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] ,
         \mem[25][3] , \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][31] ,
         \mem[24][30] , \mem[24][29] , \mem[24][28] , \mem[24][27] ,
         \mem[24][26] , \mem[24][25] , \mem[24][24] , \mem[24][23] ,
         \mem[24][22] , \mem[24][21] , \mem[24][20] , \mem[24][19] ,
         \mem[24][18] , \mem[24][17] , \mem[24][16] , \mem[24][15] ,
         \mem[24][14] , \mem[24][13] , \mem[24][12] , \mem[24][11] ,
         \mem[24][10] , \mem[24][9] , \mem[24][8] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][31] , \mem[23][30] , \mem[23][29] ,
         \mem[23][28] , \mem[23][27] , \mem[23][26] , \mem[23][25] ,
         \mem[23][24] , \mem[23][23] , \mem[23][22] , \mem[23][21] ,
         \mem[23][20] , \mem[23][19] , \mem[23][18] , \mem[23][17] ,
         \mem[23][16] , \mem[23][15] , \mem[23][14] , \mem[23][13] ,
         \mem[23][12] , \mem[23][11] , \mem[23][10] , \mem[23][9] ,
         \mem[23][8] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][31] ,
         \mem[22][30] , \mem[22][29] , \mem[22][28] , \mem[22][27] ,
         \mem[22][26] , \mem[22][25] , \mem[22][24] , \mem[22][23] ,
         \mem[22][22] , \mem[22][21] , \mem[22][20] , \mem[22][19] ,
         \mem[22][18] , \mem[22][17] , \mem[22][16] , \mem[22][15] ,
         \mem[22][14] , \mem[22][13] , \mem[22][12] , \mem[22][11] ,
         \mem[22][10] , \mem[22][9] , \mem[22][8] , \mem[22][7] , \mem[22][6] ,
         \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] , \mem[22][1] ,
         \mem[22][0] , \mem[21][31] , \mem[21][30] , \mem[21][29] ,
         \mem[21][28] , \mem[21][27] , \mem[21][26] , \mem[21][25] ,
         \mem[21][24] , \mem[21][23] , \mem[21][22] , \mem[21][21] ,
         \mem[21][20] , \mem[21][19] , \mem[21][18] , \mem[21][17] ,
         \mem[21][16] , \mem[21][15] , \mem[21][14] , \mem[21][13] ,
         \mem[21][12] , \mem[21][11] , \mem[21][10] , \mem[21][9] ,
         \mem[21][8] , \mem[21][7] , \mem[21][6] , \mem[21][5] , \mem[21][4] ,
         \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] , \mem[20][31] ,
         \mem[20][30] , \mem[20][29] , \mem[20][28] , \mem[20][27] ,
         \mem[20][26] , \mem[20][25] , \mem[20][24] , \mem[20][23] ,
         \mem[20][22] , \mem[20][21] , \mem[20][20] , \mem[20][19] ,
         \mem[20][18] , \mem[20][17] , \mem[20][16] , \mem[20][15] ,
         \mem[20][14] , \mem[20][13] , \mem[20][12] , \mem[20][11] ,
         \mem[20][10] , \mem[20][9] , \mem[20][8] , \mem[20][7] , \mem[20][6] ,
         \mem[20][5] , \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] ,
         \mem[20][0] , \mem[19][31] , \mem[19][30] , \mem[19][29] ,
         \mem[19][28] , \mem[19][27] , \mem[19][26] , \mem[19][25] ,
         \mem[19][24] , \mem[19][23] , \mem[19][22] , \mem[19][21] ,
         \mem[19][20] , \mem[19][19] , \mem[19][18] , \mem[19][17] ,
         \mem[19][16] , \mem[19][15] , \mem[19][14] , \mem[19][13] ,
         \mem[19][12] , \mem[19][11] , \mem[19][10] , \mem[19][9] ,
         \mem[19][8] , \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] ,
         \mem[19][3] , \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[18][31] ,
         \mem[18][30] , \mem[18][29] , \mem[18][28] , \mem[18][27] ,
         \mem[18][26] , \mem[18][25] , \mem[18][24] , \mem[18][23] ,
         \mem[18][22] , \mem[18][21] , \mem[18][20] , \mem[18][19] ,
         \mem[18][18] , \mem[18][17] , \mem[18][16] , \mem[18][15] ,
         \mem[18][14] , \mem[18][13] , \mem[18][12] , \mem[18][11] ,
         \mem[18][10] , \mem[18][9] , \mem[18][8] , \mem[18][7] , \mem[18][6] ,
         \mem[18][5] , \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] ,
         \mem[18][0] , \mem[17][31] , \mem[17][30] , \mem[17][29] ,
         \mem[17][28] , \mem[17][27] , \mem[17][26] , \mem[17][25] ,
         \mem[17][24] , \mem[17][23] , \mem[17][22] , \mem[17][21] ,
         \mem[17][20] , \mem[17][19] , \mem[17][18] , \mem[17][17] ,
         \mem[17][16] , \mem[17][15] , \mem[17][14] , \mem[17][13] ,
         \mem[17][12] , \mem[17][11] , \mem[17][10] , \mem[17][9] ,
         \mem[17][8] , \mem[17][7] , \mem[17][6] , \mem[17][5] , \mem[17][4] ,
         \mem[17][3] , \mem[17][2] , \mem[17][1] , \mem[17][0] , \mem[16][31] ,
         \mem[16][30] , \mem[16][29] , \mem[16][28] , \mem[16][27] ,
         \mem[16][26] , \mem[16][25] , \mem[16][24] , \mem[16][23] ,
         \mem[16][22] , \mem[16][21] , \mem[16][20] , \mem[16][19] ,
         \mem[16][18] , \mem[16][17] , \mem[16][16] , \mem[16][15] ,
         \mem[16][14] , \mem[16][13] , \mem[16][12] , \mem[16][11] ,
         \mem[16][10] , \mem[16][9] , \mem[16][8] , \mem[16][7] , \mem[16][6] ,
         \mem[16][5] , \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] ,
         \mem[16][0] , \mem[15][31] , \mem[15][30] , \mem[15][29] ,
         \mem[15][28] , \mem[15][27] , \mem[15][26] , \mem[15][25] ,
         \mem[15][24] , \mem[15][23] , \mem[15][22] , \mem[15][21] ,
         \mem[15][20] , \mem[15][19] , \mem[15][18] , \mem[15][17] ,
         \mem[15][16] , \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][31] ,
         \mem[14][30] , \mem[14][29] , \mem[14][28] , \mem[14][27] ,
         \mem[14][26] , \mem[14][25] , \mem[14][24] , \mem[14][23] ,
         \mem[14][22] , \mem[14][21] , \mem[14][20] , \mem[14][19] ,
         \mem[14][18] , \mem[14][17] , \mem[14][16] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][31] , \mem[13][30] , \mem[13][29] ,
         \mem[13][28] , \mem[13][27] , \mem[13][26] , \mem[13][25] ,
         \mem[13][24] , \mem[13][23] , \mem[13][22] , \mem[13][21] ,
         \mem[13][20] , \mem[13][19] , \mem[13][18] , \mem[13][17] ,
         \mem[13][16] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][31] ,
         \mem[12][30] , \mem[12][29] , \mem[12][28] , \mem[12][27] ,
         \mem[12][26] , \mem[12][25] , \mem[12][24] , \mem[12][23] ,
         \mem[12][22] , \mem[12][21] , \mem[12][20] , \mem[12][19] ,
         \mem[12][18] , \mem[12][17] , \mem[12][16] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][31] , \mem[11][30] , \mem[11][29] ,
         \mem[11][28] , \mem[11][27] , \mem[11][26] , \mem[11][25] ,
         \mem[11][24] , \mem[11][23] , \mem[11][22] , \mem[11][21] ,
         \mem[11][20] , \mem[11][19] , \mem[11][18] , \mem[11][17] ,
         \mem[11][16] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][31] ,
         \mem[10][30] , \mem[10][29] , \mem[10][28] , \mem[10][27] ,
         \mem[10][26] , \mem[10][25] , \mem[10][24] , \mem[10][23] ,
         \mem[10][22] , \mem[10][21] , \mem[10][20] , \mem[10][19] ,
         \mem[10][18] , \mem[10][17] , \mem[10][16] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][31] , \mem[9][30] , \mem[9][29] , \mem[9][28] ,
         \mem[9][27] , \mem[9][26] , \mem[9][25] , \mem[9][24] , \mem[9][23] ,
         \mem[9][22] , \mem[9][21] , \mem[9][20] , \mem[9][19] , \mem[9][18] ,
         \mem[9][17] , \mem[9][16] , \mem[9][15] , \mem[9][14] , \mem[9][13] ,
         \mem[9][12] , \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][31] , \mem[8][30] ,
         \mem[8][29] , \mem[8][28] , \mem[8][27] , \mem[8][26] , \mem[8][25] ,
         \mem[8][24] , \mem[8][23] , \mem[8][22] , \mem[8][21] , \mem[8][20] ,
         \mem[8][19] , \mem[8][18] , \mem[8][17] , \mem[8][16] , \mem[8][15] ,
         \mem[8][14] , \mem[8][13] , \mem[8][12] , \mem[8][11] , \mem[8][10] ,
         \mem[8][9] , \mem[8][8] , \mem[8][7] , \mem[8][6] , \mem[8][5] ,
         \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] ,
         \mem[7][31] , \mem[7][30] , \mem[7][29] , \mem[7][28] , \mem[7][27] ,
         \mem[7][26] , \mem[7][25] , \mem[7][24] , \mem[7][23] , \mem[7][22] ,
         \mem[7][21] , \mem[7][20] , \mem[7][19] , \mem[7][18] , \mem[7][17] ,
         \mem[7][16] , \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][31] , \mem[6][30] , \mem[6][29] ,
         \mem[6][28] , \mem[6][27] , \mem[6][26] , \mem[6][25] , \mem[6][24] ,
         \mem[6][23] , \mem[6][22] , \mem[6][21] , \mem[6][20] , \mem[6][19] ,
         \mem[6][18] , \mem[6][17] , \mem[6][16] , \mem[6][15] , \mem[6][14] ,
         \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] ,
         \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] ,
         \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][31] ,
         \mem[5][30] , \mem[5][29] , \mem[5][28] , \mem[5][27] , \mem[5][26] ,
         \mem[5][25] , \mem[5][24] , \mem[5][23] , \mem[5][22] , \mem[5][21] ,
         \mem[5][20] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][31] , \mem[4][30] , \mem[4][29] , \mem[4][28] ,
         \mem[4][27] , \mem[4][26] , \mem[4][25] , \mem[4][24] , \mem[4][23] ,
         \mem[4][22] , \mem[4][21] , \mem[4][20] , \mem[4][19] , \mem[4][18] ,
         \mem[4][17] , \mem[4][16] , \mem[4][15] , \mem[4][14] , \mem[4][13] ,
         \mem[4][12] , \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][31] , \mem[3][30] ,
         \mem[3][29] , \mem[3][28] , \mem[3][27] , \mem[3][26] , \mem[3][25] ,
         \mem[3][24] , \mem[3][23] , \mem[3][22] , \mem[3][21] , \mem[3][20] ,
         \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] , \mem[3][15] ,
         \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] , \mem[3][10] ,
         \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[2][31] , \mem[2][30] , \mem[2][29] , \mem[2][28] , \mem[2][27] ,
         \mem[2][26] , \mem[2][25] , \mem[2][24] , \mem[2][23] , \mem[2][22] ,
         \mem[2][21] , \mem[2][20] , \mem[2][19] , \mem[2][18] , \mem[2][17] ,
         \mem[2][16] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][31] , \mem[1][30] , \mem[1][29] ,
         \mem[1][28] , \mem[1][27] , \mem[1][26] , \mem[1][25] , \mem[1][24] ,
         \mem[1][23] , \mem[1][22] , \mem[1][21] , \mem[1][20] , \mem[1][19] ,
         \mem[1][18] , \mem[1][17] , \mem[1][16] , \mem[1][15] , \mem[1][14] ,
         \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] ,
         \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][31] ,
         \mem[0][30] , \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] ,
         \mem[0][25] , \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] ,
         \mem[0][20] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23,
         n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51,
         n53, n55, n57, n59, n61, n63, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n4406, n4407, n4408, n4409, n4410;
  assign N9 = rs[0];
  assign N10 = rs[1];
  assign N11 = rs[2];
  assign N12 = rs[3];
  assign N13 = rs[4];

  DFF_X2 \mem_reg[31][31]  ( .D(n2136), .CK(clk), .Q(\mem[31][31] ) );
  DFF_X2 \mem_reg[31][30]  ( .D(n2135), .CK(clk), .Q(\mem[31][30] ) );
  DFF_X2 \mem_reg[31][29]  ( .D(n2134), .CK(clk), .Q(\mem[31][29] ) );
  DFF_X2 \mem_reg[31][28]  ( .D(n2133), .CK(clk), .Q(\mem[31][28] ) );
  DFF_X2 \mem_reg[31][27]  ( .D(n2132), .CK(clk), .Q(\mem[31][27] ) );
  DFF_X2 \mem_reg[31][26]  ( .D(n2131), .CK(clk), .Q(\mem[31][26] ) );
  DFF_X2 \mem_reg[31][25]  ( .D(n2130), .CK(clk), .Q(\mem[31][25] ) );
  DFF_X2 \mem_reg[31][24]  ( .D(n2129), .CK(clk), .Q(\mem[31][24] ) );
  DFF_X2 \mem_reg[31][23]  ( .D(n2128), .CK(clk), .Q(\mem[31][23] ) );
  DFF_X2 \mem_reg[31][22]  ( .D(n2127), .CK(clk), .Q(\mem[31][22] ) );
  DFF_X2 \mem_reg[31][21]  ( .D(n2126), .CK(clk), .Q(\mem[31][21] ) );
  DFF_X2 \mem_reg[31][20]  ( .D(n2125), .CK(clk), .Q(\mem[31][20] ) );
  DFF_X2 \mem_reg[31][19]  ( .D(n2124), .CK(clk), .Q(\mem[31][19] ) );
  DFF_X2 \mem_reg[31][18]  ( .D(n2123), .CK(clk), .Q(\mem[31][18] ) );
  DFF_X2 \mem_reg[31][17]  ( .D(n2122), .CK(clk), .Q(\mem[31][17] ) );
  DFF_X2 \mem_reg[31][16]  ( .D(n2121), .CK(clk), .Q(\mem[31][16] ) );
  DFF_X2 \mem_reg[31][15]  ( .D(n2120), .CK(clk), .Q(\mem[31][15] ) );
  DFF_X2 \mem_reg[31][14]  ( .D(n2119), .CK(clk), .Q(\mem[31][14] ) );
  DFF_X2 \mem_reg[31][13]  ( .D(n2118), .CK(clk), .Q(\mem[31][13] ) );
  DFF_X2 \mem_reg[31][12]  ( .D(n2117), .CK(clk), .Q(\mem[31][12] ) );
  DFF_X2 \mem_reg[31][11]  ( .D(n2116), .CK(clk), .Q(\mem[31][11] ) );
  DFF_X2 \mem_reg[31][10]  ( .D(n2115), .CK(clk), .Q(\mem[31][10] ) );
  DFF_X2 \mem_reg[31][9]  ( .D(n2114), .CK(clk), .Q(\mem[31][9] ) );
  DFF_X2 \mem_reg[31][8]  ( .D(n2113), .CK(clk), .Q(\mem[31][8] ) );
  DFF_X2 \mem_reg[31][7]  ( .D(n2112), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X2 \mem_reg[31][6]  ( .D(n2111), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X2 \mem_reg[31][5]  ( .D(n2110), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X2 \mem_reg[31][4]  ( .D(n2109), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X2 \mem_reg[31][3]  ( .D(n2108), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X2 \mem_reg[31][2]  ( .D(n2107), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X2 \mem_reg[31][1]  ( .D(n2106), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X2 \mem_reg[31][0]  ( .D(n2105), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X2 \mem_reg[30][31]  ( .D(n2104), .CK(clk), .Q(\mem[30][31] ) );
  DFF_X2 \mem_reg[30][30]  ( .D(n2103), .CK(clk), .Q(\mem[30][30] ) );
  DFF_X2 \mem_reg[30][29]  ( .D(n2102), .CK(clk), .Q(\mem[30][29] ) );
  DFF_X2 \mem_reg[30][28]  ( .D(n2101), .CK(clk), .Q(\mem[30][28] ) );
  DFF_X2 \mem_reg[30][27]  ( .D(n2100), .CK(clk), .Q(\mem[30][27] ) );
  DFF_X2 \mem_reg[30][26]  ( .D(n2099), .CK(clk), .Q(\mem[30][26] ) );
  DFF_X2 \mem_reg[30][25]  ( .D(n2098), .CK(clk), .Q(\mem[30][25] ) );
  DFF_X2 \mem_reg[30][24]  ( .D(n2097), .CK(clk), .Q(\mem[30][24] ) );
  DFF_X2 \mem_reg[30][23]  ( .D(n2096), .CK(clk), .Q(\mem[30][23] ) );
  DFF_X2 \mem_reg[30][22]  ( .D(n2095), .CK(clk), .Q(\mem[30][22] ) );
  DFF_X2 \mem_reg[30][21]  ( .D(n2094), .CK(clk), .Q(\mem[30][21] ) );
  DFF_X2 \mem_reg[30][20]  ( .D(n2093), .CK(clk), .Q(\mem[30][20] ) );
  DFF_X2 \mem_reg[30][19]  ( .D(n2092), .CK(clk), .Q(\mem[30][19] ) );
  DFF_X2 \mem_reg[30][18]  ( .D(n2091), .CK(clk), .Q(\mem[30][18] ) );
  DFF_X2 \mem_reg[30][17]  ( .D(n2090), .CK(clk), .Q(\mem[30][17] ) );
  DFF_X2 \mem_reg[30][16]  ( .D(n2089), .CK(clk), .Q(\mem[30][16] ) );
  DFF_X2 \mem_reg[30][15]  ( .D(n2088), .CK(clk), .Q(\mem[30][15] ) );
  DFF_X2 \mem_reg[30][14]  ( .D(n2087), .CK(clk), .Q(\mem[30][14] ) );
  DFF_X2 \mem_reg[30][13]  ( .D(n2086), .CK(clk), .Q(\mem[30][13] ) );
  DFF_X2 \mem_reg[30][12]  ( .D(n2085), .CK(clk), .Q(\mem[30][12] ) );
  DFF_X2 \mem_reg[30][11]  ( .D(n2084), .CK(clk), .Q(\mem[30][11] ) );
  DFF_X2 \mem_reg[30][10]  ( .D(n2083), .CK(clk), .Q(\mem[30][10] ) );
  DFF_X2 \mem_reg[30][9]  ( .D(n2082), .CK(clk), .Q(\mem[30][9] ) );
  DFF_X2 \mem_reg[30][8]  ( .D(n2081), .CK(clk), .Q(\mem[30][8] ) );
  DFF_X2 \mem_reg[30][7]  ( .D(n2080), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X2 \mem_reg[30][6]  ( .D(n2079), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X2 \mem_reg[30][5]  ( .D(n2078), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X2 \mem_reg[30][4]  ( .D(n2077), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X2 \mem_reg[30][3]  ( .D(n2076), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X2 \mem_reg[30][2]  ( .D(n2075), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X2 \mem_reg[30][1]  ( .D(n2074), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X2 \mem_reg[30][0]  ( .D(n2073), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X2 \mem_reg[29][31]  ( .D(n2072), .CK(clk), .Q(\mem[29][31] ) );
  DFF_X2 \mem_reg[29][30]  ( .D(n2071), .CK(clk), .Q(\mem[29][30] ) );
  DFF_X2 \mem_reg[29][29]  ( .D(n2070), .CK(clk), .Q(\mem[29][29] ) );
  DFF_X2 \mem_reg[29][28]  ( .D(n2069), .CK(clk), .Q(\mem[29][28] ) );
  DFF_X2 \mem_reg[29][27]  ( .D(n2068), .CK(clk), .Q(\mem[29][27] ) );
  DFF_X2 \mem_reg[29][26]  ( .D(n2067), .CK(clk), .Q(\mem[29][26] ) );
  DFF_X2 \mem_reg[29][25]  ( .D(n2066), .CK(clk), .Q(\mem[29][25] ) );
  DFF_X2 \mem_reg[29][24]  ( .D(n2065), .CK(clk), .Q(\mem[29][24] ) );
  DFF_X2 \mem_reg[29][23]  ( .D(n2064), .CK(clk), .Q(\mem[29][23] ) );
  DFF_X2 \mem_reg[29][22]  ( .D(n2063), .CK(clk), .Q(\mem[29][22] ) );
  DFF_X2 \mem_reg[29][21]  ( .D(n2062), .CK(clk), .Q(\mem[29][21] ) );
  DFF_X2 \mem_reg[29][20]  ( .D(n2061), .CK(clk), .Q(\mem[29][20] ) );
  DFF_X2 \mem_reg[29][19]  ( .D(n2060), .CK(clk), .Q(\mem[29][19] ) );
  DFF_X2 \mem_reg[29][18]  ( .D(n2059), .CK(clk), .Q(\mem[29][18] ) );
  DFF_X2 \mem_reg[29][17]  ( .D(n2058), .CK(clk), .Q(\mem[29][17] ) );
  DFF_X2 \mem_reg[29][16]  ( .D(n2057), .CK(clk), .Q(\mem[29][16] ) );
  DFF_X2 \mem_reg[29][15]  ( .D(n2056), .CK(clk), .Q(\mem[29][15] ) );
  DFF_X2 \mem_reg[29][14]  ( .D(n2055), .CK(clk), .Q(\mem[29][14] ) );
  DFF_X2 \mem_reg[29][13]  ( .D(n2054), .CK(clk), .Q(\mem[29][13] ) );
  DFF_X2 \mem_reg[29][12]  ( .D(n2053), .CK(clk), .Q(\mem[29][12] ) );
  DFF_X2 \mem_reg[29][11]  ( .D(n2052), .CK(clk), .Q(\mem[29][11] ) );
  DFF_X2 \mem_reg[29][10]  ( .D(n2051), .CK(clk), .Q(\mem[29][10] ) );
  DFF_X2 \mem_reg[29][9]  ( .D(n2050), .CK(clk), .Q(\mem[29][9] ) );
  DFF_X2 \mem_reg[29][8]  ( .D(n2049), .CK(clk), .Q(\mem[29][8] ) );
  DFF_X2 \mem_reg[29][7]  ( .D(n2048), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X2 \mem_reg[29][6]  ( .D(n2047), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X2 \mem_reg[29][5]  ( .D(n2046), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X2 \mem_reg[29][4]  ( .D(n2045), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X2 \mem_reg[29][3]  ( .D(n2044), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X2 \mem_reg[29][2]  ( .D(n2043), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X2 \mem_reg[29][1]  ( .D(n2042), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X2 \mem_reg[29][0]  ( .D(n2041), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X2 \mem_reg[28][31]  ( .D(n2040), .CK(clk), .Q(\mem[28][31] ) );
  DFF_X2 \mem_reg[28][30]  ( .D(n2039), .CK(clk), .Q(\mem[28][30] ) );
  DFF_X2 \mem_reg[28][29]  ( .D(n2038), .CK(clk), .Q(\mem[28][29] ) );
  DFF_X2 \mem_reg[28][28]  ( .D(n2037), .CK(clk), .Q(\mem[28][28] ) );
  DFF_X2 \mem_reg[28][27]  ( .D(n2036), .CK(clk), .Q(\mem[28][27] ) );
  DFF_X2 \mem_reg[28][26]  ( .D(n2035), .CK(clk), .Q(\mem[28][26] ) );
  DFF_X2 \mem_reg[28][25]  ( .D(n2034), .CK(clk), .Q(\mem[28][25] ) );
  DFF_X2 \mem_reg[28][24]  ( .D(n2033), .CK(clk), .Q(\mem[28][24] ) );
  DFF_X2 \mem_reg[28][23]  ( .D(n2032), .CK(clk), .Q(\mem[28][23] ) );
  DFF_X2 \mem_reg[28][22]  ( .D(n2031), .CK(clk), .Q(\mem[28][22] ) );
  DFF_X2 \mem_reg[28][21]  ( .D(n2030), .CK(clk), .Q(\mem[28][21] ) );
  DFF_X2 \mem_reg[28][20]  ( .D(n2029), .CK(clk), .Q(\mem[28][20] ) );
  DFF_X2 \mem_reg[28][19]  ( .D(n2028), .CK(clk), .Q(\mem[28][19] ) );
  DFF_X2 \mem_reg[28][18]  ( .D(n2027), .CK(clk), .Q(\mem[28][18] ) );
  DFF_X2 \mem_reg[28][17]  ( .D(n2026), .CK(clk), .Q(\mem[28][17] ) );
  DFF_X2 \mem_reg[28][16]  ( .D(n2025), .CK(clk), .Q(\mem[28][16] ) );
  DFF_X2 \mem_reg[28][15]  ( .D(n2024), .CK(clk), .Q(\mem[28][15] ) );
  DFF_X2 \mem_reg[28][14]  ( .D(n2023), .CK(clk), .Q(\mem[28][14] ) );
  DFF_X2 \mem_reg[28][13]  ( .D(n2022), .CK(clk), .Q(\mem[28][13] ) );
  DFF_X2 \mem_reg[28][12]  ( .D(n2021), .CK(clk), .Q(\mem[28][12] ) );
  DFF_X2 \mem_reg[28][11]  ( .D(n2020), .CK(clk), .Q(\mem[28][11] ) );
  DFF_X2 \mem_reg[28][10]  ( .D(n2019), .CK(clk), .Q(\mem[28][10] ) );
  DFF_X2 \mem_reg[28][9]  ( .D(n2018), .CK(clk), .Q(\mem[28][9] ) );
  DFF_X2 \mem_reg[28][8]  ( .D(n2017), .CK(clk), .Q(\mem[28][8] ) );
  DFF_X2 \mem_reg[28][7]  ( .D(n2016), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X2 \mem_reg[28][6]  ( .D(n2015), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X2 \mem_reg[28][5]  ( .D(n2014), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X2 \mem_reg[28][4]  ( .D(n2013), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X2 \mem_reg[28][3]  ( .D(n2012), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X2 \mem_reg[28][2]  ( .D(n2011), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X2 \mem_reg[28][1]  ( .D(n2010), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X2 \mem_reg[28][0]  ( .D(n2009), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X2 \mem_reg[27][31]  ( .D(n2008), .CK(clk), .Q(\mem[27][31] ) );
  DFF_X2 \mem_reg[27][30]  ( .D(n2007), .CK(clk), .Q(\mem[27][30] ) );
  DFF_X2 \mem_reg[27][29]  ( .D(n2006), .CK(clk), .Q(\mem[27][29] ) );
  DFF_X2 \mem_reg[27][28]  ( .D(n2005), .CK(clk), .Q(\mem[27][28] ) );
  DFF_X2 \mem_reg[27][27]  ( .D(n2004), .CK(clk), .Q(\mem[27][27] ) );
  DFF_X2 \mem_reg[27][26]  ( .D(n2003), .CK(clk), .Q(\mem[27][26] ) );
  DFF_X2 \mem_reg[27][25]  ( .D(n2002), .CK(clk), .Q(\mem[27][25] ) );
  DFF_X2 \mem_reg[27][24]  ( .D(n2001), .CK(clk), .Q(\mem[27][24] ) );
  DFF_X2 \mem_reg[27][23]  ( .D(n2000), .CK(clk), .Q(\mem[27][23] ) );
  DFF_X2 \mem_reg[27][22]  ( .D(n1999), .CK(clk), .Q(\mem[27][22] ) );
  DFF_X2 \mem_reg[27][21]  ( .D(n1998), .CK(clk), .Q(\mem[27][21] ) );
  DFF_X2 \mem_reg[27][20]  ( .D(n1997), .CK(clk), .Q(\mem[27][20] ) );
  DFF_X2 \mem_reg[27][19]  ( .D(n1996), .CK(clk), .Q(\mem[27][19] ) );
  DFF_X2 \mem_reg[27][18]  ( .D(n1995), .CK(clk), .Q(\mem[27][18] ) );
  DFF_X2 \mem_reg[27][17]  ( .D(n1994), .CK(clk), .Q(\mem[27][17] ) );
  DFF_X2 \mem_reg[27][16]  ( .D(n1993), .CK(clk), .Q(\mem[27][16] ) );
  DFF_X2 \mem_reg[27][15]  ( .D(n1992), .CK(clk), .Q(\mem[27][15] ) );
  DFF_X2 \mem_reg[27][14]  ( .D(n1991), .CK(clk), .Q(\mem[27][14] ) );
  DFF_X2 \mem_reg[27][13]  ( .D(n1990), .CK(clk), .Q(\mem[27][13] ) );
  DFF_X2 \mem_reg[27][12]  ( .D(n1989), .CK(clk), .Q(\mem[27][12] ) );
  DFF_X2 \mem_reg[27][11]  ( .D(n1988), .CK(clk), .Q(\mem[27][11] ) );
  DFF_X2 \mem_reg[27][10]  ( .D(n1987), .CK(clk), .Q(\mem[27][10] ) );
  DFF_X2 \mem_reg[27][9]  ( .D(n1986), .CK(clk), .Q(\mem[27][9] ) );
  DFF_X2 \mem_reg[27][8]  ( .D(n1985), .CK(clk), .Q(\mem[27][8] ) );
  DFF_X2 \mem_reg[27][7]  ( .D(n1984), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X2 \mem_reg[27][6]  ( .D(n1983), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X2 \mem_reg[27][5]  ( .D(n1982), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X2 \mem_reg[27][4]  ( .D(n1981), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X2 \mem_reg[27][3]  ( .D(n1980), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X2 \mem_reg[27][2]  ( .D(n1979), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X2 \mem_reg[27][1]  ( .D(n1978), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X2 \mem_reg[27][0]  ( .D(n1977), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X2 \mem_reg[26][31]  ( .D(n1976), .CK(clk), .Q(\mem[26][31] ) );
  DFF_X2 \mem_reg[26][30]  ( .D(n1975), .CK(clk), .Q(\mem[26][30] ) );
  DFF_X2 \mem_reg[26][29]  ( .D(n1974), .CK(clk), .Q(\mem[26][29] ) );
  DFF_X2 \mem_reg[26][28]  ( .D(n1973), .CK(clk), .Q(\mem[26][28] ) );
  DFF_X2 \mem_reg[26][27]  ( .D(n1972), .CK(clk), .Q(\mem[26][27] ) );
  DFF_X2 \mem_reg[26][26]  ( .D(n1971), .CK(clk), .Q(\mem[26][26] ) );
  DFF_X2 \mem_reg[26][25]  ( .D(n1970), .CK(clk), .Q(\mem[26][25] ) );
  DFF_X2 \mem_reg[26][24]  ( .D(n1969), .CK(clk), .Q(\mem[26][24] ) );
  DFF_X2 \mem_reg[26][23]  ( .D(n1968), .CK(clk), .Q(\mem[26][23] ) );
  DFF_X2 \mem_reg[26][22]  ( .D(n1967), .CK(clk), .Q(\mem[26][22] ) );
  DFF_X2 \mem_reg[26][21]  ( .D(n1966), .CK(clk), .Q(\mem[26][21] ) );
  DFF_X2 \mem_reg[26][20]  ( .D(n1965), .CK(clk), .Q(\mem[26][20] ) );
  DFF_X2 \mem_reg[26][19]  ( .D(n1964), .CK(clk), .Q(\mem[26][19] ) );
  DFF_X2 \mem_reg[26][18]  ( .D(n1963), .CK(clk), .Q(\mem[26][18] ) );
  DFF_X2 \mem_reg[26][17]  ( .D(n1962), .CK(clk), .Q(\mem[26][17] ) );
  DFF_X2 \mem_reg[26][16]  ( .D(n1961), .CK(clk), .Q(\mem[26][16] ) );
  DFF_X2 \mem_reg[26][15]  ( .D(n1960), .CK(clk), .Q(\mem[26][15] ) );
  DFF_X2 \mem_reg[26][14]  ( .D(n1959), .CK(clk), .Q(\mem[26][14] ) );
  DFF_X2 \mem_reg[26][13]  ( .D(n1958), .CK(clk), .Q(\mem[26][13] ) );
  DFF_X2 \mem_reg[26][12]  ( .D(n1957), .CK(clk), .Q(\mem[26][12] ) );
  DFF_X2 \mem_reg[26][11]  ( .D(n1956), .CK(clk), .Q(\mem[26][11] ) );
  DFF_X2 \mem_reg[26][10]  ( .D(n1955), .CK(clk), .Q(\mem[26][10] ) );
  DFF_X2 \mem_reg[26][9]  ( .D(n1954), .CK(clk), .Q(\mem[26][9] ) );
  DFF_X2 \mem_reg[26][8]  ( .D(n1953), .CK(clk), .Q(\mem[26][8] ) );
  DFF_X2 \mem_reg[26][7]  ( .D(n1952), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X2 \mem_reg[26][6]  ( .D(n1951), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X2 \mem_reg[26][5]  ( .D(n1950), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X2 \mem_reg[26][4]  ( .D(n1949), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X2 \mem_reg[26][3]  ( .D(n1948), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X2 \mem_reg[26][2]  ( .D(n1947), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X2 \mem_reg[26][1]  ( .D(n1946), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X2 \mem_reg[26][0]  ( .D(n1945), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X2 \mem_reg[25][31]  ( .D(n1944), .CK(clk), .Q(\mem[25][31] ) );
  DFF_X2 \mem_reg[25][30]  ( .D(n1943), .CK(clk), .Q(\mem[25][30] ) );
  DFF_X2 \mem_reg[25][29]  ( .D(n1942), .CK(clk), .Q(\mem[25][29] ) );
  DFF_X2 \mem_reg[25][28]  ( .D(n1941), .CK(clk), .Q(\mem[25][28] ) );
  DFF_X2 \mem_reg[25][27]  ( .D(n1940), .CK(clk), .Q(\mem[25][27] ) );
  DFF_X2 \mem_reg[25][26]  ( .D(n1939), .CK(clk), .Q(\mem[25][26] ) );
  DFF_X2 \mem_reg[25][25]  ( .D(n1938), .CK(clk), .Q(\mem[25][25] ) );
  DFF_X2 \mem_reg[25][24]  ( .D(n1937), .CK(clk), .Q(\mem[25][24] ) );
  DFF_X2 \mem_reg[25][23]  ( .D(n1936), .CK(clk), .Q(\mem[25][23] ) );
  DFF_X2 \mem_reg[25][22]  ( .D(n1935), .CK(clk), .Q(\mem[25][22] ) );
  DFF_X2 \mem_reg[25][21]  ( .D(n1934), .CK(clk), .Q(\mem[25][21] ) );
  DFF_X2 \mem_reg[25][20]  ( .D(n1933), .CK(clk), .Q(\mem[25][20] ) );
  DFF_X2 \mem_reg[25][19]  ( .D(n1932), .CK(clk), .Q(\mem[25][19] ) );
  DFF_X2 \mem_reg[25][18]  ( .D(n1931), .CK(clk), .Q(\mem[25][18] ) );
  DFF_X2 \mem_reg[25][17]  ( .D(n1930), .CK(clk), .Q(\mem[25][17] ) );
  DFF_X2 \mem_reg[25][16]  ( .D(n1929), .CK(clk), .Q(\mem[25][16] ) );
  DFF_X2 \mem_reg[25][15]  ( .D(n1928), .CK(clk), .Q(\mem[25][15] ) );
  DFF_X2 \mem_reg[25][14]  ( .D(n1927), .CK(clk), .Q(\mem[25][14] ) );
  DFF_X2 \mem_reg[25][13]  ( .D(n1926), .CK(clk), .Q(\mem[25][13] ) );
  DFF_X2 \mem_reg[25][12]  ( .D(n1925), .CK(clk), .Q(\mem[25][12] ) );
  DFF_X2 \mem_reg[25][11]  ( .D(n1924), .CK(clk), .Q(\mem[25][11] ) );
  DFF_X2 \mem_reg[25][10]  ( .D(n1923), .CK(clk), .Q(\mem[25][10] ) );
  DFF_X2 \mem_reg[25][9]  ( .D(n1922), .CK(clk), .Q(\mem[25][9] ) );
  DFF_X2 \mem_reg[25][8]  ( .D(n1921), .CK(clk), .Q(\mem[25][8] ) );
  DFF_X2 \mem_reg[25][7]  ( .D(n1920), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X2 \mem_reg[25][6]  ( .D(n1919), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X2 \mem_reg[25][5]  ( .D(n1918), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X2 \mem_reg[25][4]  ( .D(n1917), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X2 \mem_reg[25][3]  ( .D(n1916), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X2 \mem_reg[25][2]  ( .D(n1915), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X2 \mem_reg[25][1]  ( .D(n1914), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X2 \mem_reg[25][0]  ( .D(n1913), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X2 \mem_reg[24][31]  ( .D(n1912), .CK(clk), .Q(\mem[24][31] ) );
  DFF_X2 \mem_reg[24][30]  ( .D(n1911), .CK(clk), .Q(\mem[24][30] ) );
  DFF_X2 \mem_reg[24][29]  ( .D(n1910), .CK(clk), .Q(\mem[24][29] ) );
  DFF_X2 \mem_reg[24][28]  ( .D(n1909), .CK(clk), .Q(\mem[24][28] ) );
  DFF_X2 \mem_reg[24][27]  ( .D(n1908), .CK(clk), .Q(\mem[24][27] ) );
  DFF_X2 \mem_reg[24][26]  ( .D(n1907), .CK(clk), .Q(\mem[24][26] ) );
  DFF_X2 \mem_reg[24][25]  ( .D(n1906), .CK(clk), .Q(\mem[24][25] ) );
  DFF_X2 \mem_reg[24][24]  ( .D(n1905), .CK(clk), .Q(\mem[24][24] ) );
  DFF_X2 \mem_reg[24][23]  ( .D(n1904), .CK(clk), .Q(\mem[24][23] ) );
  DFF_X2 \mem_reg[24][22]  ( .D(n1903), .CK(clk), .Q(\mem[24][22] ) );
  DFF_X2 \mem_reg[24][21]  ( .D(n1902), .CK(clk), .Q(\mem[24][21] ) );
  DFF_X2 \mem_reg[24][20]  ( .D(n1901), .CK(clk), .Q(\mem[24][20] ) );
  DFF_X2 \mem_reg[24][19]  ( .D(n1900), .CK(clk), .Q(\mem[24][19] ) );
  DFF_X2 \mem_reg[24][18]  ( .D(n1899), .CK(clk), .Q(\mem[24][18] ) );
  DFF_X2 \mem_reg[24][17]  ( .D(n1898), .CK(clk), .Q(\mem[24][17] ) );
  DFF_X2 \mem_reg[24][16]  ( .D(n1897), .CK(clk), .Q(\mem[24][16] ) );
  DFF_X2 \mem_reg[24][15]  ( .D(n1896), .CK(clk), .Q(\mem[24][15] ) );
  DFF_X2 \mem_reg[24][14]  ( .D(n1895), .CK(clk), .Q(\mem[24][14] ) );
  DFF_X2 \mem_reg[24][13]  ( .D(n1894), .CK(clk), .Q(\mem[24][13] ) );
  DFF_X2 \mem_reg[24][12]  ( .D(n1893), .CK(clk), .Q(\mem[24][12] ) );
  DFF_X2 \mem_reg[24][11]  ( .D(n1892), .CK(clk), .Q(\mem[24][11] ) );
  DFF_X2 \mem_reg[24][10]  ( .D(n1891), .CK(clk), .Q(\mem[24][10] ) );
  DFF_X2 \mem_reg[24][9]  ( .D(n1890), .CK(clk), .Q(\mem[24][9] ) );
  DFF_X2 \mem_reg[24][8]  ( .D(n1889), .CK(clk), .Q(\mem[24][8] ) );
  DFF_X2 \mem_reg[24][7]  ( .D(n1888), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X2 \mem_reg[24][6]  ( .D(n1887), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X2 \mem_reg[24][5]  ( .D(n1886), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X2 \mem_reg[24][4]  ( .D(n1885), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X2 \mem_reg[24][3]  ( .D(n1884), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X2 \mem_reg[24][2]  ( .D(n1883), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X2 \mem_reg[24][1]  ( .D(n1882), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X2 \mem_reg[24][0]  ( .D(n1881), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X2 \mem_reg[23][31]  ( .D(n1880), .CK(clk), .Q(\mem[23][31] ) );
  DFF_X2 \mem_reg[23][30]  ( .D(n1879), .CK(clk), .Q(\mem[23][30] ) );
  DFF_X2 \mem_reg[23][29]  ( .D(n1878), .CK(clk), .Q(\mem[23][29] ) );
  DFF_X2 \mem_reg[23][28]  ( .D(n1877), .CK(clk), .Q(\mem[23][28] ) );
  DFF_X2 \mem_reg[23][27]  ( .D(n1876), .CK(clk), .Q(\mem[23][27] ) );
  DFF_X2 \mem_reg[23][26]  ( .D(n1875), .CK(clk), .Q(\mem[23][26] ) );
  DFF_X2 \mem_reg[23][25]  ( .D(n1874), .CK(clk), .Q(\mem[23][25] ) );
  DFF_X2 \mem_reg[23][24]  ( .D(n1873), .CK(clk), .Q(\mem[23][24] ) );
  DFF_X2 \mem_reg[23][23]  ( .D(n1872), .CK(clk), .Q(\mem[23][23] ) );
  DFF_X2 \mem_reg[23][22]  ( .D(n1871), .CK(clk), .Q(\mem[23][22] ) );
  DFF_X2 \mem_reg[23][21]  ( .D(n1870), .CK(clk), .Q(\mem[23][21] ) );
  DFF_X2 \mem_reg[23][20]  ( .D(n1869), .CK(clk), .Q(\mem[23][20] ) );
  DFF_X2 \mem_reg[23][19]  ( .D(n1868), .CK(clk), .Q(\mem[23][19] ) );
  DFF_X2 \mem_reg[23][18]  ( .D(n1867), .CK(clk), .Q(\mem[23][18] ) );
  DFF_X2 \mem_reg[23][17]  ( .D(n1866), .CK(clk), .Q(\mem[23][17] ) );
  DFF_X2 \mem_reg[23][16]  ( .D(n1865), .CK(clk), .Q(\mem[23][16] ) );
  DFF_X2 \mem_reg[23][15]  ( .D(n1864), .CK(clk), .Q(\mem[23][15] ) );
  DFF_X2 \mem_reg[23][14]  ( .D(n1863), .CK(clk), .Q(\mem[23][14] ) );
  DFF_X2 \mem_reg[23][13]  ( .D(n1862), .CK(clk), .Q(\mem[23][13] ) );
  DFF_X2 \mem_reg[23][12]  ( .D(n1861), .CK(clk), .Q(\mem[23][12] ) );
  DFF_X2 \mem_reg[23][11]  ( .D(n1860), .CK(clk), .Q(\mem[23][11] ) );
  DFF_X2 \mem_reg[23][10]  ( .D(n1859), .CK(clk), .Q(\mem[23][10] ) );
  DFF_X2 \mem_reg[23][9]  ( .D(n1858), .CK(clk), .Q(\mem[23][9] ) );
  DFF_X2 \mem_reg[23][8]  ( .D(n1857), .CK(clk), .Q(\mem[23][8] ) );
  DFF_X2 \mem_reg[23][7]  ( .D(n1856), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X2 \mem_reg[23][6]  ( .D(n1855), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X2 \mem_reg[23][5]  ( .D(n1854), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X2 \mem_reg[23][4]  ( .D(n1853), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X2 \mem_reg[23][3]  ( .D(n1852), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X2 \mem_reg[23][2]  ( .D(n1851), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X2 \mem_reg[23][1]  ( .D(n1850), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X2 \mem_reg[23][0]  ( .D(n1849), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X2 \mem_reg[22][31]  ( .D(n1848), .CK(clk), .Q(\mem[22][31] ) );
  DFF_X2 \mem_reg[22][30]  ( .D(n1847), .CK(clk), .Q(\mem[22][30] ) );
  DFF_X2 \mem_reg[22][29]  ( .D(n1846), .CK(clk), .Q(\mem[22][29] ) );
  DFF_X2 \mem_reg[22][28]  ( .D(n1845), .CK(clk), .Q(\mem[22][28] ) );
  DFF_X2 \mem_reg[22][27]  ( .D(n1844), .CK(clk), .Q(\mem[22][27] ) );
  DFF_X2 \mem_reg[22][26]  ( .D(n1843), .CK(clk), .Q(\mem[22][26] ) );
  DFF_X2 \mem_reg[22][25]  ( .D(n1842), .CK(clk), .Q(\mem[22][25] ) );
  DFF_X2 \mem_reg[22][24]  ( .D(n1841), .CK(clk), .Q(\mem[22][24] ) );
  DFF_X2 \mem_reg[22][23]  ( .D(n1840), .CK(clk), .Q(\mem[22][23] ) );
  DFF_X2 \mem_reg[22][22]  ( .D(n1839), .CK(clk), .Q(\mem[22][22] ) );
  DFF_X2 \mem_reg[22][21]  ( .D(n1838), .CK(clk), .Q(\mem[22][21] ) );
  DFF_X2 \mem_reg[22][20]  ( .D(n1837), .CK(clk), .Q(\mem[22][20] ) );
  DFF_X2 \mem_reg[22][19]  ( .D(n1836), .CK(clk), .Q(\mem[22][19] ) );
  DFF_X2 \mem_reg[22][18]  ( .D(n1835), .CK(clk), .Q(\mem[22][18] ) );
  DFF_X2 \mem_reg[22][17]  ( .D(n1834), .CK(clk), .Q(\mem[22][17] ) );
  DFF_X2 \mem_reg[22][16]  ( .D(n1833), .CK(clk), .Q(\mem[22][16] ) );
  DFF_X2 \mem_reg[22][15]  ( .D(n1832), .CK(clk), .Q(\mem[22][15] ) );
  DFF_X2 \mem_reg[22][14]  ( .D(n1831), .CK(clk), .Q(\mem[22][14] ) );
  DFF_X2 \mem_reg[22][13]  ( .D(n1830), .CK(clk), .Q(\mem[22][13] ) );
  DFF_X2 \mem_reg[22][12]  ( .D(n1829), .CK(clk), .Q(\mem[22][12] ) );
  DFF_X2 \mem_reg[22][11]  ( .D(n1828), .CK(clk), .Q(\mem[22][11] ) );
  DFF_X2 \mem_reg[22][10]  ( .D(n1827), .CK(clk), .Q(\mem[22][10] ) );
  DFF_X2 \mem_reg[22][9]  ( .D(n1826), .CK(clk), .Q(\mem[22][9] ) );
  DFF_X2 \mem_reg[22][8]  ( .D(n1825), .CK(clk), .Q(\mem[22][8] ) );
  DFF_X2 \mem_reg[22][7]  ( .D(n1824), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X2 \mem_reg[22][6]  ( .D(n1823), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X2 \mem_reg[22][5]  ( .D(n1822), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X2 \mem_reg[22][4]  ( .D(n1821), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X2 \mem_reg[22][3]  ( .D(n1820), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X2 \mem_reg[22][2]  ( .D(n1819), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X2 \mem_reg[22][1]  ( .D(n1818), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X2 \mem_reg[22][0]  ( .D(n1817), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X2 \mem_reg[21][31]  ( .D(n1816), .CK(clk), .Q(\mem[21][31] ) );
  DFF_X2 \mem_reg[21][30]  ( .D(n1815), .CK(clk), .Q(\mem[21][30] ) );
  DFF_X2 \mem_reg[21][29]  ( .D(n1814), .CK(clk), .Q(\mem[21][29] ) );
  DFF_X2 \mem_reg[21][28]  ( .D(n1813), .CK(clk), .Q(\mem[21][28] ) );
  DFF_X2 \mem_reg[21][27]  ( .D(n1812), .CK(clk), .Q(\mem[21][27] ) );
  DFF_X2 \mem_reg[21][26]  ( .D(n1811), .CK(clk), .Q(\mem[21][26] ) );
  DFF_X2 \mem_reg[21][25]  ( .D(n1810), .CK(clk), .Q(\mem[21][25] ) );
  DFF_X2 \mem_reg[21][24]  ( .D(n1809), .CK(clk), .Q(\mem[21][24] ) );
  DFF_X2 \mem_reg[21][23]  ( .D(n1808), .CK(clk), .Q(\mem[21][23] ) );
  DFF_X2 \mem_reg[21][22]  ( .D(n1807), .CK(clk), .Q(\mem[21][22] ) );
  DFF_X2 \mem_reg[21][21]  ( .D(n1806), .CK(clk), .Q(\mem[21][21] ) );
  DFF_X2 \mem_reg[21][20]  ( .D(n1805), .CK(clk), .Q(\mem[21][20] ) );
  DFF_X2 \mem_reg[21][19]  ( .D(n1804), .CK(clk), .Q(\mem[21][19] ) );
  DFF_X2 \mem_reg[21][18]  ( .D(n1803), .CK(clk), .Q(\mem[21][18] ) );
  DFF_X2 \mem_reg[21][17]  ( .D(n1802), .CK(clk), .Q(\mem[21][17] ) );
  DFF_X2 \mem_reg[21][16]  ( .D(n1801), .CK(clk), .Q(\mem[21][16] ) );
  DFF_X2 \mem_reg[21][15]  ( .D(n1800), .CK(clk), .Q(\mem[21][15] ) );
  DFF_X2 \mem_reg[21][14]  ( .D(n1799), .CK(clk), .Q(\mem[21][14] ) );
  DFF_X2 \mem_reg[21][13]  ( .D(n1798), .CK(clk), .Q(\mem[21][13] ) );
  DFF_X2 \mem_reg[21][12]  ( .D(n1797), .CK(clk), .Q(\mem[21][12] ) );
  DFF_X2 \mem_reg[21][11]  ( .D(n1796), .CK(clk), .Q(\mem[21][11] ) );
  DFF_X2 \mem_reg[21][10]  ( .D(n1795), .CK(clk), .Q(\mem[21][10] ) );
  DFF_X2 \mem_reg[21][9]  ( .D(n1794), .CK(clk), .Q(\mem[21][9] ) );
  DFF_X2 \mem_reg[21][8]  ( .D(n1793), .CK(clk), .Q(\mem[21][8] ) );
  DFF_X2 \mem_reg[21][7]  ( .D(n1792), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X2 \mem_reg[21][6]  ( .D(n1791), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X2 \mem_reg[21][5]  ( .D(n1790), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X2 \mem_reg[21][4]  ( .D(n1789), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X2 \mem_reg[21][3]  ( .D(n1788), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X2 \mem_reg[21][2]  ( .D(n1787), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X2 \mem_reg[21][1]  ( .D(n1786), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X2 \mem_reg[21][0]  ( .D(n1785), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X2 \mem_reg[20][31]  ( .D(n1784), .CK(clk), .Q(\mem[20][31] ) );
  DFF_X2 \mem_reg[20][30]  ( .D(n1783), .CK(clk), .Q(\mem[20][30] ) );
  DFF_X2 \mem_reg[20][29]  ( .D(n1782), .CK(clk), .Q(\mem[20][29] ) );
  DFF_X2 \mem_reg[20][28]  ( .D(n1781), .CK(clk), .Q(\mem[20][28] ) );
  DFF_X2 \mem_reg[20][27]  ( .D(n1780), .CK(clk), .Q(\mem[20][27] ) );
  DFF_X2 \mem_reg[20][26]  ( .D(n1779), .CK(clk), .Q(\mem[20][26] ) );
  DFF_X2 \mem_reg[20][25]  ( .D(n1778), .CK(clk), .Q(\mem[20][25] ) );
  DFF_X2 \mem_reg[20][24]  ( .D(n1777), .CK(clk), .Q(\mem[20][24] ) );
  DFF_X2 \mem_reg[20][23]  ( .D(n1776), .CK(clk), .Q(\mem[20][23] ) );
  DFF_X2 \mem_reg[20][22]  ( .D(n1775), .CK(clk), .Q(\mem[20][22] ) );
  DFF_X2 \mem_reg[20][21]  ( .D(n1774), .CK(clk), .Q(\mem[20][21] ) );
  DFF_X2 \mem_reg[20][20]  ( .D(n1773), .CK(clk), .Q(\mem[20][20] ) );
  DFF_X2 \mem_reg[20][19]  ( .D(n1772), .CK(clk), .Q(\mem[20][19] ) );
  DFF_X2 \mem_reg[20][18]  ( .D(n1771), .CK(clk), .Q(\mem[20][18] ) );
  DFF_X2 \mem_reg[20][17]  ( .D(n1770), .CK(clk), .Q(\mem[20][17] ) );
  DFF_X2 \mem_reg[20][16]  ( .D(n1769), .CK(clk), .Q(\mem[20][16] ) );
  DFF_X2 \mem_reg[20][15]  ( .D(n1768), .CK(clk), .Q(\mem[20][15] ) );
  DFF_X2 \mem_reg[20][14]  ( .D(n1767), .CK(clk), .Q(\mem[20][14] ) );
  DFF_X2 \mem_reg[20][13]  ( .D(n1766), .CK(clk), .Q(\mem[20][13] ) );
  DFF_X2 \mem_reg[20][12]  ( .D(n1765), .CK(clk), .Q(\mem[20][12] ) );
  DFF_X2 \mem_reg[20][11]  ( .D(n1764), .CK(clk), .Q(\mem[20][11] ) );
  DFF_X2 \mem_reg[20][10]  ( .D(n1763), .CK(clk), .Q(\mem[20][10] ) );
  DFF_X2 \mem_reg[20][9]  ( .D(n1762), .CK(clk), .Q(\mem[20][9] ) );
  DFF_X2 \mem_reg[20][8]  ( .D(n1761), .CK(clk), .Q(\mem[20][8] ) );
  DFF_X2 \mem_reg[20][7]  ( .D(n1760), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X2 \mem_reg[20][6]  ( .D(n1759), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X2 \mem_reg[20][5]  ( .D(n1758), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X2 \mem_reg[20][4]  ( .D(n1757), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X2 \mem_reg[20][3]  ( .D(n1756), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X2 \mem_reg[20][2]  ( .D(n1755), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X2 \mem_reg[20][1]  ( .D(n1754), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X2 \mem_reg[20][0]  ( .D(n1753), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X2 \mem_reg[19][31]  ( .D(n1752), .CK(clk), .Q(\mem[19][31] ) );
  DFF_X2 \mem_reg[19][30]  ( .D(n1751), .CK(clk), .Q(\mem[19][30] ) );
  DFF_X2 \mem_reg[19][29]  ( .D(n1750), .CK(clk), .Q(\mem[19][29] ) );
  DFF_X2 \mem_reg[19][28]  ( .D(n1749), .CK(clk), .Q(\mem[19][28] ) );
  DFF_X2 \mem_reg[19][27]  ( .D(n1748), .CK(clk), .Q(\mem[19][27] ) );
  DFF_X2 \mem_reg[19][26]  ( .D(n1747), .CK(clk), .Q(\mem[19][26] ) );
  DFF_X2 \mem_reg[19][25]  ( .D(n1746), .CK(clk), .Q(\mem[19][25] ) );
  DFF_X2 \mem_reg[19][24]  ( .D(n1745), .CK(clk), .Q(\mem[19][24] ) );
  DFF_X2 \mem_reg[19][23]  ( .D(n1744), .CK(clk), .Q(\mem[19][23] ) );
  DFF_X2 \mem_reg[19][22]  ( .D(n1743), .CK(clk), .Q(\mem[19][22] ) );
  DFF_X2 \mem_reg[19][21]  ( .D(n1742), .CK(clk), .Q(\mem[19][21] ) );
  DFF_X2 \mem_reg[19][20]  ( .D(n1741), .CK(clk), .Q(\mem[19][20] ) );
  DFF_X2 \mem_reg[19][19]  ( .D(n1740), .CK(clk), .Q(\mem[19][19] ) );
  DFF_X2 \mem_reg[19][18]  ( .D(n1739), .CK(clk), .Q(\mem[19][18] ) );
  DFF_X2 \mem_reg[19][17]  ( .D(n1738), .CK(clk), .Q(\mem[19][17] ) );
  DFF_X2 \mem_reg[19][16]  ( .D(n1737), .CK(clk), .Q(\mem[19][16] ) );
  DFF_X2 \mem_reg[19][15]  ( .D(n1736), .CK(clk), .Q(\mem[19][15] ) );
  DFF_X2 \mem_reg[19][14]  ( .D(n1735), .CK(clk), .Q(\mem[19][14] ) );
  DFF_X2 \mem_reg[19][13]  ( .D(n1734), .CK(clk), .Q(\mem[19][13] ) );
  DFF_X2 \mem_reg[19][12]  ( .D(n1733), .CK(clk), .Q(\mem[19][12] ) );
  DFF_X2 \mem_reg[19][11]  ( .D(n1732), .CK(clk), .Q(\mem[19][11] ) );
  DFF_X2 \mem_reg[19][10]  ( .D(n1731), .CK(clk), .Q(\mem[19][10] ) );
  DFF_X2 \mem_reg[19][9]  ( .D(n1730), .CK(clk), .Q(\mem[19][9] ) );
  DFF_X2 \mem_reg[19][8]  ( .D(n1729), .CK(clk), .Q(\mem[19][8] ) );
  DFF_X2 \mem_reg[19][7]  ( .D(n1728), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X2 \mem_reg[19][6]  ( .D(n1727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X2 \mem_reg[19][5]  ( .D(n1726), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X2 \mem_reg[19][4]  ( .D(n1725), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X2 \mem_reg[19][3]  ( .D(n1724), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X2 \mem_reg[19][2]  ( .D(n1723), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X2 \mem_reg[19][1]  ( .D(n1722), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X2 \mem_reg[19][0]  ( .D(n1721), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X2 \mem_reg[18][31]  ( .D(n1720), .CK(clk), .Q(\mem[18][31] ) );
  DFF_X2 \mem_reg[18][30]  ( .D(n1719), .CK(clk), .Q(\mem[18][30] ) );
  DFF_X2 \mem_reg[18][29]  ( .D(n1718), .CK(clk), .Q(\mem[18][29] ) );
  DFF_X2 \mem_reg[18][28]  ( .D(n1717), .CK(clk), .Q(\mem[18][28] ) );
  DFF_X2 \mem_reg[18][27]  ( .D(n1716), .CK(clk), .Q(\mem[18][27] ) );
  DFF_X2 \mem_reg[18][26]  ( .D(n1715), .CK(clk), .Q(\mem[18][26] ) );
  DFF_X2 \mem_reg[18][25]  ( .D(n1714), .CK(clk), .Q(\mem[18][25] ) );
  DFF_X2 \mem_reg[18][24]  ( .D(n1713), .CK(clk), .Q(\mem[18][24] ) );
  DFF_X2 \mem_reg[18][23]  ( .D(n1712), .CK(clk), .Q(\mem[18][23] ) );
  DFF_X2 \mem_reg[18][22]  ( .D(n1711), .CK(clk), .Q(\mem[18][22] ) );
  DFF_X2 \mem_reg[18][21]  ( .D(n1710), .CK(clk), .Q(\mem[18][21] ) );
  DFF_X2 \mem_reg[18][20]  ( .D(n1709), .CK(clk), .Q(\mem[18][20] ) );
  DFF_X2 \mem_reg[18][19]  ( .D(n1708), .CK(clk), .Q(\mem[18][19] ) );
  DFF_X2 \mem_reg[18][18]  ( .D(n1707), .CK(clk), .Q(\mem[18][18] ) );
  DFF_X2 \mem_reg[18][17]  ( .D(n1706), .CK(clk), .Q(\mem[18][17] ) );
  DFF_X2 \mem_reg[18][16]  ( .D(n1705), .CK(clk), .Q(\mem[18][16] ) );
  DFF_X2 \mem_reg[18][15]  ( .D(n1704), .CK(clk), .Q(\mem[18][15] ) );
  DFF_X2 \mem_reg[18][14]  ( .D(n1703), .CK(clk), .Q(\mem[18][14] ) );
  DFF_X2 \mem_reg[18][13]  ( .D(n1702), .CK(clk), .Q(\mem[18][13] ) );
  DFF_X2 \mem_reg[18][12]  ( .D(n1701), .CK(clk), .Q(\mem[18][12] ) );
  DFF_X2 \mem_reg[18][11]  ( .D(n1700), .CK(clk), .Q(\mem[18][11] ) );
  DFF_X2 \mem_reg[18][10]  ( .D(n1699), .CK(clk), .Q(\mem[18][10] ) );
  DFF_X2 \mem_reg[18][9]  ( .D(n1698), .CK(clk), .Q(\mem[18][9] ) );
  DFF_X2 \mem_reg[18][8]  ( .D(n1697), .CK(clk), .Q(\mem[18][8] ) );
  DFF_X2 \mem_reg[18][7]  ( .D(n1696), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X2 \mem_reg[18][6]  ( .D(n1695), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X2 \mem_reg[18][5]  ( .D(n1694), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X2 \mem_reg[18][4]  ( .D(n1693), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X2 \mem_reg[18][3]  ( .D(n1692), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X2 \mem_reg[18][2]  ( .D(n1691), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X2 \mem_reg[18][1]  ( .D(n1690), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X2 \mem_reg[18][0]  ( .D(n1689), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X2 \mem_reg[17][31]  ( .D(n1688), .CK(clk), .Q(\mem[17][31] ) );
  DFF_X2 \mem_reg[17][30]  ( .D(n1687), .CK(clk), .Q(\mem[17][30] ) );
  DFF_X2 \mem_reg[17][29]  ( .D(n1686), .CK(clk), .Q(\mem[17][29] ) );
  DFF_X2 \mem_reg[17][28]  ( .D(n1685), .CK(clk), .Q(\mem[17][28] ) );
  DFF_X2 \mem_reg[17][27]  ( .D(n1684), .CK(clk), .Q(\mem[17][27] ) );
  DFF_X2 \mem_reg[17][26]  ( .D(n1683), .CK(clk), .Q(\mem[17][26] ) );
  DFF_X2 \mem_reg[17][25]  ( .D(n1682), .CK(clk), .Q(\mem[17][25] ) );
  DFF_X2 \mem_reg[17][24]  ( .D(n1681), .CK(clk), .Q(\mem[17][24] ) );
  DFF_X2 \mem_reg[17][23]  ( .D(n1680), .CK(clk), .Q(\mem[17][23] ) );
  DFF_X2 \mem_reg[17][22]  ( .D(n1679), .CK(clk), .Q(\mem[17][22] ) );
  DFF_X2 \mem_reg[17][21]  ( .D(n1678), .CK(clk), .Q(\mem[17][21] ) );
  DFF_X2 \mem_reg[17][20]  ( .D(n1677), .CK(clk), .Q(\mem[17][20] ) );
  DFF_X2 \mem_reg[17][19]  ( .D(n1676), .CK(clk), .Q(\mem[17][19] ) );
  DFF_X2 \mem_reg[17][18]  ( .D(n1675), .CK(clk), .Q(\mem[17][18] ) );
  DFF_X2 \mem_reg[17][17]  ( .D(n1674), .CK(clk), .Q(\mem[17][17] ) );
  DFF_X2 \mem_reg[17][16]  ( .D(n1673), .CK(clk), .Q(\mem[17][16] ) );
  DFF_X2 \mem_reg[17][15]  ( .D(n1672), .CK(clk), .Q(\mem[17][15] ) );
  DFF_X2 \mem_reg[17][14]  ( .D(n1671), .CK(clk), .Q(\mem[17][14] ) );
  DFF_X2 \mem_reg[17][13]  ( .D(n1670), .CK(clk), .Q(\mem[17][13] ) );
  DFF_X2 \mem_reg[17][12]  ( .D(n1669), .CK(clk), .Q(\mem[17][12] ) );
  DFF_X2 \mem_reg[17][11]  ( .D(n1668), .CK(clk), .Q(\mem[17][11] ) );
  DFF_X2 \mem_reg[17][10]  ( .D(n1667), .CK(clk), .Q(\mem[17][10] ) );
  DFF_X2 \mem_reg[17][9]  ( .D(n1666), .CK(clk), .Q(\mem[17][9] ) );
  DFF_X2 \mem_reg[17][8]  ( .D(n1665), .CK(clk), .Q(\mem[17][8] ) );
  DFF_X2 \mem_reg[17][7]  ( .D(n1664), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X2 \mem_reg[17][6]  ( .D(n1663), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X2 \mem_reg[17][5]  ( .D(n1662), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X2 \mem_reg[17][4]  ( .D(n1661), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X2 \mem_reg[17][3]  ( .D(n1660), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X2 \mem_reg[17][2]  ( .D(n1659), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X2 \mem_reg[17][1]  ( .D(n1658), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X2 \mem_reg[17][0]  ( .D(n1657), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X2 \mem_reg[16][31]  ( .D(n1656), .CK(clk), .Q(\mem[16][31] ) );
  DFF_X2 \mem_reg[16][30]  ( .D(n1655), .CK(clk), .Q(\mem[16][30] ) );
  DFF_X2 \mem_reg[16][29]  ( .D(n1654), .CK(clk), .Q(\mem[16][29] ) );
  DFF_X2 \mem_reg[16][28]  ( .D(n1653), .CK(clk), .Q(\mem[16][28] ) );
  DFF_X2 \mem_reg[16][27]  ( .D(n1652), .CK(clk), .Q(\mem[16][27] ) );
  DFF_X2 \mem_reg[16][26]  ( .D(n1651), .CK(clk), .Q(\mem[16][26] ) );
  DFF_X2 \mem_reg[16][25]  ( .D(n1650), .CK(clk), .Q(\mem[16][25] ) );
  DFF_X2 \mem_reg[16][24]  ( .D(n1649), .CK(clk), .Q(\mem[16][24] ) );
  DFF_X2 \mem_reg[16][23]  ( .D(n1648), .CK(clk), .Q(\mem[16][23] ) );
  DFF_X2 \mem_reg[16][22]  ( .D(n1647), .CK(clk), .Q(\mem[16][22] ) );
  DFF_X2 \mem_reg[16][21]  ( .D(n1646), .CK(clk), .Q(\mem[16][21] ) );
  DFF_X2 \mem_reg[16][20]  ( .D(n1645), .CK(clk), .Q(\mem[16][20] ) );
  DFF_X2 \mem_reg[16][19]  ( .D(n1644), .CK(clk), .Q(\mem[16][19] ) );
  DFF_X2 \mem_reg[16][18]  ( .D(n1643), .CK(clk), .Q(\mem[16][18] ) );
  DFF_X2 \mem_reg[16][17]  ( .D(n1642), .CK(clk), .Q(\mem[16][17] ) );
  DFF_X2 \mem_reg[16][16]  ( .D(n1641), .CK(clk), .Q(\mem[16][16] ) );
  DFF_X2 \mem_reg[16][15]  ( .D(n1640), .CK(clk), .Q(\mem[16][15] ) );
  DFF_X2 \mem_reg[16][14]  ( .D(n1639), .CK(clk), .Q(\mem[16][14] ) );
  DFF_X2 \mem_reg[16][13]  ( .D(n1638), .CK(clk), .Q(\mem[16][13] ) );
  DFF_X2 \mem_reg[16][12]  ( .D(n1637), .CK(clk), .Q(\mem[16][12] ) );
  DFF_X2 \mem_reg[16][11]  ( .D(n1636), .CK(clk), .Q(\mem[16][11] ) );
  DFF_X2 \mem_reg[16][10]  ( .D(n1635), .CK(clk), .Q(\mem[16][10] ) );
  DFF_X2 \mem_reg[16][9]  ( .D(n1634), .CK(clk), .Q(\mem[16][9] ) );
  DFF_X2 \mem_reg[16][8]  ( .D(n1633), .CK(clk), .Q(\mem[16][8] ) );
  DFF_X2 \mem_reg[16][7]  ( .D(n1632), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X2 \mem_reg[16][6]  ( .D(n1631), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X2 \mem_reg[16][5]  ( .D(n1630), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X2 \mem_reg[16][4]  ( .D(n1629), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X2 \mem_reg[16][3]  ( .D(n1628), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X2 \mem_reg[16][2]  ( .D(n1627), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X2 \mem_reg[16][1]  ( .D(n1626), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X2 \mem_reg[16][0]  ( .D(n1625), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X2 \mem_reg[15][31]  ( .D(n1624), .CK(clk), .Q(\mem[15][31] ) );
  DFF_X2 \mem_reg[15][30]  ( .D(n1623), .CK(clk), .Q(\mem[15][30] ) );
  DFF_X2 \mem_reg[15][29]  ( .D(n1622), .CK(clk), .Q(\mem[15][29] ) );
  DFF_X2 \mem_reg[15][28]  ( .D(n1621), .CK(clk), .Q(\mem[15][28] ) );
  DFF_X2 \mem_reg[15][27]  ( .D(n1620), .CK(clk), .Q(\mem[15][27] ) );
  DFF_X2 \mem_reg[15][26]  ( .D(n1619), .CK(clk), .Q(\mem[15][26] ) );
  DFF_X2 \mem_reg[15][25]  ( .D(n1618), .CK(clk), .Q(\mem[15][25] ) );
  DFF_X2 \mem_reg[15][24]  ( .D(n1617), .CK(clk), .Q(\mem[15][24] ) );
  DFF_X2 \mem_reg[15][23]  ( .D(n1616), .CK(clk), .Q(\mem[15][23] ) );
  DFF_X2 \mem_reg[15][22]  ( .D(n1615), .CK(clk), .Q(\mem[15][22] ) );
  DFF_X2 \mem_reg[15][21]  ( .D(n1614), .CK(clk), .Q(\mem[15][21] ) );
  DFF_X2 \mem_reg[15][20]  ( .D(n1613), .CK(clk), .Q(\mem[15][20] ) );
  DFF_X2 \mem_reg[15][19]  ( .D(n1612), .CK(clk), .Q(\mem[15][19] ) );
  DFF_X2 \mem_reg[15][18]  ( .D(n1611), .CK(clk), .Q(\mem[15][18] ) );
  DFF_X2 \mem_reg[15][17]  ( .D(n1610), .CK(clk), .Q(\mem[15][17] ) );
  DFF_X2 \mem_reg[15][16]  ( .D(n1609), .CK(clk), .Q(\mem[15][16] ) );
  DFF_X2 \mem_reg[15][15]  ( .D(n1608), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X2 \mem_reg[15][14]  ( .D(n1607), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X2 \mem_reg[15][13]  ( .D(n1606), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X2 \mem_reg[15][12]  ( .D(n1605), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X2 \mem_reg[15][11]  ( .D(n1604), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X2 \mem_reg[15][10]  ( .D(n1603), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X2 \mem_reg[15][9]  ( .D(n1602), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X2 \mem_reg[15][8]  ( .D(n1601), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X2 \mem_reg[15][7]  ( .D(n1600), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X2 \mem_reg[15][6]  ( .D(n1599), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X2 \mem_reg[15][5]  ( .D(n1598), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X2 \mem_reg[15][4]  ( .D(n1597), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X2 \mem_reg[15][3]  ( .D(n1596), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X2 \mem_reg[15][2]  ( .D(n1595), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X2 \mem_reg[15][1]  ( .D(n1594), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X2 \mem_reg[15][0]  ( .D(n1593), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X2 \mem_reg[14][31]  ( .D(n1592), .CK(clk), .Q(\mem[14][31] ) );
  DFF_X2 \mem_reg[14][30]  ( .D(n1591), .CK(clk), .Q(\mem[14][30] ) );
  DFF_X2 \mem_reg[14][29]  ( .D(n1590), .CK(clk), .Q(\mem[14][29] ) );
  DFF_X2 \mem_reg[14][28]  ( .D(n1589), .CK(clk), .Q(\mem[14][28] ) );
  DFF_X2 \mem_reg[14][27]  ( .D(n1588), .CK(clk), .Q(\mem[14][27] ) );
  DFF_X2 \mem_reg[14][26]  ( .D(n1587), .CK(clk), .Q(\mem[14][26] ) );
  DFF_X2 \mem_reg[14][25]  ( .D(n1586), .CK(clk), .Q(\mem[14][25] ) );
  DFF_X2 \mem_reg[14][24]  ( .D(n1585), .CK(clk), .Q(\mem[14][24] ) );
  DFF_X2 \mem_reg[14][23]  ( .D(n1584), .CK(clk), .Q(\mem[14][23] ) );
  DFF_X2 \mem_reg[14][22]  ( .D(n1583), .CK(clk), .Q(\mem[14][22] ) );
  DFF_X2 \mem_reg[14][21]  ( .D(n1582), .CK(clk), .Q(\mem[14][21] ) );
  DFF_X2 \mem_reg[14][20]  ( .D(n1581), .CK(clk), .Q(\mem[14][20] ) );
  DFF_X2 \mem_reg[14][19]  ( .D(n1580), .CK(clk), .Q(\mem[14][19] ) );
  DFF_X2 \mem_reg[14][18]  ( .D(n1579), .CK(clk), .Q(\mem[14][18] ) );
  DFF_X2 \mem_reg[14][17]  ( .D(n1578), .CK(clk), .Q(\mem[14][17] ) );
  DFF_X2 \mem_reg[14][16]  ( .D(n1577), .CK(clk), .Q(\mem[14][16] ) );
  DFF_X2 \mem_reg[14][15]  ( .D(n1576), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X2 \mem_reg[14][14]  ( .D(n1575), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X2 \mem_reg[14][13]  ( .D(n1574), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X2 \mem_reg[14][12]  ( .D(n1573), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X2 \mem_reg[14][11]  ( .D(n1572), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X2 \mem_reg[14][10]  ( .D(n1571), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X2 \mem_reg[14][9]  ( .D(n1570), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X2 \mem_reg[14][8]  ( .D(n1569), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X2 \mem_reg[14][7]  ( .D(n1568), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X2 \mem_reg[14][6]  ( .D(n1567), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X2 \mem_reg[14][5]  ( .D(n1566), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X2 \mem_reg[14][4]  ( .D(n1565), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X2 \mem_reg[14][3]  ( .D(n1564), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X2 \mem_reg[14][2]  ( .D(n1563), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X2 \mem_reg[14][1]  ( .D(n1562), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X2 \mem_reg[14][0]  ( .D(n1561), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X2 \mem_reg[13][31]  ( .D(n1560), .CK(clk), .Q(\mem[13][31] ) );
  DFF_X2 \mem_reg[13][30]  ( .D(n1559), .CK(clk), .Q(\mem[13][30] ) );
  DFF_X2 \mem_reg[13][29]  ( .D(n1558), .CK(clk), .Q(\mem[13][29] ) );
  DFF_X2 \mem_reg[13][28]  ( .D(n1557), .CK(clk), .Q(\mem[13][28] ) );
  DFF_X2 \mem_reg[13][27]  ( .D(n1556), .CK(clk), .Q(\mem[13][27] ) );
  DFF_X2 \mem_reg[13][26]  ( .D(n1555), .CK(clk), .Q(\mem[13][26] ) );
  DFF_X2 \mem_reg[13][25]  ( .D(n1554), .CK(clk), .Q(\mem[13][25] ) );
  DFF_X2 \mem_reg[13][24]  ( .D(n1553), .CK(clk), .Q(\mem[13][24] ) );
  DFF_X2 \mem_reg[13][23]  ( .D(n1552), .CK(clk), .Q(\mem[13][23] ) );
  DFF_X2 \mem_reg[13][22]  ( .D(n1551), .CK(clk), .Q(\mem[13][22] ) );
  DFF_X2 \mem_reg[13][21]  ( .D(n1550), .CK(clk), .Q(\mem[13][21] ) );
  DFF_X2 \mem_reg[13][20]  ( .D(n1549), .CK(clk), .Q(\mem[13][20] ) );
  DFF_X2 \mem_reg[13][19]  ( .D(n1548), .CK(clk), .Q(\mem[13][19] ) );
  DFF_X2 \mem_reg[13][18]  ( .D(n1547), .CK(clk), .Q(\mem[13][18] ) );
  DFF_X2 \mem_reg[13][17]  ( .D(n1546), .CK(clk), .Q(\mem[13][17] ) );
  DFF_X2 \mem_reg[13][16]  ( .D(n1545), .CK(clk), .Q(\mem[13][16] ) );
  DFF_X2 \mem_reg[13][15]  ( .D(n1544), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X2 \mem_reg[13][14]  ( .D(n1543), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X2 \mem_reg[13][13]  ( .D(n1542), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X2 \mem_reg[13][12]  ( .D(n1541), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X2 \mem_reg[13][11]  ( .D(n1540), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X2 \mem_reg[13][10]  ( .D(n1539), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X2 \mem_reg[13][9]  ( .D(n1538), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X2 \mem_reg[13][8]  ( .D(n1537), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X2 \mem_reg[13][7]  ( .D(n1536), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X2 \mem_reg[13][6]  ( .D(n1535), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X2 \mem_reg[13][5]  ( .D(n1534), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X2 \mem_reg[13][4]  ( .D(n1533), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X2 \mem_reg[13][3]  ( .D(n1532), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X2 \mem_reg[13][2]  ( .D(n1531), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X2 \mem_reg[13][1]  ( .D(n1530), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X2 \mem_reg[13][0]  ( .D(n1529), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X2 \mem_reg[12][31]  ( .D(n1528), .CK(clk), .Q(\mem[12][31] ) );
  DFF_X2 \mem_reg[12][30]  ( .D(n1527), .CK(clk), .Q(\mem[12][30] ) );
  DFF_X2 \mem_reg[12][29]  ( .D(n1526), .CK(clk), .Q(\mem[12][29] ) );
  DFF_X2 \mem_reg[12][28]  ( .D(n1525), .CK(clk), .Q(\mem[12][28] ) );
  DFF_X2 \mem_reg[12][27]  ( .D(n1524), .CK(clk), .Q(\mem[12][27] ) );
  DFF_X2 \mem_reg[12][26]  ( .D(n1523), .CK(clk), .Q(\mem[12][26] ) );
  DFF_X2 \mem_reg[12][25]  ( .D(n1522), .CK(clk), .Q(\mem[12][25] ) );
  DFF_X2 \mem_reg[12][24]  ( .D(n1521), .CK(clk), .Q(\mem[12][24] ) );
  DFF_X2 \mem_reg[12][23]  ( .D(n1520), .CK(clk), .Q(\mem[12][23] ) );
  DFF_X2 \mem_reg[12][22]  ( .D(n1519), .CK(clk), .Q(\mem[12][22] ) );
  DFF_X2 \mem_reg[12][21]  ( .D(n1518), .CK(clk), .Q(\mem[12][21] ) );
  DFF_X2 \mem_reg[12][20]  ( .D(n1517), .CK(clk), .Q(\mem[12][20] ) );
  DFF_X2 \mem_reg[12][19]  ( .D(n1516), .CK(clk), .Q(\mem[12][19] ) );
  DFF_X2 \mem_reg[12][18]  ( .D(n1515), .CK(clk), .Q(\mem[12][18] ) );
  DFF_X2 \mem_reg[12][17]  ( .D(n1514), .CK(clk), .Q(\mem[12][17] ) );
  DFF_X2 \mem_reg[12][16]  ( .D(n1513), .CK(clk), .Q(\mem[12][16] ) );
  DFF_X2 \mem_reg[12][15]  ( .D(n1512), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X2 \mem_reg[12][14]  ( .D(n1511), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X2 \mem_reg[12][13]  ( .D(n1510), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X2 \mem_reg[12][12]  ( .D(n1509), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X2 \mem_reg[12][11]  ( .D(n1508), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X2 \mem_reg[12][10]  ( .D(n1507), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X2 \mem_reg[12][9]  ( .D(n1506), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X2 \mem_reg[12][8]  ( .D(n1505), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X2 \mem_reg[12][7]  ( .D(n1504), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X2 \mem_reg[12][6]  ( .D(n1503), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X2 \mem_reg[12][5]  ( .D(n1502), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X2 \mem_reg[12][4]  ( .D(n1501), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X2 \mem_reg[12][3]  ( .D(n1500), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X2 \mem_reg[12][2]  ( .D(n1499), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X2 \mem_reg[12][1]  ( .D(n1498), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X2 \mem_reg[12][0]  ( .D(n1497), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X2 \mem_reg[11][31]  ( .D(n1496), .CK(clk), .Q(\mem[11][31] ) );
  DFF_X2 \mem_reg[11][30]  ( .D(n1495), .CK(clk), .Q(\mem[11][30] ) );
  DFF_X2 \mem_reg[11][29]  ( .D(n1494), .CK(clk), .Q(\mem[11][29] ) );
  DFF_X2 \mem_reg[11][28]  ( .D(n1493), .CK(clk), .Q(\mem[11][28] ) );
  DFF_X2 \mem_reg[11][27]  ( .D(n1492), .CK(clk), .Q(\mem[11][27] ) );
  DFF_X2 \mem_reg[11][26]  ( .D(n1491), .CK(clk), .Q(\mem[11][26] ) );
  DFF_X2 \mem_reg[11][25]  ( .D(n1490), .CK(clk), .Q(\mem[11][25] ) );
  DFF_X2 \mem_reg[11][24]  ( .D(n1489), .CK(clk), .Q(\mem[11][24] ) );
  DFF_X2 \mem_reg[11][23]  ( .D(n1488), .CK(clk), .Q(\mem[11][23] ) );
  DFF_X2 \mem_reg[11][22]  ( .D(n1487), .CK(clk), .Q(\mem[11][22] ) );
  DFF_X2 \mem_reg[11][21]  ( .D(n1486), .CK(clk), .Q(\mem[11][21] ) );
  DFF_X2 \mem_reg[11][20]  ( .D(n1485), .CK(clk), .Q(\mem[11][20] ) );
  DFF_X2 \mem_reg[11][19]  ( .D(n1484), .CK(clk), .Q(\mem[11][19] ) );
  DFF_X2 \mem_reg[11][18]  ( .D(n1483), .CK(clk), .Q(\mem[11][18] ) );
  DFF_X2 \mem_reg[11][17]  ( .D(n1482), .CK(clk), .Q(\mem[11][17] ) );
  DFF_X2 \mem_reg[11][16]  ( .D(n1481), .CK(clk), .Q(\mem[11][16] ) );
  DFF_X2 \mem_reg[11][15]  ( .D(n1480), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X2 \mem_reg[11][14]  ( .D(n1479), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X2 \mem_reg[11][13]  ( .D(n1478), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X2 \mem_reg[11][12]  ( .D(n1477), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X2 \mem_reg[11][11]  ( .D(n1476), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X2 \mem_reg[11][10]  ( .D(n1475), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X2 \mem_reg[11][9]  ( .D(n1474), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X2 \mem_reg[11][8]  ( .D(n1473), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X2 \mem_reg[11][7]  ( .D(n1472), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X2 \mem_reg[11][6]  ( .D(n1471), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X2 \mem_reg[11][5]  ( .D(n1470), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X2 \mem_reg[11][4]  ( .D(n1469), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X2 \mem_reg[11][3]  ( .D(n1468), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X2 \mem_reg[11][2]  ( .D(n1467), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X2 \mem_reg[11][1]  ( .D(n1466), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X2 \mem_reg[11][0]  ( .D(n1465), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X2 \mem_reg[10][31]  ( .D(n1464), .CK(clk), .Q(\mem[10][31] ) );
  DFF_X2 \mem_reg[10][30]  ( .D(n1463), .CK(clk), .Q(\mem[10][30] ) );
  DFF_X2 \mem_reg[10][29]  ( .D(n1462), .CK(clk), .Q(\mem[10][29] ) );
  DFF_X2 \mem_reg[10][28]  ( .D(n1461), .CK(clk), .Q(\mem[10][28] ) );
  DFF_X2 \mem_reg[10][27]  ( .D(n1460), .CK(clk), .Q(\mem[10][27] ) );
  DFF_X2 \mem_reg[10][26]  ( .D(n1459), .CK(clk), .Q(\mem[10][26] ) );
  DFF_X2 \mem_reg[10][25]  ( .D(n1458), .CK(clk), .Q(\mem[10][25] ) );
  DFF_X2 \mem_reg[10][24]  ( .D(n1457), .CK(clk), .Q(\mem[10][24] ) );
  DFF_X2 \mem_reg[10][23]  ( .D(n1456), .CK(clk), .Q(\mem[10][23] ) );
  DFF_X2 \mem_reg[10][22]  ( .D(n1455), .CK(clk), .Q(\mem[10][22] ) );
  DFF_X2 \mem_reg[10][21]  ( .D(n1454), .CK(clk), .Q(\mem[10][21] ) );
  DFF_X2 \mem_reg[10][20]  ( .D(n1453), .CK(clk), .Q(\mem[10][20] ) );
  DFF_X2 \mem_reg[10][19]  ( .D(n1452), .CK(clk), .Q(\mem[10][19] ) );
  DFF_X2 \mem_reg[10][18]  ( .D(n1451), .CK(clk), .Q(\mem[10][18] ) );
  DFF_X2 \mem_reg[10][17]  ( .D(n1450), .CK(clk), .Q(\mem[10][17] ) );
  DFF_X2 \mem_reg[10][16]  ( .D(n1449), .CK(clk), .Q(\mem[10][16] ) );
  DFF_X2 \mem_reg[10][15]  ( .D(n1448), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X2 \mem_reg[10][14]  ( .D(n1447), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X2 \mem_reg[10][13]  ( .D(n1446), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X2 \mem_reg[10][12]  ( .D(n1445), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X2 \mem_reg[10][11]  ( .D(n1444), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X2 \mem_reg[10][10]  ( .D(n1443), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X2 \mem_reg[10][9]  ( .D(n1442), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X2 \mem_reg[10][8]  ( .D(n1441), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X2 \mem_reg[10][7]  ( .D(n1440), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X2 \mem_reg[10][6]  ( .D(n1439), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X2 \mem_reg[10][5]  ( .D(n1438), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X2 \mem_reg[10][4]  ( .D(n1437), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X2 \mem_reg[10][3]  ( .D(n1436), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X2 \mem_reg[10][2]  ( .D(n1435), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X2 \mem_reg[10][1]  ( .D(n1434), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X2 \mem_reg[10][0]  ( .D(n1433), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X2 \mem_reg[9][31]  ( .D(n1432), .CK(clk), .Q(\mem[9][31] ) );
  DFF_X2 \mem_reg[9][30]  ( .D(n1431), .CK(clk), .Q(\mem[9][30] ) );
  DFF_X2 \mem_reg[9][29]  ( .D(n1430), .CK(clk), .Q(\mem[9][29] ) );
  DFF_X2 \mem_reg[9][28]  ( .D(n1429), .CK(clk), .Q(\mem[9][28] ) );
  DFF_X2 \mem_reg[9][27]  ( .D(n1428), .CK(clk), .Q(\mem[9][27] ) );
  DFF_X2 \mem_reg[9][26]  ( .D(n1427), .CK(clk), .Q(\mem[9][26] ) );
  DFF_X2 \mem_reg[9][25]  ( .D(n1426), .CK(clk), .Q(\mem[9][25] ) );
  DFF_X2 \mem_reg[9][24]  ( .D(n1425), .CK(clk), .Q(\mem[9][24] ) );
  DFF_X2 \mem_reg[9][23]  ( .D(n1424), .CK(clk), .Q(\mem[9][23] ) );
  DFF_X2 \mem_reg[9][22]  ( .D(n1423), .CK(clk), .Q(\mem[9][22] ) );
  DFF_X2 \mem_reg[9][21]  ( .D(n1422), .CK(clk), .Q(\mem[9][21] ) );
  DFF_X2 \mem_reg[9][20]  ( .D(n1421), .CK(clk), .Q(\mem[9][20] ) );
  DFF_X2 \mem_reg[9][19]  ( .D(n1420), .CK(clk), .Q(\mem[9][19] ) );
  DFF_X2 \mem_reg[9][18]  ( .D(n1419), .CK(clk), .Q(\mem[9][18] ) );
  DFF_X2 \mem_reg[9][17]  ( .D(n1418), .CK(clk), .Q(\mem[9][17] ) );
  DFF_X2 \mem_reg[9][16]  ( .D(n1417), .CK(clk), .Q(\mem[9][16] ) );
  DFF_X2 \mem_reg[9][15]  ( .D(n1416), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X2 \mem_reg[9][14]  ( .D(n1415), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X2 \mem_reg[9][13]  ( .D(n1414), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X2 \mem_reg[9][12]  ( .D(n1413), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X2 \mem_reg[9][11]  ( .D(n1412), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X2 \mem_reg[9][10]  ( .D(n1411), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X2 \mem_reg[9][9]  ( .D(n1410), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X2 \mem_reg[9][8]  ( .D(n1409), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X2 \mem_reg[9][7]  ( .D(n1408), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X2 \mem_reg[9][6]  ( .D(n1407), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X2 \mem_reg[9][5]  ( .D(n1406), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X2 \mem_reg[9][4]  ( .D(n1405), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X2 \mem_reg[9][3]  ( .D(n1404), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X2 \mem_reg[9][2]  ( .D(n1403), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X2 \mem_reg[9][1]  ( .D(n1402), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X2 \mem_reg[9][0]  ( .D(n1401), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X2 \mem_reg[8][31]  ( .D(n1400), .CK(clk), .Q(\mem[8][31] ) );
  DFF_X2 \mem_reg[8][30]  ( .D(n1399), .CK(clk), .Q(\mem[8][30] ) );
  DFF_X2 \mem_reg[8][29]  ( .D(n1398), .CK(clk), .Q(\mem[8][29] ) );
  DFF_X2 \mem_reg[8][28]  ( .D(n1397), .CK(clk), .Q(\mem[8][28] ) );
  DFF_X2 \mem_reg[8][27]  ( .D(n1396), .CK(clk), .Q(\mem[8][27] ) );
  DFF_X2 \mem_reg[8][26]  ( .D(n1395), .CK(clk), .Q(\mem[8][26] ) );
  DFF_X2 \mem_reg[8][25]  ( .D(n1394), .CK(clk), .Q(\mem[8][25] ) );
  DFF_X2 \mem_reg[8][24]  ( .D(n1393), .CK(clk), .Q(\mem[8][24] ) );
  DFF_X2 \mem_reg[8][23]  ( .D(n1392), .CK(clk), .Q(\mem[8][23] ) );
  DFF_X2 \mem_reg[8][22]  ( .D(n1391), .CK(clk), .Q(\mem[8][22] ) );
  DFF_X2 \mem_reg[8][21]  ( .D(n1390), .CK(clk), .Q(\mem[8][21] ) );
  DFF_X2 \mem_reg[8][20]  ( .D(n1389), .CK(clk), .Q(\mem[8][20] ) );
  DFF_X2 \mem_reg[8][19]  ( .D(n1388), .CK(clk), .Q(\mem[8][19] ) );
  DFF_X2 \mem_reg[8][18]  ( .D(n1387), .CK(clk), .Q(\mem[8][18] ) );
  DFF_X2 \mem_reg[8][17]  ( .D(n1386), .CK(clk), .Q(\mem[8][17] ) );
  DFF_X2 \mem_reg[8][16]  ( .D(n1385), .CK(clk), .Q(\mem[8][16] ) );
  DFF_X2 \mem_reg[8][15]  ( .D(n1384), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X2 \mem_reg[8][14]  ( .D(n1383), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X2 \mem_reg[8][13]  ( .D(n1382), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X2 \mem_reg[8][12]  ( .D(n1381), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X2 \mem_reg[8][11]  ( .D(n1380), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X2 \mem_reg[8][10]  ( .D(n1379), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X2 \mem_reg[8][9]  ( .D(n1378), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X2 \mem_reg[8][8]  ( .D(n1377), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X2 \mem_reg[8][7]  ( .D(n1376), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X2 \mem_reg[8][6]  ( .D(n1375), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X2 \mem_reg[8][5]  ( .D(n1374), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X2 \mem_reg[8][4]  ( .D(n1373), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X2 \mem_reg[8][3]  ( .D(n1372), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X2 \mem_reg[8][2]  ( .D(n1371), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X2 \mem_reg[8][1]  ( .D(n1370), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X2 \mem_reg[8][0]  ( .D(n1369), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X2 \mem_reg[7][31]  ( .D(n1368), .CK(clk), .Q(\mem[7][31] ) );
  DFF_X2 \mem_reg[7][30]  ( .D(n1367), .CK(clk), .Q(\mem[7][30] ) );
  DFF_X2 \mem_reg[7][29]  ( .D(n1366), .CK(clk), .Q(\mem[7][29] ) );
  DFF_X2 \mem_reg[7][28]  ( .D(n1365), .CK(clk), .Q(\mem[7][28] ) );
  DFF_X2 \mem_reg[7][27]  ( .D(n1364), .CK(clk), .Q(\mem[7][27] ) );
  DFF_X2 \mem_reg[7][26]  ( .D(n1363), .CK(clk), .Q(\mem[7][26] ) );
  DFF_X2 \mem_reg[7][25]  ( .D(n1362), .CK(clk), .Q(\mem[7][25] ) );
  DFF_X2 \mem_reg[7][24]  ( .D(n1361), .CK(clk), .Q(\mem[7][24] ) );
  DFF_X2 \mem_reg[7][23]  ( .D(n1360), .CK(clk), .Q(\mem[7][23] ) );
  DFF_X2 \mem_reg[7][22]  ( .D(n1359), .CK(clk), .Q(\mem[7][22] ) );
  DFF_X2 \mem_reg[7][21]  ( .D(n1358), .CK(clk), .Q(\mem[7][21] ) );
  DFF_X2 \mem_reg[7][20]  ( .D(n1357), .CK(clk), .Q(\mem[7][20] ) );
  DFF_X2 \mem_reg[7][19]  ( .D(n1356), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X2 \mem_reg[7][18]  ( .D(n1355), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X2 \mem_reg[7][17]  ( .D(n1354), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X2 \mem_reg[7][16]  ( .D(n1353), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X2 \mem_reg[7][15]  ( .D(n1352), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X2 \mem_reg[7][14]  ( .D(n1351), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X2 \mem_reg[7][13]  ( .D(n1350), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X2 \mem_reg[7][12]  ( .D(n1349), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X2 \mem_reg[7][11]  ( .D(n1348), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X2 \mem_reg[7][10]  ( .D(n1347), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X2 \mem_reg[7][9]  ( .D(n1346), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X2 \mem_reg[7][8]  ( .D(n1345), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X2 \mem_reg[7][7]  ( .D(n1344), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X2 \mem_reg[7][6]  ( .D(n1343), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X2 \mem_reg[7][5]  ( .D(n1342), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X2 \mem_reg[7][4]  ( .D(n1341), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X2 \mem_reg[7][3]  ( .D(n1340), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X2 \mem_reg[7][2]  ( .D(n1339), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X2 \mem_reg[7][1]  ( .D(n1338), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X2 \mem_reg[7][0]  ( .D(n1337), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X2 \mem_reg[6][31]  ( .D(n1336), .CK(clk), .Q(\mem[6][31] ) );
  DFF_X2 \mem_reg[6][30]  ( .D(n1335), .CK(clk), .Q(\mem[6][30] ) );
  DFF_X2 \mem_reg[6][29]  ( .D(n1334), .CK(clk), .Q(\mem[6][29] ) );
  DFF_X2 \mem_reg[6][28]  ( .D(n1333), .CK(clk), .Q(\mem[6][28] ) );
  DFF_X2 \mem_reg[6][27]  ( .D(n1332), .CK(clk), .Q(\mem[6][27] ) );
  DFF_X2 \mem_reg[6][26]  ( .D(n1331), .CK(clk), .Q(\mem[6][26] ) );
  DFF_X2 \mem_reg[6][25]  ( .D(n1330), .CK(clk), .Q(\mem[6][25] ) );
  DFF_X2 \mem_reg[6][24]  ( .D(n1329), .CK(clk), .Q(\mem[6][24] ) );
  DFF_X2 \mem_reg[6][23]  ( .D(n1328), .CK(clk), .Q(\mem[6][23] ) );
  DFF_X2 \mem_reg[6][22]  ( .D(n1327), .CK(clk), .Q(\mem[6][22] ) );
  DFF_X2 \mem_reg[6][21]  ( .D(n1326), .CK(clk), .Q(\mem[6][21] ) );
  DFF_X2 \mem_reg[6][20]  ( .D(n1325), .CK(clk), .Q(\mem[6][20] ) );
  DFF_X2 \mem_reg[6][19]  ( .D(n1324), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X2 \mem_reg[6][18]  ( .D(n1323), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X2 \mem_reg[6][17]  ( .D(n1322), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X2 \mem_reg[6][16]  ( .D(n1321), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X2 \mem_reg[6][15]  ( .D(n1320), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X2 \mem_reg[6][14]  ( .D(n1319), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X2 \mem_reg[6][13]  ( .D(n1318), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X2 \mem_reg[6][12]  ( .D(n1317), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X2 \mem_reg[6][11]  ( .D(n1316), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X2 \mem_reg[6][10]  ( .D(n1315), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X2 \mem_reg[6][9]  ( .D(n1314), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X2 \mem_reg[6][8]  ( .D(n1313), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X2 \mem_reg[6][7]  ( .D(n1312), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X2 \mem_reg[6][6]  ( .D(n1311), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X2 \mem_reg[6][5]  ( .D(n1310), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X2 \mem_reg[6][4]  ( .D(n1309), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X2 \mem_reg[6][3]  ( .D(n1308), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X2 \mem_reg[6][2]  ( .D(n1307), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X2 \mem_reg[6][1]  ( .D(n1306), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X2 \mem_reg[6][0]  ( .D(n1305), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X2 \mem_reg[5][31]  ( .D(n1304), .CK(clk), .Q(\mem[5][31] ) );
  DFF_X2 \mem_reg[5][30]  ( .D(n1303), .CK(clk), .Q(\mem[5][30] ) );
  DFF_X2 \mem_reg[5][29]  ( .D(n1302), .CK(clk), .Q(\mem[5][29] ) );
  DFF_X2 \mem_reg[5][28]  ( .D(n1301), .CK(clk), .Q(\mem[5][28] ) );
  DFF_X2 \mem_reg[5][27]  ( .D(n1300), .CK(clk), .Q(\mem[5][27] ) );
  DFF_X2 \mem_reg[5][26]  ( .D(n1299), .CK(clk), .Q(\mem[5][26] ) );
  DFF_X2 \mem_reg[5][25]  ( .D(n1298), .CK(clk), .Q(\mem[5][25] ) );
  DFF_X2 \mem_reg[5][24]  ( .D(n1297), .CK(clk), .Q(\mem[5][24] ) );
  DFF_X2 \mem_reg[5][23]  ( .D(n1296), .CK(clk), .Q(\mem[5][23] ) );
  DFF_X2 \mem_reg[5][22]  ( .D(n1295), .CK(clk), .Q(\mem[5][22] ) );
  DFF_X2 \mem_reg[5][21]  ( .D(n1294), .CK(clk), .Q(\mem[5][21] ) );
  DFF_X2 \mem_reg[5][20]  ( .D(n1293), .CK(clk), .Q(\mem[5][20] ) );
  DFF_X2 \mem_reg[5][19]  ( .D(n1292), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X2 \mem_reg[5][18]  ( .D(n1291), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X2 \mem_reg[5][17]  ( .D(n1290), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X2 \mem_reg[5][16]  ( .D(n1289), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X2 \mem_reg[5][15]  ( .D(n1288), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X2 \mem_reg[5][14]  ( .D(n1287), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X2 \mem_reg[5][13]  ( .D(n1286), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X2 \mem_reg[5][12]  ( .D(n1285), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X2 \mem_reg[5][11]  ( .D(n1284), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X2 \mem_reg[5][10]  ( .D(n1283), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X2 \mem_reg[5][9]  ( .D(n1282), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X2 \mem_reg[5][8]  ( .D(n1281), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X2 \mem_reg[5][7]  ( .D(n1280), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X2 \mem_reg[5][6]  ( .D(n1279), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X2 \mem_reg[5][5]  ( .D(n1278), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X2 \mem_reg[5][4]  ( .D(n1277), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X2 \mem_reg[5][3]  ( .D(n1276), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X2 \mem_reg[5][2]  ( .D(n1275), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X2 \mem_reg[5][1]  ( .D(n1274), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X2 \mem_reg[5][0]  ( .D(n1273), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X2 \mem_reg[4][31]  ( .D(n1272), .CK(clk), .Q(\mem[4][31] ) );
  DFF_X2 \mem_reg[4][30]  ( .D(n1271), .CK(clk), .Q(\mem[4][30] ) );
  DFF_X2 \mem_reg[4][29]  ( .D(n1270), .CK(clk), .Q(\mem[4][29] ) );
  DFF_X2 \mem_reg[4][28]  ( .D(n1269), .CK(clk), .Q(\mem[4][28] ) );
  DFF_X2 \mem_reg[4][27]  ( .D(n1268), .CK(clk), .Q(\mem[4][27] ) );
  DFF_X2 \mem_reg[4][26]  ( .D(n1267), .CK(clk), .Q(\mem[4][26] ) );
  DFF_X2 \mem_reg[4][25]  ( .D(n1266), .CK(clk), .Q(\mem[4][25] ) );
  DFF_X2 \mem_reg[4][24]  ( .D(n1265), .CK(clk), .Q(\mem[4][24] ) );
  DFF_X2 \mem_reg[4][23]  ( .D(n1264), .CK(clk), .Q(\mem[4][23] ) );
  DFF_X2 \mem_reg[4][22]  ( .D(n1263), .CK(clk), .Q(\mem[4][22] ) );
  DFF_X2 \mem_reg[4][21]  ( .D(n1262), .CK(clk), .Q(\mem[4][21] ) );
  DFF_X2 \mem_reg[4][20]  ( .D(n1261), .CK(clk), .Q(\mem[4][20] ) );
  DFF_X2 \mem_reg[4][19]  ( .D(n1260), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X2 \mem_reg[4][18]  ( .D(n1259), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X2 \mem_reg[4][17]  ( .D(n1258), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X2 \mem_reg[4][16]  ( .D(n1257), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X2 \mem_reg[4][15]  ( .D(n1256), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X2 \mem_reg[4][14]  ( .D(n1255), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X2 \mem_reg[4][13]  ( .D(n1254), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X2 \mem_reg[4][12]  ( .D(n1253), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X2 \mem_reg[4][11]  ( .D(n1252), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X2 \mem_reg[4][10]  ( .D(n1251), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X2 \mem_reg[4][9]  ( .D(n1250), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X2 \mem_reg[4][8]  ( .D(n1249), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X2 \mem_reg[4][7]  ( .D(n1248), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X2 \mem_reg[4][6]  ( .D(n1247), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X2 \mem_reg[4][5]  ( .D(n1246), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X2 \mem_reg[4][4]  ( .D(n1245), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X2 \mem_reg[4][3]  ( .D(n1244), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X2 \mem_reg[4][2]  ( .D(n1243), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X2 \mem_reg[4][1]  ( .D(n1242), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X2 \mem_reg[4][0]  ( .D(n1241), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X2 \mem_reg[3][31]  ( .D(n1240), .CK(clk), .Q(\mem[3][31] ) );
  DFF_X2 \mem_reg[3][30]  ( .D(n1239), .CK(clk), .Q(\mem[3][30] ) );
  DFF_X2 \mem_reg[3][29]  ( .D(n1238), .CK(clk), .Q(\mem[3][29] ) );
  DFF_X2 \mem_reg[3][28]  ( .D(n1237), .CK(clk), .Q(\mem[3][28] ) );
  DFF_X2 \mem_reg[3][27]  ( .D(n1236), .CK(clk), .Q(\mem[3][27] ) );
  DFF_X2 \mem_reg[3][26]  ( .D(n1235), .CK(clk), .Q(\mem[3][26] ) );
  DFF_X2 \mem_reg[3][25]  ( .D(n1234), .CK(clk), .Q(\mem[3][25] ) );
  DFF_X2 \mem_reg[3][24]  ( .D(n1233), .CK(clk), .Q(\mem[3][24] ) );
  DFF_X2 \mem_reg[3][23]  ( .D(n1232), .CK(clk), .Q(\mem[3][23] ) );
  DFF_X2 \mem_reg[3][22]  ( .D(n1231), .CK(clk), .Q(\mem[3][22] ) );
  DFF_X2 \mem_reg[3][21]  ( .D(n1230), .CK(clk), .Q(\mem[3][21] ) );
  DFF_X2 \mem_reg[3][20]  ( .D(n1229), .CK(clk), .Q(\mem[3][20] ) );
  DFF_X2 \mem_reg[3][19]  ( .D(n1228), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X2 \mem_reg[3][18]  ( .D(n1227), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X2 \mem_reg[3][17]  ( .D(n1226), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X2 \mem_reg[3][16]  ( .D(n1225), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X2 \mem_reg[3][15]  ( .D(n1224), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X2 \mem_reg[3][14]  ( .D(n1223), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X2 \mem_reg[3][13]  ( .D(n1222), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X2 \mem_reg[3][12]  ( .D(n1221), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X2 \mem_reg[3][11]  ( .D(n1220), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X2 \mem_reg[3][10]  ( .D(n1219), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X2 \mem_reg[3][9]  ( .D(n1218), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X2 \mem_reg[3][8]  ( .D(n1217), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X2 \mem_reg[3][7]  ( .D(n1216), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X2 \mem_reg[3][6]  ( .D(n1215), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X2 \mem_reg[3][5]  ( .D(n1214), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X2 \mem_reg[3][4]  ( .D(n1213), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X2 \mem_reg[3][3]  ( .D(n1212), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X2 \mem_reg[3][2]  ( .D(n1211), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X2 \mem_reg[3][1]  ( .D(n1210), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X2 \mem_reg[3][0]  ( .D(n1209), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X2 \mem_reg[2][31]  ( .D(n1208), .CK(clk), .Q(\mem[2][31] ) );
  DFF_X2 \mem_reg[2][30]  ( .D(n1207), .CK(clk), .Q(\mem[2][30] ) );
  DFF_X2 \mem_reg[2][29]  ( .D(n1206), .CK(clk), .Q(\mem[2][29] ) );
  DFF_X2 \mem_reg[2][28]  ( .D(n1205), .CK(clk), .Q(\mem[2][28] ) );
  DFF_X2 \mem_reg[2][27]  ( .D(n1204), .CK(clk), .Q(\mem[2][27] ) );
  DFF_X2 \mem_reg[2][26]  ( .D(n1203), .CK(clk), .Q(\mem[2][26] ) );
  DFF_X2 \mem_reg[2][25]  ( .D(n1202), .CK(clk), .Q(\mem[2][25] ) );
  DFF_X2 \mem_reg[2][24]  ( .D(n1201), .CK(clk), .Q(\mem[2][24] ) );
  DFF_X2 \mem_reg[2][23]  ( .D(n1200), .CK(clk), .Q(\mem[2][23] ) );
  DFF_X2 \mem_reg[2][22]  ( .D(n1199), .CK(clk), .Q(\mem[2][22] ) );
  DFF_X2 \mem_reg[2][21]  ( .D(n1198), .CK(clk), .Q(\mem[2][21] ) );
  DFF_X2 \mem_reg[2][20]  ( .D(n1197), .CK(clk), .Q(\mem[2][20] ) );
  DFF_X2 \mem_reg[2][19]  ( .D(n1196), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X2 \mem_reg[2][18]  ( .D(n1195), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X2 \mem_reg[2][17]  ( .D(n1194), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X2 \mem_reg[2][16]  ( .D(n1193), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X2 \mem_reg[2][15]  ( .D(n1192), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X2 \mem_reg[2][14]  ( .D(n1191), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X2 \mem_reg[2][13]  ( .D(n1190), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X2 \mem_reg[2][12]  ( .D(n1189), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X2 \mem_reg[2][11]  ( .D(n1188), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X2 \mem_reg[2][10]  ( .D(n1187), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X2 \mem_reg[2][9]  ( .D(n1186), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X2 \mem_reg[2][8]  ( .D(n1185), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X2 \mem_reg[2][7]  ( .D(n1184), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X2 \mem_reg[2][6]  ( .D(n1183), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X2 \mem_reg[2][5]  ( .D(n1182), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X2 \mem_reg[2][4]  ( .D(n1181), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X2 \mem_reg[2][3]  ( .D(n1180), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X2 \mem_reg[2][2]  ( .D(n1179), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X2 \mem_reg[2][1]  ( .D(n1178), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X2 \mem_reg[2][0]  ( .D(n1177), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X2 \mem_reg[1][31]  ( .D(n1176), .CK(clk), .Q(\mem[1][31] ) );
  DFF_X2 \mem_reg[1][30]  ( .D(n1175), .CK(clk), .Q(\mem[1][30] ) );
  DFF_X2 \mem_reg[1][29]  ( .D(n1174), .CK(clk), .Q(\mem[1][29] ) );
  DFF_X2 \mem_reg[1][28]  ( .D(n1173), .CK(clk), .Q(\mem[1][28] ) );
  DFF_X2 \mem_reg[1][27]  ( .D(n1172), .CK(clk), .Q(\mem[1][27] ) );
  DFF_X2 \mem_reg[1][26]  ( .D(n1171), .CK(clk), .Q(\mem[1][26] ) );
  DFF_X2 \mem_reg[1][25]  ( .D(n1170), .CK(clk), .Q(\mem[1][25] ) );
  DFF_X2 \mem_reg[1][24]  ( .D(n1169), .CK(clk), .Q(\mem[1][24] ) );
  DFF_X2 \mem_reg[1][23]  ( .D(n1168), .CK(clk), .Q(\mem[1][23] ) );
  DFF_X2 \mem_reg[1][22]  ( .D(n1167), .CK(clk), .Q(\mem[1][22] ) );
  DFF_X2 \mem_reg[1][21]  ( .D(n1166), .CK(clk), .Q(\mem[1][21] ) );
  DFF_X2 \mem_reg[1][20]  ( .D(n1165), .CK(clk), .Q(\mem[1][20] ) );
  DFF_X2 \mem_reg[1][19]  ( .D(n1164), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X2 \mem_reg[1][18]  ( .D(n1163), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X2 \mem_reg[1][17]  ( .D(n1162), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X2 \mem_reg[1][16]  ( .D(n1161), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X2 \mem_reg[1][15]  ( .D(n1160), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X2 \mem_reg[1][14]  ( .D(n1159), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X2 \mem_reg[1][13]  ( .D(n1158), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X2 \mem_reg[1][12]  ( .D(n1157), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X2 \mem_reg[1][11]  ( .D(n1156), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X2 \mem_reg[1][10]  ( .D(n1155), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X2 \mem_reg[1][9]  ( .D(n1154), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X2 \mem_reg[1][8]  ( .D(n1153), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X2 \mem_reg[1][7]  ( .D(n1152), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X2 \mem_reg[1][6]  ( .D(n1151), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X2 \mem_reg[1][5]  ( .D(n1150), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X2 \mem_reg[1][4]  ( .D(n1149), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X2 \mem_reg[1][3]  ( .D(n1148), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X2 \mem_reg[1][2]  ( .D(n1147), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X2 \mem_reg[1][1]  ( .D(n1146), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X2 \mem_reg[1][0]  ( .D(n1145), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X2 \mem_reg[0][31]  ( .D(n1144), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X2 \mem_reg[0][30]  ( .D(n1143), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X2 \mem_reg[0][29]  ( .D(n1142), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X2 \mem_reg[0][28]  ( .D(n1141), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X2 \mem_reg[0][27]  ( .D(n1140), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X2 \mem_reg[0][26]  ( .D(n1139), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X2 \mem_reg[0][25]  ( .D(n1138), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X2 \mem_reg[0][24]  ( .D(n1137), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X2 \mem_reg[0][23]  ( .D(n1136), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X2 \mem_reg[0][22]  ( .D(n1135), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X2 \mem_reg[0][21]  ( .D(n1134), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X2 \mem_reg[0][20]  ( .D(n1133), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X2 \mem_reg[0][19]  ( .D(n1132), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X2 \mem_reg[0][18]  ( .D(n1131), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X2 \mem_reg[0][17]  ( .D(n1130), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X2 \mem_reg[0][16]  ( .D(n1129), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X2 \mem_reg[0][15]  ( .D(n1128), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X2 \mem_reg[0][14]  ( .D(n1127), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X2 \mem_reg[0][13]  ( .D(n1126), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X2 \mem_reg[0][12]  ( .D(n1125), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X2 \mem_reg[0][11]  ( .D(n1124), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X2 \mem_reg[0][10]  ( .D(n1123), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X2 \mem_reg[0][9]  ( .D(n1122), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X2 \mem_reg[0][8]  ( .D(n1121), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X2 \mem_reg[0][7]  ( .D(n1120), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X2 \mem_reg[0][6]  ( .D(n1119), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X2 \mem_reg[0][5]  ( .D(n1118), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X2 \mem_reg[0][4]  ( .D(n1117), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X2 \mem_reg[0][3]  ( .D(n1116), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X2 \mem_reg[0][2]  ( .D(n1115), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X2 \mem_reg[0][1]  ( .D(n1114), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X2 \mem_reg[0][0]  ( .D(n1113), .CK(clk), .Q(\mem[0][0] ) );
  NAND2_X2 U3 ( .A1(\mem[9][9] ), .A2(n3380), .ZN(n3) );
  NAND2_X2 U5 ( .A1(\mem[9][8] ), .A2(n3379), .ZN(n5) );
  NAND2_X2 U7 ( .A1(\mem[9][7] ), .A2(n3380), .ZN(n7) );
  NAND2_X2 U9 ( .A1(\mem[9][6] ), .A2(n3379), .ZN(n9) );
  NAND2_X2 U11 ( .A1(\mem[9][5] ), .A2(n3380), .ZN(n11) );
  NAND2_X2 U13 ( .A1(\mem[9][4] ), .A2(n3379), .ZN(n13) );
  NAND2_X2 U15 ( .A1(\mem[9][3] ), .A2(n3380), .ZN(n15) );
  NAND2_X2 U17 ( .A1(\mem[9][31] ), .A2(n3381), .ZN(n17) );
  NAND2_X2 U19 ( .A1(\mem[9][30] ), .A2(n3381), .ZN(n19) );
  NAND2_X2 U21 ( .A1(\mem[9][2] ), .A2(n3381), .ZN(n21) );
  NAND2_X2 U23 ( .A1(\mem[9][29] ), .A2(n3381), .ZN(n23) );
  NAND2_X2 U25 ( .A1(\mem[9][28] ), .A2(n3381), .ZN(n25) );
  NAND2_X2 U27 ( .A1(\mem[9][27] ), .A2(n3381), .ZN(n27) );
  NAND2_X2 U29 ( .A1(\mem[9][26] ), .A2(n3381), .ZN(n29) );
  NAND2_X2 U31 ( .A1(\mem[9][25] ), .A2(n3381), .ZN(n31) );
  NAND2_X2 U33 ( .A1(\mem[9][24] ), .A2(n3381), .ZN(n33) );
  NAND2_X2 U35 ( .A1(\mem[9][23] ), .A2(n3381), .ZN(n35) );
  NAND2_X2 U37 ( .A1(\mem[9][22] ), .A2(n3381), .ZN(n37) );
  NAND2_X2 U39 ( .A1(\mem[9][21] ), .A2(n3381), .ZN(n39) );
  NAND2_X2 U41 ( .A1(\mem[9][20] ), .A2(n3381), .ZN(n41) );
  NAND2_X2 U43 ( .A1(\mem[9][1] ), .A2(n3381), .ZN(n43) );
  NAND2_X2 U45 ( .A1(\mem[9][19] ), .A2(n3381), .ZN(n45) );
  NAND2_X2 U47 ( .A1(\mem[9][18] ), .A2(n3381), .ZN(n47) );
  NAND2_X2 U49 ( .A1(\mem[9][17] ), .A2(n3381), .ZN(n49) );
  NAND2_X2 U51 ( .A1(\mem[9][16] ), .A2(n3381), .ZN(n51) );
  NAND2_X2 U53 ( .A1(\mem[9][15] ), .A2(n3381), .ZN(n53) );
  NAND2_X2 U55 ( .A1(\mem[9][14] ), .A2(n3381), .ZN(n55) );
  NAND2_X2 U57 ( .A1(\mem[9][13] ), .A2(n3381), .ZN(n57) );
  NAND2_X2 U59 ( .A1(\mem[9][12] ), .A2(n3381), .ZN(n59) );
  NAND2_X2 U61 ( .A1(\mem[9][11] ), .A2(n3381), .ZN(n61) );
  NAND2_X2 U63 ( .A1(\mem[9][10] ), .A2(n3381), .ZN(n63) );
  NAND2_X2 U65 ( .A1(\mem[9][0] ), .A2(n3381), .ZN(n65) );
  NAND2_X2 U66 ( .A1(n66), .A2(n67), .ZN(n1) );
  NAND2_X2 U68 ( .A1(\mem[8][9] ), .A2(n3376), .ZN(n69) );
  NAND2_X2 U70 ( .A1(\mem[8][8] ), .A2(n3375), .ZN(n70) );
  NAND2_X2 U72 ( .A1(\mem[8][7] ), .A2(n3376), .ZN(n71) );
  NAND2_X2 U74 ( .A1(\mem[8][6] ), .A2(n3375), .ZN(n72) );
  NAND2_X2 U76 ( .A1(\mem[8][5] ), .A2(n3376), .ZN(n73) );
  NAND2_X2 U78 ( .A1(\mem[8][4] ), .A2(n3375), .ZN(n74) );
  NAND2_X2 U80 ( .A1(\mem[8][3] ), .A2(n3376), .ZN(n75) );
  NAND2_X2 U82 ( .A1(\mem[8][31] ), .A2(n3377), .ZN(n76) );
  NAND2_X2 U84 ( .A1(\mem[8][30] ), .A2(n3377), .ZN(n77) );
  NAND2_X2 U86 ( .A1(\mem[8][2] ), .A2(n3377), .ZN(n78) );
  NAND2_X2 U88 ( .A1(\mem[8][29] ), .A2(n3377), .ZN(n79) );
  NAND2_X2 U90 ( .A1(\mem[8][28] ), .A2(n3377), .ZN(n80) );
  NAND2_X2 U92 ( .A1(\mem[8][27] ), .A2(n3377), .ZN(n81) );
  NAND2_X2 U94 ( .A1(\mem[8][26] ), .A2(n3377), .ZN(n82) );
  NAND2_X2 U96 ( .A1(\mem[8][25] ), .A2(n3377), .ZN(n83) );
  NAND2_X2 U98 ( .A1(\mem[8][24] ), .A2(n3377), .ZN(n84) );
  NAND2_X2 U100 ( .A1(\mem[8][23] ), .A2(n3377), .ZN(n85) );
  NAND2_X2 U102 ( .A1(\mem[8][22] ), .A2(n3377), .ZN(n86) );
  NAND2_X2 U104 ( .A1(\mem[8][21] ), .A2(n3377), .ZN(n87) );
  NAND2_X2 U106 ( .A1(\mem[8][20] ), .A2(n3377), .ZN(n88) );
  NAND2_X2 U108 ( .A1(\mem[8][1] ), .A2(n3377), .ZN(n89) );
  NAND2_X2 U110 ( .A1(\mem[8][19] ), .A2(n3377), .ZN(n90) );
  NAND2_X2 U112 ( .A1(\mem[8][18] ), .A2(n3377), .ZN(n91) );
  NAND2_X2 U114 ( .A1(\mem[8][17] ), .A2(n3377), .ZN(n92) );
  NAND2_X2 U116 ( .A1(\mem[8][16] ), .A2(n3377), .ZN(n93) );
  NAND2_X2 U118 ( .A1(\mem[8][15] ), .A2(n3377), .ZN(n94) );
  NAND2_X2 U120 ( .A1(\mem[8][14] ), .A2(n3377), .ZN(n95) );
  NAND2_X2 U122 ( .A1(\mem[8][13] ), .A2(n3377), .ZN(n96) );
  NAND2_X2 U124 ( .A1(\mem[8][12] ), .A2(n3377), .ZN(n97) );
  NAND2_X2 U126 ( .A1(\mem[8][11] ), .A2(n3377), .ZN(n98) );
  NAND2_X2 U128 ( .A1(\mem[8][10] ), .A2(n3377), .ZN(n99) );
  NAND2_X2 U130 ( .A1(\mem[8][0] ), .A2(n3377), .ZN(n100) );
  NAND2_X2 U131 ( .A1(n101), .A2(n67), .ZN(n68) );
  NAND2_X2 U133 ( .A1(\mem[7][9] ), .A2(n3372), .ZN(n103) );
  NAND2_X2 U135 ( .A1(\mem[7][8] ), .A2(n3371), .ZN(n104) );
  NAND2_X2 U137 ( .A1(\mem[7][7] ), .A2(n3372), .ZN(n105) );
  NAND2_X2 U139 ( .A1(\mem[7][6] ), .A2(n3371), .ZN(n106) );
  NAND2_X2 U141 ( .A1(\mem[7][5] ), .A2(n3372), .ZN(n107) );
  NAND2_X2 U143 ( .A1(\mem[7][4] ), .A2(n3371), .ZN(n108) );
  NAND2_X2 U145 ( .A1(\mem[7][3] ), .A2(n3372), .ZN(n109) );
  NAND2_X2 U147 ( .A1(\mem[7][31] ), .A2(n3373), .ZN(n110) );
  NAND2_X2 U149 ( .A1(\mem[7][30] ), .A2(n3373), .ZN(n111) );
  NAND2_X2 U151 ( .A1(\mem[7][2] ), .A2(n3373), .ZN(n112) );
  NAND2_X2 U153 ( .A1(\mem[7][29] ), .A2(n3373), .ZN(n113) );
  NAND2_X2 U155 ( .A1(\mem[7][28] ), .A2(n3373), .ZN(n114) );
  NAND2_X2 U157 ( .A1(\mem[7][27] ), .A2(n3373), .ZN(n115) );
  NAND2_X2 U159 ( .A1(\mem[7][26] ), .A2(n3373), .ZN(n116) );
  NAND2_X2 U161 ( .A1(\mem[7][25] ), .A2(n3373), .ZN(n117) );
  NAND2_X2 U163 ( .A1(\mem[7][24] ), .A2(n3373), .ZN(n118) );
  NAND2_X2 U165 ( .A1(\mem[7][23] ), .A2(n3373), .ZN(n119) );
  NAND2_X2 U167 ( .A1(\mem[7][22] ), .A2(n3373), .ZN(n120) );
  NAND2_X2 U169 ( .A1(\mem[7][21] ), .A2(n3373), .ZN(n121) );
  NAND2_X2 U171 ( .A1(\mem[7][20] ), .A2(n3373), .ZN(n122) );
  NAND2_X2 U173 ( .A1(\mem[7][1] ), .A2(n3373), .ZN(n123) );
  NAND2_X2 U175 ( .A1(\mem[7][19] ), .A2(n3373), .ZN(n124) );
  NAND2_X2 U177 ( .A1(\mem[7][18] ), .A2(n3373), .ZN(n125) );
  NAND2_X2 U179 ( .A1(\mem[7][17] ), .A2(n3373), .ZN(n126) );
  NAND2_X2 U181 ( .A1(\mem[7][16] ), .A2(n3373), .ZN(n127) );
  NAND2_X2 U183 ( .A1(\mem[7][15] ), .A2(n3373), .ZN(n128) );
  NAND2_X2 U185 ( .A1(\mem[7][14] ), .A2(n3373), .ZN(n129) );
  NAND2_X2 U187 ( .A1(\mem[7][13] ), .A2(n3373), .ZN(n130) );
  NAND2_X2 U189 ( .A1(\mem[7][12] ), .A2(n3373), .ZN(n131) );
  NAND2_X2 U191 ( .A1(\mem[7][11] ), .A2(n3373), .ZN(n132) );
  NAND2_X2 U193 ( .A1(\mem[7][10] ), .A2(n3373), .ZN(n133) );
  NAND2_X2 U195 ( .A1(\mem[7][0] ), .A2(n3373), .ZN(n134) );
  NAND2_X2 U196 ( .A1(n135), .A2(n136), .ZN(n102) );
  NAND2_X2 U198 ( .A1(\mem[6][9] ), .A2(n3368), .ZN(n138) );
  NAND2_X2 U200 ( .A1(\mem[6][8] ), .A2(n3367), .ZN(n139) );
  NAND2_X2 U202 ( .A1(\mem[6][7] ), .A2(n3368), .ZN(n140) );
  NAND2_X2 U204 ( .A1(\mem[6][6] ), .A2(n3367), .ZN(n141) );
  NAND2_X2 U206 ( .A1(\mem[6][5] ), .A2(n3368), .ZN(n142) );
  NAND2_X2 U208 ( .A1(\mem[6][4] ), .A2(n3367), .ZN(n143) );
  NAND2_X2 U210 ( .A1(\mem[6][3] ), .A2(n3368), .ZN(n144) );
  NAND2_X2 U212 ( .A1(\mem[6][31] ), .A2(n3369), .ZN(n145) );
  NAND2_X2 U214 ( .A1(\mem[6][30] ), .A2(n3369), .ZN(n146) );
  NAND2_X2 U216 ( .A1(\mem[6][2] ), .A2(n3369), .ZN(n147) );
  NAND2_X2 U218 ( .A1(\mem[6][29] ), .A2(n3369), .ZN(n148) );
  NAND2_X2 U220 ( .A1(\mem[6][28] ), .A2(n3369), .ZN(n149) );
  NAND2_X2 U222 ( .A1(\mem[6][27] ), .A2(n3369), .ZN(n150) );
  NAND2_X2 U224 ( .A1(\mem[6][26] ), .A2(n3369), .ZN(n151) );
  NAND2_X2 U226 ( .A1(\mem[6][25] ), .A2(n3369), .ZN(n152) );
  NAND2_X2 U228 ( .A1(\mem[6][24] ), .A2(n3369), .ZN(n153) );
  NAND2_X2 U230 ( .A1(\mem[6][23] ), .A2(n3369), .ZN(n154) );
  NAND2_X2 U232 ( .A1(\mem[6][22] ), .A2(n3369), .ZN(n155) );
  NAND2_X2 U234 ( .A1(\mem[6][21] ), .A2(n3369), .ZN(n156) );
  NAND2_X2 U236 ( .A1(\mem[6][20] ), .A2(n3369), .ZN(n157) );
  NAND2_X2 U238 ( .A1(\mem[6][1] ), .A2(n3369), .ZN(n158) );
  NAND2_X2 U240 ( .A1(\mem[6][19] ), .A2(n3369), .ZN(n159) );
  NAND2_X2 U242 ( .A1(\mem[6][18] ), .A2(n3369), .ZN(n160) );
  NAND2_X2 U244 ( .A1(\mem[6][17] ), .A2(n3369), .ZN(n161) );
  NAND2_X2 U246 ( .A1(\mem[6][16] ), .A2(n3369), .ZN(n162) );
  NAND2_X2 U248 ( .A1(\mem[6][15] ), .A2(n3369), .ZN(n163) );
  NAND2_X2 U250 ( .A1(\mem[6][14] ), .A2(n3369), .ZN(n164) );
  NAND2_X2 U252 ( .A1(\mem[6][13] ), .A2(n3369), .ZN(n165) );
  NAND2_X2 U254 ( .A1(\mem[6][12] ), .A2(n3369), .ZN(n166) );
  NAND2_X2 U256 ( .A1(\mem[6][11] ), .A2(n3369), .ZN(n167) );
  NAND2_X2 U258 ( .A1(\mem[6][10] ), .A2(n3369), .ZN(n168) );
  NAND2_X2 U260 ( .A1(\mem[6][0] ), .A2(n3369), .ZN(n169) );
  NAND2_X2 U261 ( .A1(n170), .A2(n136), .ZN(n137) );
  NAND2_X2 U263 ( .A1(\mem[5][9] ), .A2(n3364), .ZN(n172) );
  NAND2_X2 U265 ( .A1(\mem[5][8] ), .A2(n3362), .ZN(n173) );
  NAND2_X2 U267 ( .A1(\mem[5][7] ), .A2(n3363), .ZN(n174) );
  NAND2_X2 U269 ( .A1(\mem[5][6] ), .A2(n3362), .ZN(n175) );
  NAND2_X2 U271 ( .A1(\mem[5][5] ), .A2(n3363), .ZN(n176) );
  NAND2_X2 U273 ( .A1(\mem[5][4] ), .A2(n3362), .ZN(n177) );
  NAND2_X2 U275 ( .A1(\mem[5][3] ), .A2(n3363), .ZN(n178) );
  NAND2_X2 U277 ( .A1(\mem[5][31] ), .A2(n3364), .ZN(n179) );
  NAND2_X2 U279 ( .A1(\mem[5][30] ), .A2(n3364), .ZN(n180) );
  NAND2_X2 U281 ( .A1(\mem[5][2] ), .A2(n3364), .ZN(n181) );
  NAND2_X2 U283 ( .A1(\mem[5][29] ), .A2(n3364), .ZN(n182) );
  NAND2_X2 U285 ( .A1(\mem[5][28] ), .A2(n3364), .ZN(n183) );
  NAND2_X2 U287 ( .A1(\mem[5][27] ), .A2(n3364), .ZN(n184) );
  NAND2_X2 U289 ( .A1(\mem[5][26] ), .A2(n3364), .ZN(n185) );
  NAND2_X2 U291 ( .A1(\mem[5][25] ), .A2(n3364), .ZN(n186) );
  NAND2_X2 U293 ( .A1(\mem[5][24] ), .A2(n3364), .ZN(n187) );
  NAND2_X2 U295 ( .A1(\mem[5][23] ), .A2(n3364), .ZN(n188) );
  NAND2_X2 U297 ( .A1(\mem[5][22] ), .A2(n3364), .ZN(n189) );
  NAND2_X2 U299 ( .A1(\mem[5][21] ), .A2(n3364), .ZN(n190) );
  NAND2_X2 U301 ( .A1(\mem[5][20] ), .A2(n3364), .ZN(n191) );
  NAND2_X2 U303 ( .A1(\mem[5][1] ), .A2(n3364), .ZN(n192) );
  NAND2_X2 U305 ( .A1(\mem[5][19] ), .A2(n3364), .ZN(n193) );
  NAND2_X2 U307 ( .A1(\mem[5][18] ), .A2(n3364), .ZN(n194) );
  NAND2_X2 U309 ( .A1(\mem[5][17] ), .A2(n3364), .ZN(n195) );
  NAND2_X2 U311 ( .A1(\mem[5][16] ), .A2(n3364), .ZN(n196) );
  NAND2_X2 U313 ( .A1(\mem[5][15] ), .A2(n3364), .ZN(n197) );
  NAND2_X2 U315 ( .A1(\mem[5][14] ), .A2(n3364), .ZN(n198) );
  NAND2_X2 U317 ( .A1(\mem[5][13] ), .A2(n3364), .ZN(n199) );
  NAND2_X2 U319 ( .A1(\mem[5][12] ), .A2(n3363), .ZN(n200) );
  NAND2_X2 U321 ( .A1(\mem[5][11] ), .A2(n3364), .ZN(n201) );
  NAND2_X2 U323 ( .A1(\mem[5][10] ), .A2(n3362), .ZN(n202) );
  NAND2_X2 U325 ( .A1(\mem[5][0] ), .A2(n3364), .ZN(n203) );
  NAND2_X2 U326 ( .A1(n136), .A2(n66), .ZN(n171) );
  NAND2_X2 U328 ( .A1(\mem[4][9] ), .A2(n3360), .ZN(n205) );
  NAND2_X2 U330 ( .A1(\mem[4][8] ), .A2(n3358), .ZN(n206) );
  NAND2_X2 U332 ( .A1(\mem[4][7] ), .A2(n3359), .ZN(n207) );
  NAND2_X2 U334 ( .A1(\mem[4][6] ), .A2(n3358), .ZN(n208) );
  NAND2_X2 U336 ( .A1(\mem[4][5] ), .A2(n3359), .ZN(n209) );
  NAND2_X2 U338 ( .A1(\mem[4][4] ), .A2(n3358), .ZN(n210) );
  NAND2_X2 U340 ( .A1(\mem[4][3] ), .A2(n3359), .ZN(n211) );
  NAND2_X2 U342 ( .A1(\mem[4][31] ), .A2(n3360), .ZN(n212) );
  NAND2_X2 U344 ( .A1(\mem[4][30] ), .A2(n3360), .ZN(n213) );
  NAND2_X2 U346 ( .A1(\mem[4][2] ), .A2(n3360), .ZN(n214) );
  NAND2_X2 U348 ( .A1(\mem[4][29] ), .A2(n3360), .ZN(n215) );
  NAND2_X2 U350 ( .A1(\mem[4][28] ), .A2(n3360), .ZN(n216) );
  NAND2_X2 U352 ( .A1(\mem[4][27] ), .A2(n3360), .ZN(n217) );
  NAND2_X2 U354 ( .A1(\mem[4][26] ), .A2(n3360), .ZN(n218) );
  NAND2_X2 U356 ( .A1(\mem[4][25] ), .A2(n3360), .ZN(n219) );
  NAND2_X2 U358 ( .A1(\mem[4][24] ), .A2(n3360), .ZN(n220) );
  NAND2_X2 U360 ( .A1(\mem[4][23] ), .A2(n3360), .ZN(n221) );
  NAND2_X2 U362 ( .A1(\mem[4][22] ), .A2(n3360), .ZN(n222) );
  NAND2_X2 U364 ( .A1(\mem[4][21] ), .A2(n3360), .ZN(n223) );
  NAND2_X2 U366 ( .A1(\mem[4][20] ), .A2(n3360), .ZN(n224) );
  NAND2_X2 U368 ( .A1(\mem[4][1] ), .A2(n3360), .ZN(n225) );
  NAND2_X2 U370 ( .A1(\mem[4][19] ), .A2(n3360), .ZN(n226) );
  NAND2_X2 U372 ( .A1(\mem[4][18] ), .A2(n3360), .ZN(n227) );
  NAND2_X2 U374 ( .A1(\mem[4][17] ), .A2(n3360), .ZN(n228) );
  NAND2_X2 U376 ( .A1(\mem[4][16] ), .A2(n3360), .ZN(n229) );
  NAND2_X2 U378 ( .A1(\mem[4][15] ), .A2(n3360), .ZN(n230) );
  NAND2_X2 U380 ( .A1(\mem[4][14] ), .A2(n3360), .ZN(n231) );
  NAND2_X2 U382 ( .A1(\mem[4][13] ), .A2(n3360), .ZN(n232) );
  NAND2_X2 U384 ( .A1(\mem[4][12] ), .A2(n3359), .ZN(n233) );
  NAND2_X2 U386 ( .A1(\mem[4][11] ), .A2(n3360), .ZN(n234) );
  NAND2_X2 U388 ( .A1(\mem[4][10] ), .A2(n3358), .ZN(n235) );
  NAND2_X2 U390 ( .A1(\mem[4][0] ), .A2(n3360), .ZN(n236) );
  NAND2_X2 U391 ( .A1(n136), .A2(n101), .ZN(n204) );
  AND2_X2 U392 ( .A1(n237), .A2(n238), .ZN(n136) );
  NAND2_X2 U394 ( .A1(\mem[3][9] ), .A2(n3356), .ZN(n240) );
  NAND2_X2 U396 ( .A1(\mem[3][8] ), .A2(n3355), .ZN(n241) );
  NAND2_X2 U398 ( .A1(\mem[3][7] ), .A2(n3356), .ZN(n242) );
  NAND2_X2 U400 ( .A1(\mem[3][6] ), .A2(n3355), .ZN(n243) );
  NAND2_X2 U402 ( .A1(\mem[3][5] ), .A2(n3356), .ZN(n244) );
  NAND2_X2 U404 ( .A1(\mem[3][4] ), .A2(n3355), .ZN(n245) );
  NAND2_X2 U406 ( .A1(\mem[3][3] ), .A2(n3356), .ZN(n246) );
  NAND2_X2 U408 ( .A1(\mem[3][31] ), .A2(n3357), .ZN(n247) );
  NAND2_X2 U410 ( .A1(\mem[3][30] ), .A2(n3357), .ZN(n248) );
  NAND2_X2 U412 ( .A1(\mem[3][2] ), .A2(n3357), .ZN(n249) );
  NAND2_X2 U414 ( .A1(\mem[3][29] ), .A2(n3357), .ZN(n250) );
  NAND2_X2 U416 ( .A1(\mem[3][28] ), .A2(n3357), .ZN(n251) );
  NAND2_X2 U418 ( .A1(\mem[3][27] ), .A2(n3357), .ZN(n252) );
  NAND2_X2 U420 ( .A1(\mem[3][26] ), .A2(n3357), .ZN(n253) );
  NAND2_X2 U422 ( .A1(\mem[3][25] ), .A2(n3357), .ZN(n254) );
  NAND2_X2 U424 ( .A1(\mem[3][24] ), .A2(n3357), .ZN(n255) );
  NAND2_X2 U426 ( .A1(\mem[3][23] ), .A2(n3357), .ZN(n256) );
  NAND2_X2 U428 ( .A1(\mem[3][22] ), .A2(n3357), .ZN(n257) );
  NAND2_X2 U430 ( .A1(\mem[3][21] ), .A2(n3357), .ZN(n258) );
  NAND2_X2 U432 ( .A1(\mem[3][20] ), .A2(n3357), .ZN(n259) );
  NAND2_X2 U434 ( .A1(\mem[3][1] ), .A2(n3357), .ZN(n260) );
  NAND2_X2 U436 ( .A1(\mem[3][19] ), .A2(n3357), .ZN(n261) );
  NAND2_X2 U438 ( .A1(\mem[3][18] ), .A2(n3357), .ZN(n262) );
  NAND2_X2 U440 ( .A1(\mem[3][17] ), .A2(n3357), .ZN(n263) );
  NAND2_X2 U442 ( .A1(\mem[3][16] ), .A2(n3357), .ZN(n264) );
  NAND2_X2 U444 ( .A1(\mem[3][15] ), .A2(n3357), .ZN(n265) );
  NAND2_X2 U446 ( .A1(\mem[3][14] ), .A2(n3357), .ZN(n266) );
  NAND2_X2 U448 ( .A1(\mem[3][13] ), .A2(n3357), .ZN(n267) );
  NAND2_X2 U450 ( .A1(\mem[3][12] ), .A2(n3357), .ZN(n268) );
  NAND2_X2 U452 ( .A1(\mem[3][11] ), .A2(n3357), .ZN(n269) );
  NAND2_X2 U454 ( .A1(\mem[3][10] ), .A2(n3357), .ZN(n270) );
  NAND2_X2 U456 ( .A1(\mem[3][0] ), .A2(n3357), .ZN(n271) );
  NAND2_X2 U457 ( .A1(n272), .A2(n135), .ZN(n239) );
  NAND2_X2 U459 ( .A1(\mem[31][9] ), .A2(n3352), .ZN(n274) );
  NAND2_X2 U461 ( .A1(\mem[31][8] ), .A2(n3351), .ZN(n275) );
  NAND2_X2 U463 ( .A1(\mem[31][7] ), .A2(n3352), .ZN(n276) );
  NAND2_X2 U465 ( .A1(\mem[31][6] ), .A2(n3351), .ZN(n277) );
  NAND2_X2 U467 ( .A1(\mem[31][5] ), .A2(n3352), .ZN(n278) );
  NAND2_X2 U469 ( .A1(\mem[31][4] ), .A2(n3351), .ZN(n279) );
  NAND2_X2 U471 ( .A1(\mem[31][3] ), .A2(n3352), .ZN(n280) );
  NAND2_X2 U473 ( .A1(\mem[31][31] ), .A2(n3353), .ZN(n281) );
  NAND2_X2 U475 ( .A1(\mem[31][30] ), .A2(n3353), .ZN(n282) );
  NAND2_X2 U477 ( .A1(\mem[31][2] ), .A2(n3353), .ZN(n283) );
  NAND2_X2 U479 ( .A1(\mem[31][29] ), .A2(n3353), .ZN(n284) );
  NAND2_X2 U481 ( .A1(\mem[31][28] ), .A2(n3353), .ZN(n285) );
  NAND2_X2 U483 ( .A1(\mem[31][27] ), .A2(n3353), .ZN(n286) );
  NAND2_X2 U485 ( .A1(\mem[31][26] ), .A2(n3353), .ZN(n287) );
  NAND2_X2 U487 ( .A1(\mem[31][25] ), .A2(n3353), .ZN(n288) );
  NAND2_X2 U489 ( .A1(\mem[31][24] ), .A2(n3353), .ZN(n289) );
  NAND2_X2 U491 ( .A1(\mem[31][23] ), .A2(n3353), .ZN(n290) );
  NAND2_X2 U493 ( .A1(\mem[31][22] ), .A2(n3353), .ZN(n291) );
  NAND2_X2 U495 ( .A1(\mem[31][21] ), .A2(n3353), .ZN(n292) );
  NAND2_X2 U497 ( .A1(\mem[31][20] ), .A2(n3353), .ZN(n293) );
  NAND2_X2 U499 ( .A1(\mem[31][1] ), .A2(n3353), .ZN(n294) );
  NAND2_X2 U501 ( .A1(\mem[31][19] ), .A2(n3353), .ZN(n295) );
  NAND2_X2 U503 ( .A1(\mem[31][18] ), .A2(n3353), .ZN(n296) );
  NAND2_X2 U505 ( .A1(\mem[31][17] ), .A2(n3353), .ZN(n297) );
  NAND2_X2 U507 ( .A1(\mem[31][16] ), .A2(n3353), .ZN(n298) );
  NAND2_X2 U509 ( .A1(\mem[31][15] ), .A2(n3353), .ZN(n299) );
  NAND2_X2 U511 ( .A1(\mem[31][14] ), .A2(n3353), .ZN(n300) );
  NAND2_X2 U513 ( .A1(\mem[31][13] ), .A2(n3353), .ZN(n301) );
  NAND2_X2 U515 ( .A1(\mem[31][12] ), .A2(n3353), .ZN(n302) );
  NAND2_X2 U517 ( .A1(\mem[31][11] ), .A2(n3353), .ZN(n303) );
  NAND2_X2 U519 ( .A1(\mem[31][10] ), .A2(n3353), .ZN(n304) );
  NAND2_X2 U521 ( .A1(\mem[31][0] ), .A2(n3353), .ZN(n305) );
  NAND2_X2 U522 ( .A1(n306), .A2(n135), .ZN(n273) );
  NAND2_X2 U524 ( .A1(\mem[30][9] ), .A2(n3348), .ZN(n308) );
  NAND2_X2 U526 ( .A1(\mem[30][8] ), .A2(n3347), .ZN(n309) );
  NAND2_X2 U528 ( .A1(\mem[30][7] ), .A2(n3348), .ZN(n310) );
  NAND2_X2 U530 ( .A1(\mem[30][6] ), .A2(n3347), .ZN(n311) );
  NAND2_X2 U532 ( .A1(\mem[30][5] ), .A2(n3348), .ZN(n312) );
  NAND2_X2 U534 ( .A1(\mem[30][4] ), .A2(n3347), .ZN(n313) );
  NAND2_X2 U536 ( .A1(\mem[30][3] ), .A2(n3348), .ZN(n314) );
  NAND2_X2 U538 ( .A1(\mem[30][31] ), .A2(n3349), .ZN(n315) );
  NAND2_X2 U540 ( .A1(\mem[30][30] ), .A2(n3349), .ZN(n316) );
  NAND2_X2 U542 ( .A1(\mem[30][2] ), .A2(n3349), .ZN(n317) );
  NAND2_X2 U544 ( .A1(\mem[30][29] ), .A2(n3349), .ZN(n318) );
  NAND2_X2 U546 ( .A1(\mem[30][28] ), .A2(n3349), .ZN(n319) );
  NAND2_X2 U548 ( .A1(\mem[30][27] ), .A2(n3349), .ZN(n320) );
  NAND2_X2 U550 ( .A1(\mem[30][26] ), .A2(n3349), .ZN(n321) );
  NAND2_X2 U552 ( .A1(\mem[30][25] ), .A2(n3349), .ZN(n322) );
  NAND2_X2 U554 ( .A1(\mem[30][24] ), .A2(n3349), .ZN(n323) );
  NAND2_X2 U556 ( .A1(\mem[30][23] ), .A2(n3349), .ZN(n324) );
  NAND2_X2 U558 ( .A1(\mem[30][22] ), .A2(n3349), .ZN(n325) );
  NAND2_X2 U560 ( .A1(\mem[30][21] ), .A2(n3349), .ZN(n326) );
  NAND2_X2 U562 ( .A1(\mem[30][20] ), .A2(n3349), .ZN(n327) );
  NAND2_X2 U564 ( .A1(\mem[30][1] ), .A2(n3349), .ZN(n328) );
  NAND2_X2 U566 ( .A1(\mem[30][19] ), .A2(n3349), .ZN(n329) );
  NAND2_X2 U568 ( .A1(\mem[30][18] ), .A2(n3349), .ZN(n330) );
  NAND2_X2 U570 ( .A1(\mem[30][17] ), .A2(n3349), .ZN(n331) );
  NAND2_X2 U572 ( .A1(\mem[30][16] ), .A2(n3349), .ZN(n332) );
  NAND2_X2 U574 ( .A1(\mem[30][15] ), .A2(n3349), .ZN(n333) );
  NAND2_X2 U576 ( .A1(\mem[30][14] ), .A2(n3349), .ZN(n334) );
  NAND2_X2 U578 ( .A1(\mem[30][13] ), .A2(n3349), .ZN(n335) );
  NAND2_X2 U580 ( .A1(\mem[30][12] ), .A2(n3349), .ZN(n336) );
  NAND2_X2 U582 ( .A1(\mem[30][11] ), .A2(n3349), .ZN(n337) );
  NAND2_X2 U584 ( .A1(\mem[30][10] ), .A2(n3349), .ZN(n338) );
  NAND2_X2 U586 ( .A1(\mem[30][0] ), .A2(n3349), .ZN(n339) );
  NAND2_X2 U587 ( .A1(n306), .A2(n170), .ZN(n307) );
  NAND2_X2 U589 ( .A1(\mem[2][9] ), .A2(n3344), .ZN(n341) );
  NAND2_X2 U591 ( .A1(\mem[2][8] ), .A2(n3343), .ZN(n342) );
  NAND2_X2 U593 ( .A1(\mem[2][7] ), .A2(n3344), .ZN(n343) );
  NAND2_X2 U595 ( .A1(\mem[2][6] ), .A2(n3343), .ZN(n344) );
  NAND2_X2 U597 ( .A1(\mem[2][5] ), .A2(n3344), .ZN(n345) );
  NAND2_X2 U599 ( .A1(\mem[2][4] ), .A2(n3343), .ZN(n346) );
  NAND2_X2 U601 ( .A1(\mem[2][3] ), .A2(n3344), .ZN(n347) );
  NAND2_X2 U603 ( .A1(\mem[2][31] ), .A2(n3345), .ZN(n348) );
  NAND2_X2 U605 ( .A1(\mem[2][30] ), .A2(n3345), .ZN(n349) );
  NAND2_X2 U607 ( .A1(\mem[2][2] ), .A2(n3345), .ZN(n350) );
  NAND2_X2 U609 ( .A1(\mem[2][29] ), .A2(n3345), .ZN(n351) );
  NAND2_X2 U611 ( .A1(\mem[2][28] ), .A2(n3345), .ZN(n352) );
  NAND2_X2 U613 ( .A1(\mem[2][27] ), .A2(n3345), .ZN(n353) );
  NAND2_X2 U615 ( .A1(\mem[2][26] ), .A2(n3345), .ZN(n354) );
  NAND2_X2 U617 ( .A1(\mem[2][25] ), .A2(n3345), .ZN(n355) );
  NAND2_X2 U619 ( .A1(\mem[2][24] ), .A2(n3345), .ZN(n356) );
  NAND2_X2 U621 ( .A1(\mem[2][23] ), .A2(n3345), .ZN(n357) );
  NAND2_X2 U623 ( .A1(\mem[2][22] ), .A2(n3345), .ZN(n358) );
  NAND2_X2 U625 ( .A1(\mem[2][21] ), .A2(n3345), .ZN(n359) );
  NAND2_X2 U627 ( .A1(\mem[2][20] ), .A2(n3345), .ZN(n360) );
  NAND2_X2 U629 ( .A1(\mem[2][1] ), .A2(n3345), .ZN(n361) );
  NAND2_X2 U631 ( .A1(\mem[2][19] ), .A2(n3345), .ZN(n362) );
  NAND2_X2 U633 ( .A1(\mem[2][18] ), .A2(n3345), .ZN(n363) );
  NAND2_X2 U635 ( .A1(\mem[2][17] ), .A2(n3345), .ZN(n364) );
  NAND2_X2 U637 ( .A1(\mem[2][16] ), .A2(n3345), .ZN(n365) );
  NAND2_X2 U639 ( .A1(\mem[2][15] ), .A2(n3345), .ZN(n366) );
  NAND2_X2 U641 ( .A1(\mem[2][14] ), .A2(n3345), .ZN(n367) );
  NAND2_X2 U643 ( .A1(\mem[2][13] ), .A2(n3345), .ZN(n368) );
  NAND2_X2 U645 ( .A1(\mem[2][12] ), .A2(n3345), .ZN(n369) );
  NAND2_X2 U647 ( .A1(\mem[2][11] ), .A2(n3345), .ZN(n370) );
  NAND2_X2 U649 ( .A1(\mem[2][10] ), .A2(n3345), .ZN(n371) );
  NAND2_X2 U651 ( .A1(\mem[2][0] ), .A2(n3345), .ZN(n372) );
  NAND2_X2 U652 ( .A1(n272), .A2(n170), .ZN(n340) );
  NAND2_X2 U654 ( .A1(\mem[29][9] ), .A2(n3340), .ZN(n374) );
  NAND2_X2 U656 ( .A1(\mem[29][8] ), .A2(n3338), .ZN(n375) );
  NAND2_X2 U658 ( .A1(\mem[29][7] ), .A2(n3339), .ZN(n376) );
  NAND2_X2 U660 ( .A1(\mem[29][6] ), .A2(n3338), .ZN(n377) );
  NAND2_X2 U662 ( .A1(\mem[29][5] ), .A2(n3339), .ZN(n378) );
  NAND2_X2 U664 ( .A1(\mem[29][4] ), .A2(n3338), .ZN(n379) );
  NAND2_X2 U666 ( .A1(\mem[29][3] ), .A2(n3339), .ZN(n380) );
  NAND2_X2 U668 ( .A1(\mem[29][31] ), .A2(n3340), .ZN(n381) );
  NAND2_X2 U670 ( .A1(\mem[29][30] ), .A2(n3340), .ZN(n382) );
  NAND2_X2 U672 ( .A1(\mem[29][2] ), .A2(n3340), .ZN(n383) );
  NAND2_X2 U674 ( .A1(\mem[29][29] ), .A2(n3340), .ZN(n384) );
  NAND2_X2 U676 ( .A1(\mem[29][28] ), .A2(n3340), .ZN(n385) );
  NAND2_X2 U678 ( .A1(\mem[29][27] ), .A2(n3340), .ZN(n386) );
  NAND2_X2 U680 ( .A1(\mem[29][26] ), .A2(n3340), .ZN(n387) );
  NAND2_X2 U682 ( .A1(\mem[29][25] ), .A2(n3340), .ZN(n388) );
  NAND2_X2 U684 ( .A1(\mem[29][24] ), .A2(n3340), .ZN(n389) );
  NAND2_X2 U686 ( .A1(\mem[29][23] ), .A2(n3340), .ZN(n390) );
  NAND2_X2 U688 ( .A1(\mem[29][22] ), .A2(n3340), .ZN(n391) );
  NAND2_X2 U690 ( .A1(\mem[29][21] ), .A2(n3340), .ZN(n392) );
  NAND2_X2 U692 ( .A1(\mem[29][20] ), .A2(n3340), .ZN(n393) );
  NAND2_X2 U694 ( .A1(\mem[29][1] ), .A2(n3340), .ZN(n394) );
  NAND2_X2 U696 ( .A1(\mem[29][19] ), .A2(n3340), .ZN(n395) );
  NAND2_X2 U698 ( .A1(\mem[29][18] ), .A2(n3340), .ZN(n396) );
  NAND2_X2 U700 ( .A1(\mem[29][17] ), .A2(n3340), .ZN(n397) );
  NAND2_X2 U702 ( .A1(\mem[29][16] ), .A2(n3340), .ZN(n398) );
  NAND2_X2 U704 ( .A1(\mem[29][15] ), .A2(n3340), .ZN(n399) );
  NAND2_X2 U706 ( .A1(\mem[29][14] ), .A2(n3340), .ZN(n400) );
  NAND2_X2 U708 ( .A1(\mem[29][13] ), .A2(n3340), .ZN(n401) );
  NAND2_X2 U710 ( .A1(\mem[29][12] ), .A2(n3339), .ZN(n402) );
  NAND2_X2 U712 ( .A1(\mem[29][11] ), .A2(n3340), .ZN(n403) );
  NAND2_X2 U714 ( .A1(\mem[29][10] ), .A2(n3338), .ZN(n404) );
  NAND2_X2 U716 ( .A1(\mem[29][0] ), .A2(n3340), .ZN(n405) );
  NAND2_X2 U717 ( .A1(n306), .A2(n66), .ZN(n373) );
  NAND2_X2 U719 ( .A1(\mem[28][9] ), .A2(n3336), .ZN(n407) );
  NAND2_X2 U721 ( .A1(\mem[28][8] ), .A2(n3334), .ZN(n408) );
  NAND2_X2 U723 ( .A1(\mem[28][7] ), .A2(n3335), .ZN(n409) );
  NAND2_X2 U725 ( .A1(\mem[28][6] ), .A2(n3334), .ZN(n410) );
  NAND2_X2 U727 ( .A1(\mem[28][5] ), .A2(n3335), .ZN(n411) );
  NAND2_X2 U729 ( .A1(\mem[28][4] ), .A2(n3334), .ZN(n412) );
  NAND2_X2 U731 ( .A1(\mem[28][3] ), .A2(n3335), .ZN(n413) );
  NAND2_X2 U733 ( .A1(\mem[28][31] ), .A2(n3336), .ZN(n414) );
  NAND2_X2 U735 ( .A1(\mem[28][30] ), .A2(n3336), .ZN(n415) );
  NAND2_X2 U737 ( .A1(\mem[28][2] ), .A2(n3336), .ZN(n416) );
  NAND2_X2 U739 ( .A1(\mem[28][29] ), .A2(n3336), .ZN(n417) );
  NAND2_X2 U741 ( .A1(\mem[28][28] ), .A2(n3336), .ZN(n418) );
  NAND2_X2 U743 ( .A1(\mem[28][27] ), .A2(n3336), .ZN(n419) );
  NAND2_X2 U745 ( .A1(\mem[28][26] ), .A2(n3336), .ZN(n420) );
  NAND2_X2 U747 ( .A1(\mem[28][25] ), .A2(n3336), .ZN(n421) );
  NAND2_X2 U749 ( .A1(\mem[28][24] ), .A2(n3336), .ZN(n422) );
  NAND2_X2 U751 ( .A1(\mem[28][23] ), .A2(n3336), .ZN(n423) );
  NAND2_X2 U753 ( .A1(\mem[28][22] ), .A2(n3336), .ZN(n424) );
  NAND2_X2 U755 ( .A1(\mem[28][21] ), .A2(n3336), .ZN(n425) );
  NAND2_X2 U757 ( .A1(\mem[28][20] ), .A2(n3336), .ZN(n426) );
  NAND2_X2 U759 ( .A1(\mem[28][1] ), .A2(n3336), .ZN(n427) );
  NAND2_X2 U761 ( .A1(\mem[28][19] ), .A2(n3336), .ZN(n428) );
  NAND2_X2 U763 ( .A1(\mem[28][18] ), .A2(n3336), .ZN(n429) );
  NAND2_X2 U765 ( .A1(\mem[28][17] ), .A2(n3336), .ZN(n430) );
  NAND2_X2 U767 ( .A1(\mem[28][16] ), .A2(n3336), .ZN(n431) );
  NAND2_X2 U769 ( .A1(\mem[28][15] ), .A2(n3336), .ZN(n432) );
  NAND2_X2 U771 ( .A1(\mem[28][14] ), .A2(n3336), .ZN(n433) );
  NAND2_X2 U773 ( .A1(\mem[28][13] ), .A2(n3336), .ZN(n434) );
  NAND2_X2 U775 ( .A1(\mem[28][12] ), .A2(n3335), .ZN(n435) );
  NAND2_X2 U777 ( .A1(\mem[28][11] ), .A2(n3336), .ZN(n436) );
  NAND2_X2 U779 ( .A1(\mem[28][10] ), .A2(n3334), .ZN(n437) );
  NAND2_X2 U781 ( .A1(\mem[28][0] ), .A2(n3336), .ZN(n438) );
  NAND2_X2 U782 ( .A1(n306), .A2(n101), .ZN(n406) );
  AND2_X2 U783 ( .A1(n439), .A2(n440), .ZN(n306) );
  NAND2_X2 U785 ( .A1(\mem[27][9] ), .A2(n3332), .ZN(n442) );
  NAND2_X2 U787 ( .A1(\mem[27][8] ), .A2(n3331), .ZN(n443) );
  NAND2_X2 U789 ( .A1(\mem[27][7] ), .A2(n3332), .ZN(n444) );
  NAND2_X2 U791 ( .A1(\mem[27][6] ), .A2(n3331), .ZN(n445) );
  NAND2_X2 U793 ( .A1(\mem[27][5] ), .A2(n3332), .ZN(n446) );
  NAND2_X2 U795 ( .A1(\mem[27][4] ), .A2(n3331), .ZN(n447) );
  NAND2_X2 U797 ( .A1(\mem[27][3] ), .A2(n3332), .ZN(n448) );
  NAND2_X2 U799 ( .A1(\mem[27][31] ), .A2(n3333), .ZN(n449) );
  NAND2_X2 U801 ( .A1(\mem[27][30] ), .A2(n3333), .ZN(n450) );
  NAND2_X2 U803 ( .A1(\mem[27][2] ), .A2(n3333), .ZN(n451) );
  NAND2_X2 U805 ( .A1(\mem[27][29] ), .A2(n3333), .ZN(n452) );
  NAND2_X2 U807 ( .A1(\mem[27][28] ), .A2(n3333), .ZN(n453) );
  NAND2_X2 U809 ( .A1(\mem[27][27] ), .A2(n3333), .ZN(n454) );
  NAND2_X2 U811 ( .A1(\mem[27][26] ), .A2(n3333), .ZN(n455) );
  NAND2_X2 U813 ( .A1(\mem[27][25] ), .A2(n3333), .ZN(n456) );
  NAND2_X2 U815 ( .A1(\mem[27][24] ), .A2(n3333), .ZN(n457) );
  NAND2_X2 U817 ( .A1(\mem[27][23] ), .A2(n3333), .ZN(n458) );
  NAND2_X2 U819 ( .A1(\mem[27][22] ), .A2(n3333), .ZN(n459) );
  NAND2_X2 U821 ( .A1(\mem[27][21] ), .A2(n3333), .ZN(n460) );
  NAND2_X2 U823 ( .A1(\mem[27][20] ), .A2(n3333), .ZN(n461) );
  NAND2_X2 U825 ( .A1(\mem[27][1] ), .A2(n3333), .ZN(n462) );
  NAND2_X2 U827 ( .A1(\mem[27][19] ), .A2(n3333), .ZN(n463) );
  NAND2_X2 U829 ( .A1(\mem[27][18] ), .A2(n3333), .ZN(n464) );
  NAND2_X2 U831 ( .A1(\mem[27][17] ), .A2(n3333), .ZN(n465) );
  NAND2_X2 U833 ( .A1(\mem[27][16] ), .A2(n3333), .ZN(n466) );
  NAND2_X2 U835 ( .A1(\mem[27][15] ), .A2(n3333), .ZN(n467) );
  NAND2_X2 U837 ( .A1(\mem[27][14] ), .A2(n3333), .ZN(n468) );
  NAND2_X2 U839 ( .A1(\mem[27][13] ), .A2(n3333), .ZN(n469) );
  NAND2_X2 U841 ( .A1(\mem[27][12] ), .A2(n3333), .ZN(n470) );
  NAND2_X2 U843 ( .A1(\mem[27][11] ), .A2(n3333), .ZN(n471) );
  NAND2_X2 U845 ( .A1(\mem[27][10] ), .A2(n3333), .ZN(n472) );
  NAND2_X2 U847 ( .A1(\mem[27][0] ), .A2(n3333), .ZN(n473) );
  NAND2_X2 U848 ( .A1(n474), .A2(n135), .ZN(n441) );
  NAND2_X2 U850 ( .A1(\mem[26][9] ), .A2(n3328), .ZN(n476) );
  NAND2_X2 U852 ( .A1(\mem[26][8] ), .A2(n3327), .ZN(n477) );
  NAND2_X2 U854 ( .A1(\mem[26][7] ), .A2(n3328), .ZN(n478) );
  NAND2_X2 U856 ( .A1(\mem[26][6] ), .A2(n3327), .ZN(n479) );
  NAND2_X2 U858 ( .A1(\mem[26][5] ), .A2(n3328), .ZN(n480) );
  NAND2_X2 U860 ( .A1(\mem[26][4] ), .A2(n3327), .ZN(n481) );
  NAND2_X2 U862 ( .A1(\mem[26][3] ), .A2(n3328), .ZN(n482) );
  NAND2_X2 U864 ( .A1(\mem[26][31] ), .A2(n3329), .ZN(n483) );
  NAND2_X2 U866 ( .A1(\mem[26][30] ), .A2(n3329), .ZN(n484) );
  NAND2_X2 U868 ( .A1(\mem[26][2] ), .A2(n3329), .ZN(n485) );
  NAND2_X2 U870 ( .A1(\mem[26][29] ), .A2(n3329), .ZN(n486) );
  NAND2_X2 U872 ( .A1(\mem[26][28] ), .A2(n3329), .ZN(n487) );
  NAND2_X2 U874 ( .A1(\mem[26][27] ), .A2(n3329), .ZN(n488) );
  NAND2_X2 U876 ( .A1(\mem[26][26] ), .A2(n3329), .ZN(n489) );
  NAND2_X2 U878 ( .A1(\mem[26][25] ), .A2(n3329), .ZN(n490) );
  NAND2_X2 U880 ( .A1(\mem[26][24] ), .A2(n3329), .ZN(n491) );
  NAND2_X2 U882 ( .A1(\mem[26][23] ), .A2(n3329), .ZN(n492) );
  NAND2_X2 U884 ( .A1(\mem[26][22] ), .A2(n3329), .ZN(n493) );
  NAND2_X2 U886 ( .A1(\mem[26][21] ), .A2(n3329), .ZN(n494) );
  NAND2_X2 U888 ( .A1(\mem[26][20] ), .A2(n3329), .ZN(n495) );
  NAND2_X2 U890 ( .A1(\mem[26][1] ), .A2(n3329), .ZN(n496) );
  NAND2_X2 U892 ( .A1(\mem[26][19] ), .A2(n3329), .ZN(n497) );
  NAND2_X2 U894 ( .A1(\mem[26][18] ), .A2(n3329), .ZN(n498) );
  NAND2_X2 U896 ( .A1(\mem[26][17] ), .A2(n3329), .ZN(n499) );
  NAND2_X2 U898 ( .A1(\mem[26][16] ), .A2(n3329), .ZN(n500) );
  NAND2_X2 U900 ( .A1(\mem[26][15] ), .A2(n3329), .ZN(n501) );
  NAND2_X2 U902 ( .A1(\mem[26][14] ), .A2(n3329), .ZN(n502) );
  NAND2_X2 U904 ( .A1(\mem[26][13] ), .A2(n3329), .ZN(n503) );
  NAND2_X2 U906 ( .A1(\mem[26][12] ), .A2(n3329), .ZN(n504) );
  NAND2_X2 U908 ( .A1(\mem[26][11] ), .A2(n3329), .ZN(n505) );
  NAND2_X2 U910 ( .A1(\mem[26][10] ), .A2(n3329), .ZN(n506) );
  NAND2_X2 U912 ( .A1(\mem[26][0] ), .A2(n3329), .ZN(n507) );
  NAND2_X2 U913 ( .A1(n474), .A2(n170), .ZN(n475) );
  NAND2_X2 U915 ( .A1(\mem[25][9] ), .A2(n3324), .ZN(n509) );
  NAND2_X2 U917 ( .A1(\mem[25][8] ), .A2(n3322), .ZN(n510) );
  NAND2_X2 U919 ( .A1(\mem[25][7] ), .A2(n3323), .ZN(n511) );
  NAND2_X2 U921 ( .A1(\mem[25][6] ), .A2(n3322), .ZN(n512) );
  NAND2_X2 U923 ( .A1(\mem[25][5] ), .A2(n3323), .ZN(n513) );
  NAND2_X2 U925 ( .A1(\mem[25][4] ), .A2(n3322), .ZN(n514) );
  NAND2_X2 U927 ( .A1(\mem[25][3] ), .A2(n3323), .ZN(n515) );
  NAND2_X2 U929 ( .A1(\mem[25][31] ), .A2(n3324), .ZN(n516) );
  NAND2_X2 U931 ( .A1(\mem[25][30] ), .A2(n3324), .ZN(n517) );
  NAND2_X2 U933 ( .A1(\mem[25][2] ), .A2(n3324), .ZN(n518) );
  NAND2_X2 U935 ( .A1(\mem[25][29] ), .A2(n3324), .ZN(n519) );
  NAND2_X2 U937 ( .A1(\mem[25][28] ), .A2(n3324), .ZN(n520) );
  NAND2_X2 U939 ( .A1(\mem[25][27] ), .A2(n3324), .ZN(n521) );
  NAND2_X2 U941 ( .A1(\mem[25][26] ), .A2(n3324), .ZN(n522) );
  NAND2_X2 U943 ( .A1(\mem[25][25] ), .A2(n3324), .ZN(n523) );
  NAND2_X2 U945 ( .A1(\mem[25][24] ), .A2(n3324), .ZN(n524) );
  NAND2_X2 U947 ( .A1(\mem[25][23] ), .A2(n3324), .ZN(n525) );
  NAND2_X2 U949 ( .A1(\mem[25][22] ), .A2(n3324), .ZN(n526) );
  NAND2_X2 U951 ( .A1(\mem[25][21] ), .A2(n3324), .ZN(n527) );
  NAND2_X2 U953 ( .A1(\mem[25][20] ), .A2(n3324), .ZN(n528) );
  NAND2_X2 U955 ( .A1(\mem[25][1] ), .A2(n3324), .ZN(n529) );
  NAND2_X2 U957 ( .A1(\mem[25][19] ), .A2(n3324), .ZN(n530) );
  NAND2_X2 U959 ( .A1(\mem[25][18] ), .A2(n3324), .ZN(n531) );
  NAND2_X2 U961 ( .A1(\mem[25][17] ), .A2(n3324), .ZN(n532) );
  NAND2_X2 U963 ( .A1(\mem[25][16] ), .A2(n3324), .ZN(n533) );
  NAND2_X2 U965 ( .A1(\mem[25][15] ), .A2(n3324), .ZN(n534) );
  NAND2_X2 U967 ( .A1(\mem[25][14] ), .A2(n3324), .ZN(n535) );
  NAND2_X2 U969 ( .A1(\mem[25][13] ), .A2(n3324), .ZN(n536) );
  NAND2_X2 U971 ( .A1(\mem[25][12] ), .A2(n3323), .ZN(n537) );
  NAND2_X2 U973 ( .A1(\mem[25][11] ), .A2(n3324), .ZN(n538) );
  NAND2_X2 U975 ( .A1(\mem[25][10] ), .A2(n3322), .ZN(n539) );
  NAND2_X2 U977 ( .A1(\mem[25][0] ), .A2(n3324), .ZN(n540) );
  NAND2_X2 U978 ( .A1(n474), .A2(n66), .ZN(n508) );
  NAND2_X2 U980 ( .A1(\mem[24][9] ), .A2(n3320), .ZN(n542) );
  NAND2_X2 U982 ( .A1(\mem[24][8] ), .A2(n3318), .ZN(n543) );
  NAND2_X2 U984 ( .A1(\mem[24][7] ), .A2(n3319), .ZN(n544) );
  NAND2_X2 U986 ( .A1(\mem[24][6] ), .A2(n3318), .ZN(n545) );
  NAND2_X2 U988 ( .A1(\mem[24][5] ), .A2(n3319), .ZN(n546) );
  NAND2_X2 U990 ( .A1(\mem[24][4] ), .A2(n3318), .ZN(n547) );
  NAND2_X2 U992 ( .A1(\mem[24][3] ), .A2(n3319), .ZN(n548) );
  NAND2_X2 U994 ( .A1(\mem[24][31] ), .A2(n3320), .ZN(n549) );
  NAND2_X2 U996 ( .A1(\mem[24][30] ), .A2(n3320), .ZN(n550) );
  NAND2_X2 U998 ( .A1(\mem[24][2] ), .A2(n3320), .ZN(n551) );
  NAND2_X2 U1000 ( .A1(\mem[24][29] ), .A2(n3320), .ZN(n552) );
  NAND2_X2 U1002 ( .A1(\mem[24][28] ), .A2(n3320), .ZN(n553) );
  NAND2_X2 U1004 ( .A1(\mem[24][27] ), .A2(n3320), .ZN(n554) );
  NAND2_X2 U1006 ( .A1(\mem[24][26] ), .A2(n3320), .ZN(n555) );
  NAND2_X2 U1008 ( .A1(\mem[24][25] ), .A2(n3320), .ZN(n556) );
  NAND2_X2 U1010 ( .A1(\mem[24][24] ), .A2(n3320), .ZN(n557) );
  NAND2_X2 U1012 ( .A1(\mem[24][23] ), .A2(n3320), .ZN(n558) );
  NAND2_X2 U1014 ( .A1(\mem[24][22] ), .A2(n3320), .ZN(n559) );
  NAND2_X2 U1016 ( .A1(\mem[24][21] ), .A2(n3320), .ZN(n560) );
  NAND2_X2 U1018 ( .A1(\mem[24][20] ), .A2(n3320), .ZN(n561) );
  NAND2_X2 U1020 ( .A1(\mem[24][1] ), .A2(n3320), .ZN(n562) );
  NAND2_X2 U1022 ( .A1(\mem[24][19] ), .A2(n3320), .ZN(n563) );
  NAND2_X2 U1024 ( .A1(\mem[24][18] ), .A2(n3320), .ZN(n564) );
  NAND2_X2 U1026 ( .A1(\mem[24][17] ), .A2(n3320), .ZN(n565) );
  NAND2_X2 U1028 ( .A1(\mem[24][16] ), .A2(n3320), .ZN(n566) );
  NAND2_X2 U1030 ( .A1(\mem[24][15] ), .A2(n3320), .ZN(n567) );
  NAND2_X2 U1032 ( .A1(\mem[24][14] ), .A2(n3320), .ZN(n568) );
  NAND2_X2 U1034 ( .A1(\mem[24][13] ), .A2(n3320), .ZN(n569) );
  NAND2_X2 U1036 ( .A1(\mem[24][12] ), .A2(n3319), .ZN(n570) );
  NAND2_X2 U1038 ( .A1(\mem[24][11] ), .A2(n3320), .ZN(n571) );
  NAND2_X2 U1040 ( .A1(\mem[24][10] ), .A2(n3318), .ZN(n572) );
  NAND2_X2 U1042 ( .A1(\mem[24][0] ), .A2(n3320), .ZN(n573) );
  NAND2_X2 U1043 ( .A1(n474), .A2(n101), .ZN(n541) );
  AND2_X2 U1044 ( .A1(n439), .A2(n574), .ZN(n474) );
  NAND2_X2 U1046 ( .A1(\mem[23][9] ), .A2(n3316), .ZN(n576) );
  NAND2_X2 U1048 ( .A1(\mem[23][8] ), .A2(n3315), .ZN(n577) );
  NAND2_X2 U1050 ( .A1(\mem[23][7] ), .A2(n3316), .ZN(n578) );
  NAND2_X2 U1052 ( .A1(\mem[23][6] ), .A2(n3315), .ZN(n579) );
  NAND2_X2 U1054 ( .A1(\mem[23][5] ), .A2(n3316), .ZN(n580) );
  NAND2_X2 U1056 ( .A1(\mem[23][4] ), .A2(n3315), .ZN(n581) );
  NAND2_X2 U1058 ( .A1(\mem[23][3] ), .A2(n3316), .ZN(n582) );
  NAND2_X2 U1060 ( .A1(\mem[23][31] ), .A2(n3317), .ZN(n583) );
  NAND2_X2 U1062 ( .A1(\mem[23][30] ), .A2(n3317), .ZN(n584) );
  NAND2_X2 U1064 ( .A1(\mem[23][2] ), .A2(n3317), .ZN(n585) );
  NAND2_X2 U1066 ( .A1(\mem[23][29] ), .A2(n3317), .ZN(n586) );
  NAND2_X2 U1068 ( .A1(\mem[23][28] ), .A2(n3317), .ZN(n587) );
  NAND2_X2 U1070 ( .A1(\mem[23][27] ), .A2(n3317), .ZN(n588) );
  NAND2_X2 U1072 ( .A1(\mem[23][26] ), .A2(n3317), .ZN(n589) );
  NAND2_X2 U1074 ( .A1(\mem[23][25] ), .A2(n3317), .ZN(n590) );
  NAND2_X2 U1076 ( .A1(\mem[23][24] ), .A2(n3317), .ZN(n591) );
  NAND2_X2 U1078 ( .A1(\mem[23][23] ), .A2(n3317), .ZN(n592) );
  NAND2_X2 U1080 ( .A1(\mem[23][22] ), .A2(n3317), .ZN(n593) );
  NAND2_X2 U1082 ( .A1(\mem[23][21] ), .A2(n3317), .ZN(n594) );
  NAND2_X2 U1084 ( .A1(\mem[23][20] ), .A2(n3317), .ZN(n595) );
  NAND2_X2 U1086 ( .A1(\mem[23][1] ), .A2(n3317), .ZN(n596) );
  NAND2_X2 U1088 ( .A1(\mem[23][19] ), .A2(n3317), .ZN(n597) );
  NAND2_X2 U1090 ( .A1(\mem[23][18] ), .A2(n3317), .ZN(n598) );
  NAND2_X2 U1092 ( .A1(\mem[23][17] ), .A2(n3317), .ZN(n599) );
  NAND2_X2 U1094 ( .A1(\mem[23][16] ), .A2(n3317), .ZN(n600) );
  NAND2_X2 U1096 ( .A1(\mem[23][15] ), .A2(n3317), .ZN(n601) );
  NAND2_X2 U1098 ( .A1(\mem[23][14] ), .A2(n3317), .ZN(n602) );
  NAND2_X2 U1100 ( .A1(\mem[23][13] ), .A2(n3317), .ZN(n603) );
  NAND2_X2 U1102 ( .A1(\mem[23][12] ), .A2(n3317), .ZN(n604) );
  NAND2_X2 U1104 ( .A1(\mem[23][11] ), .A2(n3317), .ZN(n605) );
  NAND2_X2 U1106 ( .A1(\mem[23][10] ), .A2(n3317), .ZN(n606) );
  NAND2_X2 U1108 ( .A1(\mem[23][0] ), .A2(n3317), .ZN(n607) );
  NAND2_X2 U1109 ( .A1(n608), .A2(n135), .ZN(n575) );
  NAND2_X2 U1111 ( .A1(\mem[22][9] ), .A2(n3312), .ZN(n610) );
  NAND2_X2 U1113 ( .A1(\mem[22][8] ), .A2(n3311), .ZN(n611) );
  NAND2_X2 U1115 ( .A1(\mem[22][7] ), .A2(n3312), .ZN(n612) );
  NAND2_X2 U1117 ( .A1(\mem[22][6] ), .A2(n3311), .ZN(n613) );
  NAND2_X2 U1119 ( .A1(\mem[22][5] ), .A2(n3312), .ZN(n614) );
  NAND2_X2 U1121 ( .A1(\mem[22][4] ), .A2(n3311), .ZN(n615) );
  NAND2_X2 U1123 ( .A1(\mem[22][3] ), .A2(n3312), .ZN(n616) );
  NAND2_X2 U1125 ( .A1(\mem[22][31] ), .A2(n3313), .ZN(n617) );
  NAND2_X2 U1127 ( .A1(\mem[22][30] ), .A2(n3313), .ZN(n618) );
  NAND2_X2 U1129 ( .A1(\mem[22][2] ), .A2(n3313), .ZN(n619) );
  NAND2_X2 U1131 ( .A1(\mem[22][29] ), .A2(n3313), .ZN(n620) );
  NAND2_X2 U1133 ( .A1(\mem[22][28] ), .A2(n3313), .ZN(n621) );
  NAND2_X2 U1135 ( .A1(\mem[22][27] ), .A2(n3313), .ZN(n622) );
  NAND2_X2 U1137 ( .A1(\mem[22][26] ), .A2(n3313), .ZN(n623) );
  NAND2_X2 U1139 ( .A1(\mem[22][25] ), .A2(n3313), .ZN(n624) );
  NAND2_X2 U1141 ( .A1(\mem[22][24] ), .A2(n3313), .ZN(n625) );
  NAND2_X2 U1143 ( .A1(\mem[22][23] ), .A2(n3313), .ZN(n626) );
  NAND2_X2 U1145 ( .A1(\mem[22][22] ), .A2(n3313), .ZN(n627) );
  NAND2_X2 U1147 ( .A1(\mem[22][21] ), .A2(n3313), .ZN(n628) );
  NAND2_X2 U1149 ( .A1(\mem[22][20] ), .A2(n3313), .ZN(n629) );
  NAND2_X2 U1151 ( .A1(\mem[22][1] ), .A2(n3313), .ZN(n630) );
  NAND2_X2 U1153 ( .A1(\mem[22][19] ), .A2(n3313), .ZN(n631) );
  NAND2_X2 U1155 ( .A1(\mem[22][18] ), .A2(n3313), .ZN(n632) );
  NAND2_X2 U1157 ( .A1(\mem[22][17] ), .A2(n3313), .ZN(n633) );
  NAND2_X2 U1159 ( .A1(\mem[22][16] ), .A2(n3313), .ZN(n634) );
  NAND2_X2 U1161 ( .A1(\mem[22][15] ), .A2(n3313), .ZN(n635) );
  NAND2_X2 U1163 ( .A1(\mem[22][14] ), .A2(n3313), .ZN(n636) );
  NAND2_X2 U1165 ( .A1(\mem[22][13] ), .A2(n3313), .ZN(n637) );
  NAND2_X2 U1167 ( .A1(\mem[22][12] ), .A2(n3313), .ZN(n638) );
  NAND2_X2 U1169 ( .A1(\mem[22][11] ), .A2(n3313), .ZN(n639) );
  NAND2_X2 U1171 ( .A1(\mem[22][10] ), .A2(n3313), .ZN(n640) );
  NAND2_X2 U1173 ( .A1(\mem[22][0] ), .A2(n3313), .ZN(n641) );
  NAND2_X2 U1174 ( .A1(n608), .A2(n170), .ZN(n609) );
  NAND2_X2 U1176 ( .A1(\mem[21][9] ), .A2(n3308), .ZN(n643) );
  NAND2_X2 U1178 ( .A1(\mem[21][8] ), .A2(n3306), .ZN(n644) );
  NAND2_X2 U1180 ( .A1(\mem[21][7] ), .A2(n3307), .ZN(n645) );
  NAND2_X2 U1182 ( .A1(\mem[21][6] ), .A2(n3306), .ZN(n646) );
  NAND2_X2 U1184 ( .A1(\mem[21][5] ), .A2(n3307), .ZN(n647) );
  NAND2_X2 U1186 ( .A1(\mem[21][4] ), .A2(n3306), .ZN(n648) );
  NAND2_X2 U1188 ( .A1(\mem[21][3] ), .A2(n3307), .ZN(n649) );
  NAND2_X2 U1190 ( .A1(\mem[21][31] ), .A2(n3308), .ZN(n650) );
  NAND2_X2 U1192 ( .A1(\mem[21][30] ), .A2(n3308), .ZN(n651) );
  NAND2_X2 U1194 ( .A1(\mem[21][2] ), .A2(n3308), .ZN(n652) );
  NAND2_X2 U1196 ( .A1(\mem[21][29] ), .A2(n3308), .ZN(n653) );
  NAND2_X2 U1198 ( .A1(\mem[21][28] ), .A2(n3308), .ZN(n654) );
  NAND2_X2 U1200 ( .A1(\mem[21][27] ), .A2(n3308), .ZN(n655) );
  NAND2_X2 U1202 ( .A1(\mem[21][26] ), .A2(n3308), .ZN(n656) );
  NAND2_X2 U1204 ( .A1(\mem[21][25] ), .A2(n3308), .ZN(n657) );
  NAND2_X2 U1206 ( .A1(\mem[21][24] ), .A2(n3308), .ZN(n658) );
  NAND2_X2 U1208 ( .A1(\mem[21][23] ), .A2(n3308), .ZN(n659) );
  NAND2_X2 U1210 ( .A1(\mem[21][22] ), .A2(n3308), .ZN(n660) );
  NAND2_X2 U1212 ( .A1(\mem[21][21] ), .A2(n3308), .ZN(n661) );
  NAND2_X2 U1214 ( .A1(\mem[21][20] ), .A2(n3308), .ZN(n662) );
  NAND2_X2 U1216 ( .A1(\mem[21][1] ), .A2(n3308), .ZN(n663) );
  NAND2_X2 U1218 ( .A1(\mem[21][19] ), .A2(n3308), .ZN(n664) );
  NAND2_X2 U1220 ( .A1(\mem[21][18] ), .A2(n3308), .ZN(n665) );
  NAND2_X2 U1222 ( .A1(\mem[21][17] ), .A2(n3308), .ZN(n666) );
  NAND2_X2 U1224 ( .A1(\mem[21][16] ), .A2(n3308), .ZN(n667) );
  NAND2_X2 U1226 ( .A1(\mem[21][15] ), .A2(n3308), .ZN(n668) );
  NAND2_X2 U1228 ( .A1(\mem[21][14] ), .A2(n3308), .ZN(n669) );
  NAND2_X2 U1230 ( .A1(\mem[21][13] ), .A2(n3308), .ZN(n670) );
  NAND2_X2 U1232 ( .A1(\mem[21][12] ), .A2(n3307), .ZN(n671) );
  NAND2_X2 U1234 ( .A1(\mem[21][11] ), .A2(n3308), .ZN(n672) );
  NAND2_X2 U1236 ( .A1(\mem[21][10] ), .A2(n3306), .ZN(n673) );
  NAND2_X2 U1238 ( .A1(\mem[21][0] ), .A2(n3308), .ZN(n674) );
  NAND2_X2 U1239 ( .A1(n608), .A2(n66), .ZN(n642) );
  NAND2_X2 U1241 ( .A1(\mem[20][9] ), .A2(n3304), .ZN(n676) );
  NAND2_X2 U1243 ( .A1(\mem[20][8] ), .A2(n3302), .ZN(n677) );
  NAND2_X2 U1245 ( .A1(\mem[20][7] ), .A2(n3303), .ZN(n678) );
  NAND2_X2 U1247 ( .A1(\mem[20][6] ), .A2(n3302), .ZN(n679) );
  NAND2_X2 U1249 ( .A1(\mem[20][5] ), .A2(n3303), .ZN(n680) );
  NAND2_X2 U1251 ( .A1(\mem[20][4] ), .A2(n3302), .ZN(n681) );
  NAND2_X2 U1253 ( .A1(\mem[20][3] ), .A2(n3303), .ZN(n682) );
  NAND2_X2 U1255 ( .A1(\mem[20][31] ), .A2(n3304), .ZN(n683) );
  NAND2_X2 U1257 ( .A1(\mem[20][30] ), .A2(n3304), .ZN(n684) );
  NAND2_X2 U1259 ( .A1(\mem[20][2] ), .A2(n3304), .ZN(n685) );
  NAND2_X2 U1261 ( .A1(\mem[20][29] ), .A2(n3304), .ZN(n686) );
  NAND2_X2 U1263 ( .A1(\mem[20][28] ), .A2(n3304), .ZN(n687) );
  NAND2_X2 U1265 ( .A1(\mem[20][27] ), .A2(n3304), .ZN(n688) );
  NAND2_X2 U1267 ( .A1(\mem[20][26] ), .A2(n3304), .ZN(n689) );
  NAND2_X2 U1269 ( .A1(\mem[20][25] ), .A2(n3304), .ZN(n690) );
  NAND2_X2 U1271 ( .A1(\mem[20][24] ), .A2(n3304), .ZN(n691) );
  NAND2_X2 U1273 ( .A1(\mem[20][23] ), .A2(n3304), .ZN(n692) );
  NAND2_X2 U1275 ( .A1(\mem[20][22] ), .A2(n3304), .ZN(n693) );
  NAND2_X2 U1277 ( .A1(\mem[20][21] ), .A2(n3304), .ZN(n694) );
  NAND2_X2 U1279 ( .A1(\mem[20][20] ), .A2(n3304), .ZN(n695) );
  NAND2_X2 U1281 ( .A1(\mem[20][1] ), .A2(n3304), .ZN(n696) );
  NAND2_X2 U1283 ( .A1(\mem[20][19] ), .A2(n3304), .ZN(n697) );
  NAND2_X2 U1285 ( .A1(\mem[20][18] ), .A2(n3304), .ZN(n698) );
  NAND2_X2 U1287 ( .A1(\mem[20][17] ), .A2(n3304), .ZN(n699) );
  NAND2_X2 U1289 ( .A1(\mem[20][16] ), .A2(n3304), .ZN(n700) );
  NAND2_X2 U1291 ( .A1(\mem[20][15] ), .A2(n3304), .ZN(n701) );
  NAND2_X2 U1293 ( .A1(\mem[20][14] ), .A2(n3304), .ZN(n702) );
  NAND2_X2 U1295 ( .A1(\mem[20][13] ), .A2(n3304), .ZN(n703) );
  NAND2_X2 U1297 ( .A1(\mem[20][12] ), .A2(n3303), .ZN(n704) );
  NAND2_X2 U1299 ( .A1(\mem[20][11] ), .A2(n3304), .ZN(n705) );
  NAND2_X2 U1301 ( .A1(\mem[20][10] ), .A2(n3302), .ZN(n706) );
  NAND2_X2 U1303 ( .A1(\mem[20][0] ), .A2(n3304), .ZN(n707) );
  NAND2_X2 U1304 ( .A1(n608), .A2(n101), .ZN(n675) );
  AND2_X2 U1305 ( .A1(n439), .A2(n237), .ZN(n608) );
  NAND2_X2 U1308 ( .A1(\mem[1][9] ), .A2(n3300), .ZN(n710) );
  NAND2_X2 U1310 ( .A1(\mem[1][8] ), .A2(n3298), .ZN(n711) );
  NAND2_X2 U1312 ( .A1(\mem[1][7] ), .A2(n3299), .ZN(n712) );
  NAND2_X2 U1314 ( .A1(\mem[1][6] ), .A2(n3298), .ZN(n713) );
  NAND2_X2 U1316 ( .A1(\mem[1][5] ), .A2(n3299), .ZN(n714) );
  NAND2_X2 U1318 ( .A1(\mem[1][4] ), .A2(n3298), .ZN(n715) );
  NAND2_X2 U1320 ( .A1(\mem[1][3] ), .A2(n3299), .ZN(n716) );
  NAND2_X2 U1322 ( .A1(\mem[1][31] ), .A2(n3300), .ZN(n717) );
  NAND2_X2 U1324 ( .A1(\mem[1][30] ), .A2(n3300), .ZN(n718) );
  NAND2_X2 U1326 ( .A1(\mem[1][2] ), .A2(n3300), .ZN(n719) );
  NAND2_X2 U1328 ( .A1(\mem[1][29] ), .A2(n3300), .ZN(n720) );
  NAND2_X2 U1330 ( .A1(\mem[1][28] ), .A2(n3300), .ZN(n721) );
  NAND2_X2 U1332 ( .A1(\mem[1][27] ), .A2(n3300), .ZN(n722) );
  NAND2_X2 U1334 ( .A1(\mem[1][26] ), .A2(n3300), .ZN(n723) );
  NAND2_X2 U1336 ( .A1(\mem[1][25] ), .A2(n3300), .ZN(n724) );
  NAND2_X2 U1338 ( .A1(\mem[1][24] ), .A2(n3300), .ZN(n725) );
  NAND2_X2 U1340 ( .A1(\mem[1][23] ), .A2(n3300), .ZN(n726) );
  NAND2_X2 U1342 ( .A1(\mem[1][22] ), .A2(n3300), .ZN(n727) );
  NAND2_X2 U1344 ( .A1(\mem[1][21] ), .A2(n3300), .ZN(n728) );
  NAND2_X2 U1346 ( .A1(\mem[1][20] ), .A2(n3300), .ZN(n729) );
  NAND2_X2 U1348 ( .A1(\mem[1][1] ), .A2(n3300), .ZN(n730) );
  NAND2_X2 U1350 ( .A1(\mem[1][19] ), .A2(n3300), .ZN(n731) );
  NAND2_X2 U1352 ( .A1(\mem[1][18] ), .A2(n3300), .ZN(n732) );
  NAND2_X2 U1354 ( .A1(\mem[1][17] ), .A2(n3300), .ZN(n733) );
  NAND2_X2 U1356 ( .A1(\mem[1][16] ), .A2(n3300), .ZN(n734) );
  NAND2_X2 U1358 ( .A1(\mem[1][15] ), .A2(n3300), .ZN(n735) );
  NAND2_X2 U1360 ( .A1(\mem[1][14] ), .A2(n3300), .ZN(n736) );
  NAND2_X2 U1362 ( .A1(\mem[1][13] ), .A2(n3300), .ZN(n737) );
  NAND2_X2 U1364 ( .A1(\mem[1][12] ), .A2(n3299), .ZN(n738) );
  NAND2_X2 U1366 ( .A1(\mem[1][11] ), .A2(n3300), .ZN(n739) );
  NAND2_X2 U1368 ( .A1(\mem[1][10] ), .A2(n3298), .ZN(n740) );
  NAND2_X2 U1370 ( .A1(\mem[1][0] ), .A2(n3300), .ZN(n741) );
  NAND2_X2 U1371 ( .A1(n272), .A2(n66), .ZN(n709) );
  NAND2_X2 U1373 ( .A1(\mem[19][9] ), .A2(n3296), .ZN(n743) );
  NAND2_X2 U1375 ( .A1(\mem[19][8] ), .A2(n3295), .ZN(n744) );
  NAND2_X2 U1377 ( .A1(\mem[19][7] ), .A2(n3296), .ZN(n745) );
  NAND2_X2 U1379 ( .A1(\mem[19][6] ), .A2(n3295), .ZN(n746) );
  NAND2_X2 U1381 ( .A1(\mem[19][5] ), .A2(n3296), .ZN(n747) );
  NAND2_X2 U1383 ( .A1(\mem[19][4] ), .A2(n3295), .ZN(n748) );
  NAND2_X2 U1385 ( .A1(\mem[19][3] ), .A2(n3296), .ZN(n749) );
  NAND2_X2 U1387 ( .A1(\mem[19][31] ), .A2(n3297), .ZN(n750) );
  NAND2_X2 U1389 ( .A1(\mem[19][30] ), .A2(n3297), .ZN(n751) );
  NAND2_X2 U1391 ( .A1(\mem[19][2] ), .A2(n3297), .ZN(n752) );
  NAND2_X2 U1393 ( .A1(\mem[19][29] ), .A2(n3297), .ZN(n753) );
  NAND2_X2 U1395 ( .A1(\mem[19][28] ), .A2(n3297), .ZN(n754) );
  NAND2_X2 U1397 ( .A1(\mem[19][27] ), .A2(n3297), .ZN(n755) );
  NAND2_X2 U1399 ( .A1(\mem[19][26] ), .A2(n3297), .ZN(n756) );
  NAND2_X2 U1401 ( .A1(\mem[19][25] ), .A2(n3297), .ZN(n757) );
  NAND2_X2 U1403 ( .A1(\mem[19][24] ), .A2(n3297), .ZN(n758) );
  NAND2_X2 U1405 ( .A1(\mem[19][23] ), .A2(n3297), .ZN(n759) );
  NAND2_X2 U1407 ( .A1(\mem[19][22] ), .A2(n3297), .ZN(n760) );
  NAND2_X2 U1409 ( .A1(\mem[19][21] ), .A2(n3297), .ZN(n761) );
  NAND2_X2 U1411 ( .A1(\mem[19][20] ), .A2(n3297), .ZN(n762) );
  NAND2_X2 U1413 ( .A1(\mem[19][1] ), .A2(n3297), .ZN(n763) );
  NAND2_X2 U1415 ( .A1(\mem[19][19] ), .A2(n3297), .ZN(n764) );
  NAND2_X2 U1417 ( .A1(\mem[19][18] ), .A2(n3297), .ZN(n765) );
  NAND2_X2 U1419 ( .A1(\mem[19][17] ), .A2(n3297), .ZN(n766) );
  NAND2_X2 U1421 ( .A1(\mem[19][16] ), .A2(n3297), .ZN(n767) );
  NAND2_X2 U1423 ( .A1(\mem[19][15] ), .A2(n3297), .ZN(n768) );
  NAND2_X2 U1425 ( .A1(\mem[19][14] ), .A2(n3297), .ZN(n769) );
  NAND2_X2 U1427 ( .A1(\mem[19][13] ), .A2(n3297), .ZN(n770) );
  NAND2_X2 U1429 ( .A1(\mem[19][12] ), .A2(n3297), .ZN(n771) );
  NAND2_X2 U1431 ( .A1(\mem[19][11] ), .A2(n3297), .ZN(n772) );
  NAND2_X2 U1433 ( .A1(\mem[19][10] ), .A2(n3297), .ZN(n773) );
  NAND2_X2 U1435 ( .A1(\mem[19][0] ), .A2(n3297), .ZN(n774) );
  NAND2_X2 U1436 ( .A1(n775), .A2(n135), .ZN(n742) );
  NAND2_X2 U1438 ( .A1(\mem[18][9] ), .A2(n3292), .ZN(n777) );
  NAND2_X2 U1440 ( .A1(\mem[18][8] ), .A2(n3291), .ZN(n778) );
  NAND2_X2 U1442 ( .A1(\mem[18][7] ), .A2(n3292), .ZN(n779) );
  NAND2_X2 U1444 ( .A1(\mem[18][6] ), .A2(n3291), .ZN(n780) );
  NAND2_X2 U1446 ( .A1(\mem[18][5] ), .A2(n3292), .ZN(n781) );
  NAND2_X2 U1448 ( .A1(\mem[18][4] ), .A2(n3291), .ZN(n782) );
  NAND2_X2 U1450 ( .A1(\mem[18][3] ), .A2(n3292), .ZN(n783) );
  NAND2_X2 U1452 ( .A1(\mem[18][31] ), .A2(n3293), .ZN(n784) );
  NAND2_X2 U1454 ( .A1(\mem[18][30] ), .A2(n3293), .ZN(n785) );
  NAND2_X2 U1456 ( .A1(\mem[18][2] ), .A2(n3293), .ZN(n786) );
  NAND2_X2 U1458 ( .A1(\mem[18][29] ), .A2(n3293), .ZN(n787) );
  NAND2_X2 U1460 ( .A1(\mem[18][28] ), .A2(n3293), .ZN(n788) );
  NAND2_X2 U1462 ( .A1(\mem[18][27] ), .A2(n3293), .ZN(n789) );
  NAND2_X2 U1464 ( .A1(\mem[18][26] ), .A2(n3293), .ZN(n790) );
  NAND2_X2 U1466 ( .A1(\mem[18][25] ), .A2(n3293), .ZN(n791) );
  NAND2_X2 U1468 ( .A1(\mem[18][24] ), .A2(n3293), .ZN(n792) );
  NAND2_X2 U1470 ( .A1(\mem[18][23] ), .A2(n3293), .ZN(n793) );
  NAND2_X2 U1472 ( .A1(\mem[18][22] ), .A2(n3293), .ZN(n794) );
  NAND2_X2 U1474 ( .A1(\mem[18][21] ), .A2(n3293), .ZN(n795) );
  NAND2_X2 U1476 ( .A1(\mem[18][20] ), .A2(n3293), .ZN(n796) );
  NAND2_X2 U1478 ( .A1(\mem[18][1] ), .A2(n3293), .ZN(n797) );
  NAND2_X2 U1480 ( .A1(\mem[18][19] ), .A2(n3293), .ZN(n798) );
  NAND2_X2 U1482 ( .A1(\mem[18][18] ), .A2(n3293), .ZN(n799) );
  NAND2_X2 U1484 ( .A1(\mem[18][17] ), .A2(n3293), .ZN(n800) );
  NAND2_X2 U1486 ( .A1(\mem[18][16] ), .A2(n3293), .ZN(n801) );
  NAND2_X2 U1488 ( .A1(\mem[18][15] ), .A2(n3293), .ZN(n802) );
  NAND2_X2 U1490 ( .A1(\mem[18][14] ), .A2(n3293), .ZN(n803) );
  NAND2_X2 U1492 ( .A1(\mem[18][13] ), .A2(n3293), .ZN(n804) );
  NAND2_X2 U1494 ( .A1(\mem[18][12] ), .A2(n3293), .ZN(n805) );
  NAND2_X2 U1496 ( .A1(\mem[18][11] ), .A2(n3293), .ZN(n806) );
  NAND2_X2 U1498 ( .A1(\mem[18][10] ), .A2(n3293), .ZN(n807) );
  NAND2_X2 U1500 ( .A1(\mem[18][0] ), .A2(n3293), .ZN(n808) );
  NAND2_X2 U1501 ( .A1(n775), .A2(n170), .ZN(n776) );
  NAND2_X2 U1503 ( .A1(\mem[17][9] ), .A2(n3288), .ZN(n810) );
  NAND2_X2 U1505 ( .A1(\mem[17][8] ), .A2(n3286), .ZN(n811) );
  NAND2_X2 U1507 ( .A1(\mem[17][7] ), .A2(n3287), .ZN(n812) );
  NAND2_X2 U1509 ( .A1(\mem[17][6] ), .A2(n3286), .ZN(n813) );
  NAND2_X2 U1511 ( .A1(\mem[17][5] ), .A2(n3287), .ZN(n814) );
  NAND2_X2 U1513 ( .A1(\mem[17][4] ), .A2(n3286), .ZN(n815) );
  NAND2_X2 U1515 ( .A1(\mem[17][3] ), .A2(n3287), .ZN(n816) );
  NAND2_X2 U1517 ( .A1(\mem[17][31] ), .A2(n3288), .ZN(n817) );
  NAND2_X2 U1519 ( .A1(\mem[17][30] ), .A2(n3288), .ZN(n818) );
  NAND2_X2 U1521 ( .A1(\mem[17][2] ), .A2(n3288), .ZN(n819) );
  NAND2_X2 U1523 ( .A1(\mem[17][29] ), .A2(n3288), .ZN(n820) );
  NAND2_X2 U1525 ( .A1(\mem[17][28] ), .A2(n3288), .ZN(n821) );
  NAND2_X2 U1527 ( .A1(\mem[17][27] ), .A2(n3288), .ZN(n822) );
  NAND2_X2 U1529 ( .A1(\mem[17][26] ), .A2(n3288), .ZN(n823) );
  NAND2_X2 U1531 ( .A1(\mem[17][25] ), .A2(n3288), .ZN(n824) );
  NAND2_X2 U1533 ( .A1(\mem[17][24] ), .A2(n3288), .ZN(n825) );
  NAND2_X2 U1535 ( .A1(\mem[17][23] ), .A2(n3288), .ZN(n826) );
  NAND2_X2 U1537 ( .A1(\mem[17][22] ), .A2(n3288), .ZN(n827) );
  NAND2_X2 U1539 ( .A1(\mem[17][21] ), .A2(n3288), .ZN(n828) );
  NAND2_X2 U1541 ( .A1(\mem[17][20] ), .A2(n3288), .ZN(n829) );
  NAND2_X2 U1543 ( .A1(\mem[17][1] ), .A2(n3288), .ZN(n830) );
  NAND2_X2 U1545 ( .A1(\mem[17][19] ), .A2(n3288), .ZN(n831) );
  NAND2_X2 U1547 ( .A1(\mem[17][18] ), .A2(n3288), .ZN(n832) );
  NAND2_X2 U1549 ( .A1(\mem[17][17] ), .A2(n3288), .ZN(n833) );
  NAND2_X2 U1551 ( .A1(\mem[17][16] ), .A2(n3288), .ZN(n834) );
  NAND2_X2 U1553 ( .A1(\mem[17][15] ), .A2(n3288), .ZN(n835) );
  NAND2_X2 U1555 ( .A1(\mem[17][14] ), .A2(n3288), .ZN(n836) );
  NAND2_X2 U1557 ( .A1(\mem[17][13] ), .A2(n3288), .ZN(n837) );
  NAND2_X2 U1559 ( .A1(\mem[17][12] ), .A2(n3287), .ZN(n838) );
  NAND2_X2 U1561 ( .A1(\mem[17][11] ), .A2(n3288), .ZN(n839) );
  NAND2_X2 U1563 ( .A1(\mem[17][10] ), .A2(n3286), .ZN(n840) );
  NAND2_X2 U1565 ( .A1(\mem[17][0] ), .A2(n3288), .ZN(n841) );
  NAND2_X2 U1566 ( .A1(n775), .A2(n66), .ZN(n809) );
  NAND2_X2 U1568 ( .A1(\mem[16][9] ), .A2(n3284), .ZN(n843) );
  NAND2_X2 U1570 ( .A1(\mem[16][8] ), .A2(n3282), .ZN(n844) );
  NAND2_X2 U1572 ( .A1(\mem[16][7] ), .A2(n3283), .ZN(n845) );
  NAND2_X2 U1574 ( .A1(\mem[16][6] ), .A2(n3282), .ZN(n846) );
  NAND2_X2 U1576 ( .A1(\mem[16][5] ), .A2(n3283), .ZN(n847) );
  NAND2_X2 U1578 ( .A1(\mem[16][4] ), .A2(n3282), .ZN(n848) );
  NAND2_X2 U1580 ( .A1(\mem[16][3] ), .A2(n3283), .ZN(n849) );
  NAND2_X2 U1582 ( .A1(\mem[16][31] ), .A2(n3284), .ZN(n850) );
  NAND2_X2 U1584 ( .A1(\mem[16][30] ), .A2(n3284), .ZN(n851) );
  NAND2_X2 U1586 ( .A1(\mem[16][2] ), .A2(n3284), .ZN(n852) );
  NAND2_X2 U1588 ( .A1(\mem[16][29] ), .A2(n3284), .ZN(n853) );
  NAND2_X2 U1590 ( .A1(\mem[16][28] ), .A2(n3284), .ZN(n854) );
  NAND2_X2 U1592 ( .A1(\mem[16][27] ), .A2(n3284), .ZN(n855) );
  NAND2_X2 U1594 ( .A1(\mem[16][26] ), .A2(n3284), .ZN(n856) );
  NAND2_X2 U1596 ( .A1(\mem[16][25] ), .A2(n3284), .ZN(n857) );
  NAND2_X2 U1598 ( .A1(\mem[16][24] ), .A2(n3284), .ZN(n858) );
  NAND2_X2 U1600 ( .A1(\mem[16][23] ), .A2(n3284), .ZN(n859) );
  NAND2_X2 U1602 ( .A1(\mem[16][22] ), .A2(n3284), .ZN(n860) );
  NAND2_X2 U1604 ( .A1(\mem[16][21] ), .A2(n3284), .ZN(n861) );
  NAND2_X2 U1606 ( .A1(\mem[16][20] ), .A2(n3284), .ZN(n862) );
  NAND2_X2 U1608 ( .A1(\mem[16][1] ), .A2(n3284), .ZN(n863) );
  NAND2_X2 U1610 ( .A1(\mem[16][19] ), .A2(n3284), .ZN(n864) );
  NAND2_X2 U1612 ( .A1(\mem[16][18] ), .A2(n3284), .ZN(n865) );
  NAND2_X2 U1614 ( .A1(\mem[16][17] ), .A2(n3284), .ZN(n866) );
  NAND2_X2 U1616 ( .A1(\mem[16][16] ), .A2(n3284), .ZN(n867) );
  NAND2_X2 U1618 ( .A1(\mem[16][15] ), .A2(n3284), .ZN(n868) );
  NAND2_X2 U1620 ( .A1(\mem[16][14] ), .A2(n3284), .ZN(n869) );
  NAND2_X2 U1622 ( .A1(\mem[16][13] ), .A2(n3284), .ZN(n870) );
  NAND2_X2 U1624 ( .A1(\mem[16][12] ), .A2(n3283), .ZN(n871) );
  NAND2_X2 U1626 ( .A1(\mem[16][11] ), .A2(n3284), .ZN(n872) );
  NAND2_X2 U1628 ( .A1(\mem[16][10] ), .A2(n3282), .ZN(n873) );
  NAND2_X2 U1630 ( .A1(\mem[16][0] ), .A2(n3284), .ZN(n874) );
  NAND2_X2 U1631 ( .A1(n775), .A2(n101), .ZN(n842) );
  AND2_X2 U1632 ( .A1(n439), .A2(n875), .ZN(n775) );
  NAND2_X2 U1636 ( .A1(\mem[15][9] ), .A2(n3280), .ZN(n879) );
  NAND2_X2 U1638 ( .A1(\mem[15][8] ), .A2(n3279), .ZN(n880) );
  NAND2_X2 U1640 ( .A1(\mem[15][7] ), .A2(n3280), .ZN(n881) );
  NAND2_X2 U1642 ( .A1(\mem[15][6] ), .A2(n3279), .ZN(n882) );
  NAND2_X2 U1644 ( .A1(\mem[15][5] ), .A2(n3280), .ZN(n883) );
  NAND2_X2 U1646 ( .A1(\mem[15][4] ), .A2(n3279), .ZN(n884) );
  NAND2_X2 U1648 ( .A1(\mem[15][3] ), .A2(n3280), .ZN(n885) );
  NAND2_X2 U1650 ( .A1(\mem[15][31] ), .A2(n3281), .ZN(n886) );
  NAND2_X2 U1652 ( .A1(\mem[15][30] ), .A2(n3281), .ZN(n887) );
  NAND2_X2 U1654 ( .A1(\mem[15][2] ), .A2(n3281), .ZN(n888) );
  NAND2_X2 U1656 ( .A1(\mem[15][29] ), .A2(n3281), .ZN(n889) );
  NAND2_X2 U1658 ( .A1(\mem[15][28] ), .A2(n3281), .ZN(n890) );
  NAND2_X2 U1660 ( .A1(\mem[15][27] ), .A2(n3281), .ZN(n891) );
  NAND2_X2 U1662 ( .A1(\mem[15][26] ), .A2(n3281), .ZN(n892) );
  NAND2_X2 U1664 ( .A1(\mem[15][25] ), .A2(n3281), .ZN(n893) );
  NAND2_X2 U1666 ( .A1(\mem[15][24] ), .A2(n3281), .ZN(n894) );
  NAND2_X2 U1668 ( .A1(\mem[15][23] ), .A2(n3281), .ZN(n895) );
  NAND2_X2 U1670 ( .A1(\mem[15][22] ), .A2(n3281), .ZN(n896) );
  NAND2_X2 U1672 ( .A1(\mem[15][21] ), .A2(n3281), .ZN(n897) );
  NAND2_X2 U1674 ( .A1(\mem[15][20] ), .A2(n3281), .ZN(n898) );
  NAND2_X2 U1676 ( .A1(\mem[15][1] ), .A2(n3281), .ZN(n899) );
  NAND2_X2 U1678 ( .A1(\mem[15][19] ), .A2(n3281), .ZN(n900) );
  NAND2_X2 U1680 ( .A1(\mem[15][18] ), .A2(n3281), .ZN(n901) );
  NAND2_X2 U1682 ( .A1(\mem[15][17] ), .A2(n3281), .ZN(n902) );
  NAND2_X2 U1684 ( .A1(\mem[15][16] ), .A2(n3281), .ZN(n903) );
  NAND2_X2 U1686 ( .A1(\mem[15][15] ), .A2(n3281), .ZN(n904) );
  NAND2_X2 U1688 ( .A1(\mem[15][14] ), .A2(n3281), .ZN(n905) );
  NAND2_X2 U1690 ( .A1(\mem[15][13] ), .A2(n3281), .ZN(n906) );
  NAND2_X2 U1692 ( .A1(\mem[15][12] ), .A2(n3281), .ZN(n907) );
  NAND2_X2 U1694 ( .A1(\mem[15][11] ), .A2(n3281), .ZN(n908) );
  NAND2_X2 U1696 ( .A1(\mem[15][10] ), .A2(n3281), .ZN(n909) );
  NAND2_X2 U1698 ( .A1(\mem[15][0] ), .A2(n3281), .ZN(n910) );
  NAND2_X2 U1699 ( .A1(n911), .A2(n135), .ZN(n878) );
  NAND2_X2 U1701 ( .A1(\mem[14][9] ), .A2(n3276), .ZN(n913) );
  NAND2_X2 U1703 ( .A1(\mem[14][8] ), .A2(n3275), .ZN(n914) );
  NAND2_X2 U1705 ( .A1(\mem[14][7] ), .A2(n3276), .ZN(n915) );
  NAND2_X2 U1707 ( .A1(\mem[14][6] ), .A2(n3275), .ZN(n916) );
  NAND2_X2 U1709 ( .A1(\mem[14][5] ), .A2(n3276), .ZN(n917) );
  NAND2_X2 U1711 ( .A1(\mem[14][4] ), .A2(n3275), .ZN(n918) );
  NAND2_X2 U1713 ( .A1(\mem[14][3] ), .A2(n3276), .ZN(n919) );
  NAND2_X2 U1715 ( .A1(\mem[14][31] ), .A2(n3277), .ZN(n920) );
  NAND2_X2 U1717 ( .A1(\mem[14][30] ), .A2(n3277), .ZN(n921) );
  NAND2_X2 U1719 ( .A1(\mem[14][2] ), .A2(n3277), .ZN(n922) );
  NAND2_X2 U1721 ( .A1(\mem[14][29] ), .A2(n3277), .ZN(n923) );
  NAND2_X2 U1723 ( .A1(\mem[14][28] ), .A2(n3277), .ZN(n924) );
  NAND2_X2 U1725 ( .A1(\mem[14][27] ), .A2(n3277), .ZN(n925) );
  NAND2_X2 U1727 ( .A1(\mem[14][26] ), .A2(n3277), .ZN(n926) );
  NAND2_X2 U1729 ( .A1(\mem[14][25] ), .A2(n3277), .ZN(n927) );
  NAND2_X2 U1731 ( .A1(\mem[14][24] ), .A2(n3277), .ZN(n928) );
  NAND2_X2 U1733 ( .A1(\mem[14][23] ), .A2(n3277), .ZN(n929) );
  NAND2_X2 U1735 ( .A1(\mem[14][22] ), .A2(n3277), .ZN(n930) );
  NAND2_X2 U1737 ( .A1(\mem[14][21] ), .A2(n3277), .ZN(n931) );
  NAND2_X2 U1739 ( .A1(\mem[14][20] ), .A2(n3277), .ZN(n932) );
  NAND2_X2 U1741 ( .A1(\mem[14][1] ), .A2(n3277), .ZN(n933) );
  NAND2_X2 U1743 ( .A1(\mem[14][19] ), .A2(n3277), .ZN(n934) );
  NAND2_X2 U1745 ( .A1(\mem[14][18] ), .A2(n3277), .ZN(n935) );
  NAND2_X2 U1747 ( .A1(\mem[14][17] ), .A2(n3277), .ZN(n936) );
  NAND2_X2 U1749 ( .A1(\mem[14][16] ), .A2(n3277), .ZN(n937) );
  NAND2_X2 U1751 ( .A1(\mem[14][15] ), .A2(n3277), .ZN(n938) );
  NAND2_X2 U1753 ( .A1(\mem[14][14] ), .A2(n3277), .ZN(n939) );
  NAND2_X2 U1755 ( .A1(\mem[14][13] ), .A2(n3277), .ZN(n940) );
  NAND2_X2 U1757 ( .A1(\mem[14][12] ), .A2(n3277), .ZN(n941) );
  NAND2_X2 U1759 ( .A1(\mem[14][11] ), .A2(n3277), .ZN(n942) );
  NAND2_X2 U1761 ( .A1(\mem[14][10] ), .A2(n3277), .ZN(n943) );
  NAND2_X2 U1763 ( .A1(\mem[14][0] ), .A2(n3277), .ZN(n944) );
  NAND2_X2 U1764 ( .A1(n911), .A2(n170), .ZN(n912) );
  NAND2_X2 U1766 ( .A1(\mem[13][9] ), .A2(n3272), .ZN(n946) );
  NAND2_X2 U1768 ( .A1(\mem[13][8] ), .A2(n3270), .ZN(n947) );
  NAND2_X2 U1770 ( .A1(\mem[13][7] ), .A2(n3271), .ZN(n948) );
  NAND2_X2 U1772 ( .A1(\mem[13][6] ), .A2(n3270), .ZN(n949) );
  NAND2_X2 U1774 ( .A1(\mem[13][5] ), .A2(n3271), .ZN(n950) );
  NAND2_X2 U1776 ( .A1(\mem[13][4] ), .A2(n3270), .ZN(n951) );
  NAND2_X2 U1778 ( .A1(\mem[13][3] ), .A2(n3271), .ZN(n952) );
  NAND2_X2 U1780 ( .A1(\mem[13][31] ), .A2(n3272), .ZN(n953) );
  NAND2_X2 U1782 ( .A1(\mem[13][30] ), .A2(n3272), .ZN(n954) );
  NAND2_X2 U1784 ( .A1(\mem[13][2] ), .A2(n3272), .ZN(n955) );
  NAND2_X2 U1786 ( .A1(\mem[13][29] ), .A2(n3272), .ZN(n956) );
  NAND2_X2 U1788 ( .A1(\mem[13][28] ), .A2(n3272), .ZN(n957) );
  NAND2_X2 U1790 ( .A1(\mem[13][27] ), .A2(n3272), .ZN(n958) );
  NAND2_X2 U1792 ( .A1(\mem[13][26] ), .A2(n3272), .ZN(n959) );
  NAND2_X2 U1794 ( .A1(\mem[13][25] ), .A2(n3272), .ZN(n960) );
  NAND2_X2 U1796 ( .A1(\mem[13][24] ), .A2(n3272), .ZN(n961) );
  NAND2_X2 U1798 ( .A1(\mem[13][23] ), .A2(n3272), .ZN(n962) );
  NAND2_X2 U1800 ( .A1(\mem[13][22] ), .A2(n3272), .ZN(n963) );
  NAND2_X2 U1802 ( .A1(\mem[13][21] ), .A2(n3272), .ZN(n964) );
  NAND2_X2 U1804 ( .A1(\mem[13][20] ), .A2(n3272), .ZN(n965) );
  NAND2_X2 U1806 ( .A1(\mem[13][1] ), .A2(n3272), .ZN(n966) );
  NAND2_X2 U1808 ( .A1(\mem[13][19] ), .A2(n3272), .ZN(n967) );
  NAND2_X2 U1810 ( .A1(\mem[13][18] ), .A2(n3272), .ZN(n968) );
  NAND2_X2 U1812 ( .A1(\mem[13][17] ), .A2(n3272), .ZN(n969) );
  NAND2_X2 U1814 ( .A1(\mem[13][16] ), .A2(n3272), .ZN(n970) );
  NAND2_X2 U1816 ( .A1(\mem[13][15] ), .A2(n3272), .ZN(n971) );
  NAND2_X2 U1818 ( .A1(\mem[13][14] ), .A2(n3272), .ZN(n972) );
  NAND2_X2 U1820 ( .A1(\mem[13][13] ), .A2(n3272), .ZN(n973) );
  NAND2_X2 U1822 ( .A1(\mem[13][12] ), .A2(n3271), .ZN(n974) );
  NAND2_X2 U1824 ( .A1(\mem[13][11] ), .A2(n3272), .ZN(n975) );
  NAND2_X2 U1826 ( .A1(\mem[13][10] ), .A2(n3270), .ZN(n976) );
  NAND2_X2 U1828 ( .A1(\mem[13][0] ), .A2(n3272), .ZN(n977) );
  NAND2_X2 U1829 ( .A1(n911), .A2(n66), .ZN(n945) );
  NAND2_X2 U1832 ( .A1(\mem[12][9] ), .A2(n3268), .ZN(n980) );
  NAND2_X2 U1834 ( .A1(\mem[12][8] ), .A2(n3266), .ZN(n981) );
  NAND2_X2 U1836 ( .A1(\mem[12][7] ), .A2(n3267), .ZN(n982) );
  NAND2_X2 U1838 ( .A1(\mem[12][6] ), .A2(n3266), .ZN(n983) );
  NAND2_X2 U1840 ( .A1(\mem[12][5] ), .A2(n3267), .ZN(n984) );
  NAND2_X2 U1842 ( .A1(\mem[12][4] ), .A2(n3266), .ZN(n985) );
  NAND2_X2 U1844 ( .A1(\mem[12][3] ), .A2(n3267), .ZN(n986) );
  NAND2_X2 U1846 ( .A1(\mem[12][31] ), .A2(n3268), .ZN(n987) );
  NAND2_X2 U1848 ( .A1(\mem[12][30] ), .A2(n3268), .ZN(n988) );
  NAND2_X2 U1850 ( .A1(\mem[12][2] ), .A2(n3268), .ZN(n989) );
  NAND2_X2 U1852 ( .A1(\mem[12][29] ), .A2(n3268), .ZN(n990) );
  NAND2_X2 U1854 ( .A1(\mem[12][28] ), .A2(n3268), .ZN(n991) );
  NAND2_X2 U1856 ( .A1(\mem[12][27] ), .A2(n3268), .ZN(n992) );
  NAND2_X2 U1858 ( .A1(\mem[12][26] ), .A2(n3268), .ZN(n993) );
  NAND2_X2 U1860 ( .A1(\mem[12][25] ), .A2(n3268), .ZN(n994) );
  NAND2_X2 U1862 ( .A1(\mem[12][24] ), .A2(n3268), .ZN(n995) );
  NAND2_X2 U1864 ( .A1(\mem[12][23] ), .A2(n3268), .ZN(n996) );
  NAND2_X2 U1866 ( .A1(\mem[12][22] ), .A2(n3268), .ZN(n997) );
  NAND2_X2 U1868 ( .A1(\mem[12][21] ), .A2(n3268), .ZN(n998) );
  NAND2_X2 U1870 ( .A1(\mem[12][20] ), .A2(n3268), .ZN(n999) );
  NAND2_X2 U1872 ( .A1(\mem[12][1] ), .A2(n3268), .ZN(n1000) );
  NAND2_X2 U1874 ( .A1(\mem[12][19] ), .A2(n3268), .ZN(n1001) );
  NAND2_X2 U1876 ( .A1(\mem[12][18] ), .A2(n3268), .ZN(n1002) );
  NAND2_X2 U1878 ( .A1(\mem[12][17] ), .A2(n3268), .ZN(n1003) );
  NAND2_X2 U1880 ( .A1(\mem[12][16] ), .A2(n3268), .ZN(n1004) );
  NAND2_X2 U1882 ( .A1(\mem[12][15] ), .A2(n3268), .ZN(n1005) );
  NAND2_X2 U1884 ( .A1(\mem[12][14] ), .A2(n3268), .ZN(n1006) );
  NAND2_X2 U1886 ( .A1(\mem[12][13] ), .A2(n3268), .ZN(n1007) );
  NAND2_X2 U1888 ( .A1(\mem[12][12] ), .A2(n3267), .ZN(n1008) );
  NAND2_X2 U1890 ( .A1(\mem[12][11] ), .A2(n3268), .ZN(n1009) );
  NAND2_X2 U1892 ( .A1(\mem[12][10] ), .A2(n3266), .ZN(n1010) );
  NAND2_X2 U1894 ( .A1(\mem[12][0] ), .A2(n3268), .ZN(n1011) );
  NAND2_X2 U1895 ( .A1(n911), .A2(n101), .ZN(n979) );
  AND2_X2 U1896 ( .A1(n440), .A2(n238), .ZN(n911) );
  NAND2_X2 U1900 ( .A1(\mem[11][9] ), .A2(n3264), .ZN(n1014) );
  NAND2_X2 U1902 ( .A1(\mem[11][8] ), .A2(n3263), .ZN(n1015) );
  NAND2_X2 U1904 ( .A1(\mem[11][7] ), .A2(n3264), .ZN(n1016) );
  NAND2_X2 U1906 ( .A1(\mem[11][6] ), .A2(n3263), .ZN(n1017) );
  NAND2_X2 U1908 ( .A1(\mem[11][5] ), .A2(n3264), .ZN(n1018) );
  NAND2_X2 U1910 ( .A1(\mem[11][4] ), .A2(n3263), .ZN(n1019) );
  NAND2_X2 U1912 ( .A1(\mem[11][3] ), .A2(n3264), .ZN(n1020) );
  NAND2_X2 U1914 ( .A1(\mem[11][31] ), .A2(n3265), .ZN(n1021) );
  NAND2_X2 U1916 ( .A1(\mem[11][30] ), .A2(n3265), .ZN(n1022) );
  NAND2_X2 U1918 ( .A1(\mem[11][2] ), .A2(n3265), .ZN(n1023) );
  NAND2_X2 U1920 ( .A1(\mem[11][29] ), .A2(n3265), .ZN(n1024) );
  NAND2_X2 U1922 ( .A1(\mem[11][28] ), .A2(n3265), .ZN(n1025) );
  NAND2_X2 U1924 ( .A1(\mem[11][27] ), .A2(n3265), .ZN(n1026) );
  NAND2_X2 U1926 ( .A1(\mem[11][26] ), .A2(n3265), .ZN(n1027) );
  NAND2_X2 U1928 ( .A1(\mem[11][25] ), .A2(n3265), .ZN(n1028) );
  NAND2_X2 U1930 ( .A1(\mem[11][24] ), .A2(n3265), .ZN(n1029) );
  NAND2_X2 U1932 ( .A1(\mem[11][23] ), .A2(n3265), .ZN(n1030) );
  NAND2_X2 U1934 ( .A1(\mem[11][22] ), .A2(n3265), .ZN(n1031) );
  NAND2_X2 U1936 ( .A1(\mem[11][21] ), .A2(n3265), .ZN(n1032) );
  NAND2_X2 U1938 ( .A1(\mem[11][20] ), .A2(n3265), .ZN(n1033) );
  NAND2_X2 U1940 ( .A1(\mem[11][1] ), .A2(n3265), .ZN(n1034) );
  NAND2_X2 U1942 ( .A1(\mem[11][19] ), .A2(n3265), .ZN(n1035) );
  NAND2_X2 U1944 ( .A1(\mem[11][18] ), .A2(n3265), .ZN(n1036) );
  NAND2_X2 U1946 ( .A1(\mem[11][17] ), .A2(n3265), .ZN(n1037) );
  NAND2_X2 U1948 ( .A1(\mem[11][16] ), .A2(n3265), .ZN(n1038) );
  NAND2_X2 U1950 ( .A1(\mem[11][15] ), .A2(n3265), .ZN(n1039) );
  NAND2_X2 U1952 ( .A1(\mem[11][14] ), .A2(n3265), .ZN(n1040) );
  NAND2_X2 U1954 ( .A1(\mem[11][13] ), .A2(n3265), .ZN(n1041) );
  NAND2_X2 U1956 ( .A1(\mem[11][12] ), .A2(n3265), .ZN(n1042) );
  NAND2_X2 U1958 ( .A1(\mem[11][11] ), .A2(n3265), .ZN(n1043) );
  NAND2_X2 U1960 ( .A1(\mem[11][10] ), .A2(n3265), .ZN(n1044) );
  NAND2_X2 U1962 ( .A1(\mem[11][0] ), .A2(n3265), .ZN(n1045) );
  NAND2_X2 U1963 ( .A1(n135), .A2(n67), .ZN(n1013) );
  AND2_X2 U1964 ( .A1(rd[1]), .A2(rd[0]), .ZN(n135) );
  NAND2_X2 U1966 ( .A1(\mem[10][9] ), .A2(n3260), .ZN(n1047) );
  NAND2_X2 U1968 ( .A1(\mem[10][8] ), .A2(n3259), .ZN(n1048) );
  NAND2_X2 U1970 ( .A1(\mem[10][7] ), .A2(n3260), .ZN(n1049) );
  NAND2_X2 U1972 ( .A1(\mem[10][6] ), .A2(n3259), .ZN(n1050) );
  NAND2_X2 U1974 ( .A1(\mem[10][5] ), .A2(n3260), .ZN(n1051) );
  NAND2_X2 U1976 ( .A1(\mem[10][4] ), .A2(n3259), .ZN(n1052) );
  NAND2_X2 U1978 ( .A1(\mem[10][3] ), .A2(n3260), .ZN(n1053) );
  NAND2_X2 U1980 ( .A1(\mem[10][31] ), .A2(n3261), .ZN(n1054) );
  NAND2_X2 U1982 ( .A1(\mem[10][30] ), .A2(n3261), .ZN(n1055) );
  NAND2_X2 U1984 ( .A1(\mem[10][2] ), .A2(n3261), .ZN(n1056) );
  NAND2_X2 U1986 ( .A1(\mem[10][29] ), .A2(n3261), .ZN(n1057) );
  NAND2_X2 U1988 ( .A1(\mem[10][28] ), .A2(n3261), .ZN(n1058) );
  NAND2_X2 U1990 ( .A1(\mem[10][27] ), .A2(n3261), .ZN(n1059) );
  NAND2_X2 U1992 ( .A1(\mem[10][26] ), .A2(n3261), .ZN(n1060) );
  NAND2_X2 U1994 ( .A1(\mem[10][25] ), .A2(n3261), .ZN(n1061) );
  NAND2_X2 U1996 ( .A1(\mem[10][24] ), .A2(n3261), .ZN(n1062) );
  NAND2_X2 U1998 ( .A1(\mem[10][23] ), .A2(n3261), .ZN(n1063) );
  NAND2_X2 U2000 ( .A1(\mem[10][22] ), .A2(n3261), .ZN(n1064) );
  NAND2_X2 U2002 ( .A1(\mem[10][21] ), .A2(n3261), .ZN(n1065) );
  NAND2_X2 U2004 ( .A1(\mem[10][20] ), .A2(n3261), .ZN(n1066) );
  NAND2_X2 U2006 ( .A1(\mem[10][1] ), .A2(n3261), .ZN(n1067) );
  NAND2_X2 U2008 ( .A1(\mem[10][19] ), .A2(n3261), .ZN(n1068) );
  NAND2_X2 U2010 ( .A1(\mem[10][18] ), .A2(n3261), .ZN(n1069) );
  NAND2_X2 U2012 ( .A1(\mem[10][17] ), .A2(n3261), .ZN(n1070) );
  NAND2_X2 U2014 ( .A1(\mem[10][16] ), .A2(n3261), .ZN(n1071) );
  NAND2_X2 U2016 ( .A1(\mem[10][15] ), .A2(n3261), .ZN(n1072) );
  NAND2_X2 U2018 ( .A1(\mem[10][14] ), .A2(n3261), .ZN(n1073) );
  NAND2_X2 U2020 ( .A1(\mem[10][13] ), .A2(n3261), .ZN(n1074) );
  NAND2_X2 U2022 ( .A1(\mem[10][12] ), .A2(n3261), .ZN(n1075) );
  NAND2_X2 U2024 ( .A1(\mem[10][11] ), .A2(n3261), .ZN(n1076) );
  NAND2_X2 U2026 ( .A1(\mem[10][10] ), .A2(n3261), .ZN(n1077) );
  NAND2_X2 U2028 ( .A1(\mem[10][0] ), .A2(n3261), .ZN(n1078) );
  NAND2_X2 U2029 ( .A1(n170), .A2(n67), .ZN(n1046) );
  AND2_X2 U2030 ( .A1(n238), .A2(n574), .ZN(n67) );
  AND2_X2 U2033 ( .A1(rd[1]), .A2(n4409), .ZN(n170) );
  NAND2_X2 U2036 ( .A1(\mem[0][9] ), .A2(n3256), .ZN(n1080) );
  NAND2_X2 U2039 ( .A1(\mem[0][8] ), .A2(n3254), .ZN(n1081) );
  NAND2_X2 U2042 ( .A1(\mem[0][7] ), .A2(n3255), .ZN(n1082) );
  NAND2_X2 U2045 ( .A1(\mem[0][6] ), .A2(n3254), .ZN(n1083) );
  NAND2_X2 U2048 ( .A1(\mem[0][5] ), .A2(n3255), .ZN(n1084) );
  NAND2_X2 U2051 ( .A1(\mem[0][4] ), .A2(n3254), .ZN(n1085) );
  NAND2_X2 U2054 ( .A1(\mem[0][3] ), .A2(n3255), .ZN(n1086) );
  NAND2_X2 U2057 ( .A1(\mem[0][31] ), .A2(n3256), .ZN(n1087) );
  NAND2_X2 U2060 ( .A1(\mem[0][30] ), .A2(n3256), .ZN(n1088) );
  NAND2_X2 U2063 ( .A1(\mem[0][2] ), .A2(n3256), .ZN(n1089) );
  NAND2_X2 U2066 ( .A1(\mem[0][29] ), .A2(n3256), .ZN(n1090) );
  NAND2_X2 U2069 ( .A1(\mem[0][28] ), .A2(n3256), .ZN(n1091) );
  NAND2_X2 U2072 ( .A1(\mem[0][27] ), .A2(n3256), .ZN(n1092) );
  NAND2_X2 U2075 ( .A1(\mem[0][26] ), .A2(n3256), .ZN(n1093) );
  NAND2_X2 U2078 ( .A1(\mem[0][25] ), .A2(n3256), .ZN(n1094) );
  NAND2_X2 U2081 ( .A1(\mem[0][24] ), .A2(n3256), .ZN(n1095) );
  NAND2_X2 U2084 ( .A1(\mem[0][23] ), .A2(n3256), .ZN(n1096) );
  NAND2_X2 U2087 ( .A1(\mem[0][22] ), .A2(n3256), .ZN(n1097) );
  NAND2_X2 U2090 ( .A1(\mem[0][21] ), .A2(n3256), .ZN(n1098) );
  NAND2_X2 U2093 ( .A1(\mem[0][20] ), .A2(n3256), .ZN(n1099) );
  NAND2_X2 U2096 ( .A1(\mem[0][1] ), .A2(n3256), .ZN(n1100) );
  NAND2_X2 U2099 ( .A1(\mem[0][19] ), .A2(n3256), .ZN(n1101) );
  NAND2_X2 U2102 ( .A1(\mem[0][18] ), .A2(n3256), .ZN(n1102) );
  NAND2_X2 U2105 ( .A1(\mem[0][17] ), .A2(n3256), .ZN(n1103) );
  NAND2_X2 U2108 ( .A1(\mem[0][16] ), .A2(n3256), .ZN(n1104) );
  NAND2_X2 U2111 ( .A1(\mem[0][15] ), .A2(n3256), .ZN(n1105) );
  NAND2_X2 U2114 ( .A1(\mem[0][14] ), .A2(n3256), .ZN(n1106) );
  NAND2_X2 U2117 ( .A1(\mem[0][13] ), .A2(n3256), .ZN(n1107) );
  NAND2_X2 U2120 ( .A1(\mem[0][12] ), .A2(n3255), .ZN(n1108) );
  NAND2_X2 U2123 ( .A1(\mem[0][11] ), .A2(n3256), .ZN(n1109) );
  NAND2_X2 U2126 ( .A1(\mem[0][10] ), .A2(n3254), .ZN(n1110) );
  NAND2_X2 U2129 ( .A1(\mem[0][0] ), .A2(n3256), .ZN(n1111) );
  NAND2_X2 U2130 ( .A1(n272), .A2(n101), .ZN(n1079) );
  AND2_X2 U2132 ( .A1(n875), .A2(n238), .ZN(n272) );
  NAND2_X2 U2134 ( .A1(fp), .A2(n4410), .ZN(n877) );
  NOR2_X2 U2138 ( .A1(rd[0]), .A2(rd[1]), .ZN(n101) );
  NOR2_X2 U2139 ( .A1(n4409), .A2(rd[1]), .ZN(n66) );
  BUF_X4 U2140 ( .A(N9), .Z(n3106) );
  BUF_X4 U2141 ( .A(N9), .Z(n3105) );
  BUF_X4 U2142 ( .A(N9), .Z(n3104) );
  BUF_X4 U2143 ( .A(N9), .Z(n3103) );
  BUF_X4 U2144 ( .A(N9), .Z(n3102) );
  BUF_X4 U2145 ( .A(N9), .Z(n3101) );
  BUF_X4 U2146 ( .A(N9), .Z(n3100) );
  BUF_X4 U2147 ( .A(N9), .Z(n3099) );
  BUF_X4 U2148 ( .A(N9), .Z(n3098) );
  BUF_X4 U2149 ( .A(N9), .Z(n3097) );
  NOR2_X2 U2150 ( .A1(n877), .A2(rd[4]), .ZN(n238) );
  NOR2_X2 U2151 ( .A1(rd[2]), .A2(rd[3]), .ZN(n875) );
  NOR2_X2 U2152 ( .A1(n4408), .A2(rd[3]), .ZN(n237) );
  NOR2_X2 U2153 ( .A1(n4407), .A2(rd[2]), .ZN(n574) );
  NOR2_X2 U2154 ( .A1(n4406), .A2(n877), .ZN(n439) );
  NOR2_X2 U2155 ( .A1(n4408), .A2(n4407), .ZN(n440) );
  BUF_X4 U2156 ( .A(n3106), .Z(n3107) );
  BUF_X4 U2157 ( .A(n3106), .Z(n3108) );
  BUF_X4 U2158 ( .A(n3106), .Z(n3109) );
  BUF_X4 U2159 ( .A(N10), .Z(n3154) );
  BUF_X4 U2160 ( .A(n3105), .Z(n3110) );
  BUF_X4 U2161 ( .A(n3105), .Z(n3111) );
  BUF_X4 U2162 ( .A(N10), .Z(n3155) );
  BUF_X4 U2163 ( .A(n3105), .Z(n3112) );
  BUF_X4 U2164 ( .A(n3104), .Z(n3113) );
  BUF_X4 U2165 ( .A(N10), .Z(n3156) );
  BUF_X4 U2166 ( .A(n3104), .Z(n3114) );
  BUF_X4 U2167 ( .A(n3104), .Z(n3115) );
  BUF_X4 U2168 ( .A(N10), .Z(n3157) );
  BUF_X4 U2169 ( .A(n3103), .Z(n3116) );
  BUF_X4 U2170 ( .A(n3103), .Z(n3117) );
  BUF_X4 U2171 ( .A(N10), .Z(n3158) );
  BUF_X4 U2172 ( .A(n3103), .Z(n3118) );
  BUF_X4 U2173 ( .A(n3102), .Z(n3119) );
  BUF_X4 U2174 ( .A(N10), .Z(n3159) );
  BUF_X4 U2175 ( .A(n3102), .Z(n3120) );
  BUF_X4 U2176 ( .A(n3102), .Z(n3121) );
  BUF_X4 U2177 ( .A(N10), .Z(n3160) );
  BUF_X4 U2178 ( .A(n3101), .Z(n3122) );
  BUF_X4 U2179 ( .A(n3101), .Z(n3123) );
  BUF_X4 U2180 ( .A(N10), .Z(n3161) );
  BUF_X4 U2181 ( .A(n3101), .Z(n3124) );
  BUF_X4 U2182 ( .A(n3100), .Z(n3125) );
  BUF_X4 U2183 ( .A(N10), .Z(n3162) );
  BUF_X4 U2184 ( .A(n3100), .Z(n3126) );
  BUF_X4 U2185 ( .A(n3100), .Z(n3127) );
  BUF_X4 U2186 ( .A(N10), .Z(n3163) );
  BUF_X4 U2187 ( .A(n3099), .Z(n3128) );
  BUF_X4 U2188 ( .A(n3099), .Z(n3129) );
  BUF_X4 U2189 ( .A(N10), .Z(n3164) );
  BUF_X4 U2190 ( .A(n3099), .Z(n3130) );
  BUF_X4 U2191 ( .A(n3098), .Z(n3131) );
  BUF_X4 U2192 ( .A(N10), .Z(n3165) );
  BUF_X4 U2193 ( .A(n3098), .Z(n3132) );
  BUF_X4 U2194 ( .A(n3098), .Z(n3133) );
  BUF_X4 U2195 ( .A(N10), .Z(n3166) );
  BUF_X4 U2196 ( .A(n3097), .Z(n3134) );
  BUF_X4 U2197 ( .A(n3097), .Z(n3135) );
  BUF_X4 U2198 ( .A(N10), .Z(n3167) );
  BUF_X4 U2199 ( .A(n3097), .Z(n3136) );
  BUF_X4 U2200 ( .A(n3152), .Z(n3137) );
  BUF_X4 U2201 ( .A(N10), .Z(n3168) );
  BUF_X4 U2202 ( .A(n3152), .Z(n3138) );
  BUF_X4 U2203 ( .A(n3152), .Z(n3139) );
  BUF_X4 U2204 ( .A(N10), .Z(n3169) );
  BUF_X4 U2205 ( .A(n3152), .Z(n3140) );
  BUF_X4 U2206 ( .A(n3152), .Z(n3141) );
  BUF_X4 U2207 ( .A(N10), .Z(n3170) );
  BUF_X4 U2208 ( .A(n3152), .Z(n3142) );
  BUF_X4 U2209 ( .A(n3152), .Z(n3143) );
  BUF_X4 U2210 ( .A(N10), .Z(n3171) );
  BUF_X4 U2211 ( .A(n3152), .Z(n3144) );
  BUF_X4 U2212 ( .A(n3152), .Z(n3145) );
  BUF_X4 U2213 ( .A(n3152), .Z(n3146) );
  BUF_X4 U2214 ( .A(n3152), .Z(n3147) );
  BUF_X4 U2215 ( .A(n3152), .Z(n3148) );
  BUF_X4 U2216 ( .A(N9), .Z(n3149) );
  BUF_X4 U2217 ( .A(n3152), .Z(n3150) );
  BUF_X4 U2218 ( .A(N9), .Z(n3151) );
  BUF_X4 U2219 ( .A(N9), .Z(n3153) );
  INV_X4 U2220 ( .A(n3172), .ZN(n3181) );
  INV_X4 U2221 ( .A(n3172), .ZN(n3182) );
  OAI21_X2 U2222 ( .B1(n3252), .B2(n3254), .A(n1111), .ZN(n1113) );
  OAI21_X2 U2223 ( .B1(n3250), .B2(n3255), .A(n1100), .ZN(n1114) );
  OAI21_X2 U2224 ( .B1(n3248), .B2(n3255), .A(n1089), .ZN(n1115) );
  OAI21_X2 U2225 ( .B1(n3246), .B2(n3254), .A(n1086), .ZN(n1116) );
  OAI21_X2 U2226 ( .B1(n3244), .B2(n3254), .A(n1085), .ZN(n1117) );
  OAI21_X2 U2227 ( .B1(n3242), .B2(n3254), .A(n1084), .ZN(n1118) );
  OAI21_X2 U2228 ( .B1(n3240), .B2(n3254), .A(n1083), .ZN(n1119) );
  OAI21_X2 U2229 ( .B1(n3238), .B2(n3254), .A(n1082), .ZN(n1120) );
  OAI21_X2 U2230 ( .B1(n3236), .B2(n3254), .A(n1081), .ZN(n1121) );
  OAI21_X2 U2231 ( .B1(n3234), .B2(n3254), .A(n1080), .ZN(n1122) );
  OAI21_X2 U2232 ( .B1(n3232), .B2(n3254), .A(n1110), .ZN(n1123) );
  OAI21_X2 U2233 ( .B1(n3230), .B2(n3254), .A(n1109), .ZN(n1124) );
  OAI21_X2 U2234 ( .B1(n3228), .B2(n3254), .A(n1108), .ZN(n1125) );
  OAI21_X2 U2235 ( .B1(n3226), .B2(n3255), .A(n1107), .ZN(n1126) );
  OAI21_X2 U2236 ( .B1(n3224), .B2(n3255), .A(n1106), .ZN(n1127) );
  OAI21_X2 U2237 ( .B1(n3222), .B2(n3255), .A(n1105), .ZN(n1128) );
  OAI21_X2 U2238 ( .B1(n3220), .B2(n1079), .A(n1104), .ZN(n1129) );
  OAI21_X2 U2239 ( .B1(n3218), .B2(n3256), .A(n1103), .ZN(n1130) );
  OAI21_X2 U2240 ( .B1(n3216), .B2(n1079), .A(n1102), .ZN(n1131) );
  OAI21_X2 U2241 ( .B1(n3214), .B2(n1079), .A(n1101), .ZN(n1132) );
  OAI21_X2 U2242 ( .B1(n3212), .B2(n3254), .A(n1099), .ZN(n1133) );
  OAI21_X2 U2243 ( .B1(n3210), .B2(n3255), .A(n1098), .ZN(n1134) );
  OAI21_X2 U2244 ( .B1(n3208), .B2(n1079), .A(n1097), .ZN(n1135) );
  OAI21_X2 U2245 ( .B1(n3206), .B2(n1079), .A(n1096), .ZN(n1136) );
  OAI21_X2 U2246 ( .B1(n3204), .B2(n3255), .A(n1095), .ZN(n1137) );
  OAI21_X2 U2247 ( .B1(n3202), .B2(n3255), .A(n1094), .ZN(n1138) );
  OAI21_X2 U2248 ( .B1(n3200), .B2(n3255), .A(n1093), .ZN(n1139) );
  OAI21_X2 U2249 ( .B1(n3198), .B2(n3255), .A(n1092), .ZN(n1140) );
  OAI21_X2 U2250 ( .B1(n3196), .B2(n3255), .A(n1091), .ZN(n1141) );
  OAI21_X2 U2251 ( .B1(n3194), .B2(n3255), .A(n1090), .ZN(n1142) );
  OAI21_X2 U2252 ( .B1(n3192), .B2(n3255), .A(n1088), .ZN(n1143) );
  OAI21_X2 U2253 ( .B1(n3190), .B2(n3254), .A(n1087), .ZN(n1144) );
  OAI21_X2 U2254 ( .B1(n3252), .B2(n3298), .A(n741), .ZN(n1145) );
  OAI21_X2 U2255 ( .B1(n3250), .B2(n3299), .A(n730), .ZN(n1146) );
  OAI21_X2 U2256 ( .B1(n3248), .B2(n3299), .A(n719), .ZN(n1147) );
  OAI21_X2 U2257 ( .B1(n3246), .B2(n3298), .A(n716), .ZN(n1148) );
  OAI21_X2 U2258 ( .B1(n3244), .B2(n3298), .A(n715), .ZN(n1149) );
  OAI21_X2 U2259 ( .B1(n3242), .B2(n3298), .A(n714), .ZN(n1150) );
  OAI21_X2 U2260 ( .B1(n3240), .B2(n3298), .A(n713), .ZN(n1151) );
  OAI21_X2 U2261 ( .B1(n3238), .B2(n3298), .A(n712), .ZN(n1152) );
  OAI21_X2 U2262 ( .B1(n3236), .B2(n3298), .A(n711), .ZN(n1153) );
  OAI21_X2 U2263 ( .B1(n3234), .B2(n3298), .A(n710), .ZN(n1154) );
  OAI21_X2 U2264 ( .B1(n3232), .B2(n3298), .A(n740), .ZN(n1155) );
  OAI21_X2 U2265 ( .B1(n3230), .B2(n3298), .A(n739), .ZN(n1156) );
  OAI21_X2 U2266 ( .B1(n3228), .B2(n3298), .A(n738), .ZN(n1157) );
  OAI21_X2 U2267 ( .B1(n3226), .B2(n3299), .A(n737), .ZN(n1158) );
  OAI21_X2 U2268 ( .B1(n3224), .B2(n3299), .A(n736), .ZN(n1159) );
  OAI21_X2 U2269 ( .B1(n3222), .B2(n3299), .A(n735), .ZN(n1160) );
  OAI21_X2 U2270 ( .B1(n3220), .B2(n709), .A(n734), .ZN(n1161) );
  OAI21_X2 U2271 ( .B1(n3218), .B2(n3300), .A(n733), .ZN(n1162) );
  OAI21_X2 U2272 ( .B1(n3216), .B2(n709), .A(n732), .ZN(n1163) );
  OAI21_X2 U2273 ( .B1(n3214), .B2(n709), .A(n731), .ZN(n1164) );
  OAI21_X2 U2274 ( .B1(n3212), .B2(n3298), .A(n729), .ZN(n1165) );
  OAI21_X2 U2275 ( .B1(n3210), .B2(n3299), .A(n728), .ZN(n1166) );
  OAI21_X2 U2276 ( .B1(n3208), .B2(n709), .A(n727), .ZN(n1167) );
  OAI21_X2 U2277 ( .B1(n3206), .B2(n709), .A(n726), .ZN(n1168) );
  OAI21_X2 U2278 ( .B1(n3204), .B2(n3299), .A(n725), .ZN(n1169) );
  OAI21_X2 U2279 ( .B1(n3202), .B2(n3299), .A(n724), .ZN(n1170) );
  OAI21_X2 U2280 ( .B1(n3200), .B2(n3299), .A(n723), .ZN(n1171) );
  OAI21_X2 U2281 ( .B1(n3198), .B2(n3299), .A(n722), .ZN(n1172) );
  OAI21_X2 U2282 ( .B1(n3196), .B2(n3299), .A(n721), .ZN(n1173) );
  OAI21_X2 U2283 ( .B1(n3194), .B2(n3299), .A(n720), .ZN(n1174) );
  OAI21_X2 U2284 ( .B1(n3192), .B2(n3299), .A(n718), .ZN(n1175) );
  OAI21_X2 U2285 ( .B1(n3190), .B2(n3298), .A(n717), .ZN(n1176) );
  OAI21_X2 U2286 ( .B1(n3253), .B2(n3343), .A(n372), .ZN(n1177) );
  OAI21_X2 U2287 ( .B1(n3251), .B2(n3343), .A(n361), .ZN(n1178) );
  OAI21_X2 U2288 ( .B1(n3249), .B2(n3344), .A(n350), .ZN(n1179) );
  OAI21_X2 U2289 ( .B1(n3247), .B2(n3343), .A(n347), .ZN(n1180) );
  OAI21_X2 U2290 ( .B1(n3245), .B2(n3343), .A(n346), .ZN(n1181) );
  OAI21_X2 U2291 ( .B1(n3243), .B2(n3343), .A(n345), .ZN(n1182) );
  OAI21_X2 U2292 ( .B1(n3241), .B2(n3343), .A(n344), .ZN(n1183) );
  OAI21_X2 U2293 ( .B1(n3239), .B2(n3343), .A(n343), .ZN(n1184) );
  OAI21_X2 U2294 ( .B1(n3237), .B2(n3343), .A(n342), .ZN(n1185) );
  OAI21_X2 U2295 ( .B1(n3235), .B2(n3343), .A(n341), .ZN(n1186) );
  OAI21_X2 U2296 ( .B1(n3233), .B2(n3343), .A(n371), .ZN(n1187) );
  OAI21_X2 U2297 ( .B1(n3231), .B2(n3343), .A(n370), .ZN(n1188) );
  OAI21_X2 U2298 ( .B1(n3229), .B2(n3343), .A(n369), .ZN(n1189) );
  OAI21_X2 U2299 ( .B1(n3227), .B2(n3344), .A(n368), .ZN(n1190) );
  OAI21_X2 U2300 ( .B1(n3225), .B2(n3344), .A(n367), .ZN(n1191) );
  OAI21_X2 U2301 ( .B1(n3223), .B2(n3344), .A(n366), .ZN(n1192) );
  OAI21_X2 U2302 ( .B1(n3221), .B2(n340), .A(n365), .ZN(n1193) );
  OAI21_X2 U2303 ( .B1(n3219), .B2(n3344), .A(n364), .ZN(n1194) );
  OAI21_X2 U2304 ( .B1(n3217), .B2(n340), .A(n363), .ZN(n1195) );
  OAI21_X2 U2305 ( .B1(n3215), .B2(n340), .A(n362), .ZN(n1196) );
  OAI21_X2 U2306 ( .B1(n3213), .B2(n3345), .A(n360), .ZN(n1197) );
  OAI21_X2 U2307 ( .B1(n3211), .B2(n3344), .A(n359), .ZN(n1198) );
  OAI21_X2 U2308 ( .B1(n3209), .B2(n340), .A(n358), .ZN(n1199) );
  OAI21_X2 U2309 ( .B1(n3207), .B2(n340), .A(n357), .ZN(n1200) );
  OAI21_X2 U2310 ( .B1(n3205), .B2(n3344), .A(n356), .ZN(n1201) );
  OAI21_X2 U2311 ( .B1(n3203), .B2(n3344), .A(n355), .ZN(n1202) );
  OAI21_X2 U2312 ( .B1(n3201), .B2(n3344), .A(n354), .ZN(n1203) );
  OAI21_X2 U2313 ( .B1(n3199), .B2(n3344), .A(n353), .ZN(n1204) );
  OAI21_X2 U2314 ( .B1(n3197), .B2(n3344), .A(n352), .ZN(n1205) );
  OAI21_X2 U2315 ( .B1(n3195), .B2(n3344), .A(n351), .ZN(n1206) );
  OAI21_X2 U2316 ( .B1(n3193), .B2(n3344), .A(n349), .ZN(n1207) );
  OAI21_X2 U2317 ( .B1(n3191), .B2(n3343), .A(n348), .ZN(n1208) );
  OAI21_X2 U2318 ( .B1(n3253), .B2(n3355), .A(n271), .ZN(n1209) );
  OAI21_X2 U2319 ( .B1(n3251), .B2(n3355), .A(n260), .ZN(n1210) );
  OAI21_X2 U2320 ( .B1(n3249), .B2(n3356), .A(n249), .ZN(n1211) );
  OAI21_X2 U2321 ( .B1(n3247), .B2(n3355), .A(n246), .ZN(n1212) );
  OAI21_X2 U2322 ( .B1(n3245), .B2(n3355), .A(n245), .ZN(n1213) );
  OAI21_X2 U2323 ( .B1(n3243), .B2(n3355), .A(n244), .ZN(n1214) );
  OAI21_X2 U2324 ( .B1(n3241), .B2(n3355), .A(n243), .ZN(n1215) );
  OAI21_X2 U2325 ( .B1(n3239), .B2(n3355), .A(n242), .ZN(n1216) );
  OAI21_X2 U2326 ( .B1(n3237), .B2(n3355), .A(n241), .ZN(n1217) );
  OAI21_X2 U2327 ( .B1(n3235), .B2(n3355), .A(n240), .ZN(n1218) );
  OAI21_X2 U2328 ( .B1(n3233), .B2(n3355), .A(n270), .ZN(n1219) );
  OAI21_X2 U2329 ( .B1(n3231), .B2(n3355), .A(n269), .ZN(n1220) );
  OAI21_X2 U2330 ( .B1(n3229), .B2(n3355), .A(n268), .ZN(n1221) );
  OAI21_X2 U2331 ( .B1(n3227), .B2(n3356), .A(n267), .ZN(n1222) );
  OAI21_X2 U2332 ( .B1(n3225), .B2(n3356), .A(n266), .ZN(n1223) );
  OAI21_X2 U2333 ( .B1(n3223), .B2(n3356), .A(n265), .ZN(n1224) );
  OAI21_X2 U2334 ( .B1(n3221), .B2(n239), .A(n264), .ZN(n1225) );
  OAI21_X2 U2335 ( .B1(n3219), .B2(n3356), .A(n263), .ZN(n1226) );
  OAI21_X2 U2336 ( .B1(n3217), .B2(n239), .A(n262), .ZN(n1227) );
  OAI21_X2 U2337 ( .B1(n3215), .B2(n239), .A(n261), .ZN(n1228) );
  OAI21_X2 U2338 ( .B1(n3213), .B2(n3357), .A(n259), .ZN(n1229) );
  OAI21_X2 U2339 ( .B1(n3211), .B2(n3356), .A(n258), .ZN(n1230) );
  OAI21_X2 U2340 ( .B1(n3209), .B2(n239), .A(n257), .ZN(n1231) );
  OAI21_X2 U2341 ( .B1(n3207), .B2(n239), .A(n256), .ZN(n1232) );
  OAI21_X2 U2342 ( .B1(n3205), .B2(n3356), .A(n255), .ZN(n1233) );
  OAI21_X2 U2343 ( .B1(n3203), .B2(n3356), .A(n254), .ZN(n1234) );
  OAI21_X2 U2344 ( .B1(n3201), .B2(n3356), .A(n253), .ZN(n1235) );
  OAI21_X2 U2345 ( .B1(n3199), .B2(n3356), .A(n252), .ZN(n1236) );
  OAI21_X2 U2346 ( .B1(n3197), .B2(n3356), .A(n251), .ZN(n1237) );
  OAI21_X2 U2347 ( .B1(n3195), .B2(n3356), .A(n250), .ZN(n1238) );
  OAI21_X2 U2348 ( .B1(n3193), .B2(n3356), .A(n248), .ZN(n1239) );
  OAI21_X2 U2349 ( .B1(n3191), .B2(n3355), .A(n247), .ZN(n1240) );
  OAI21_X2 U2350 ( .B1(n3253), .B2(n3358), .A(n236), .ZN(n1241) );
  OAI21_X2 U2351 ( .B1(n3251), .B2(n3359), .A(n225), .ZN(n1242) );
  OAI21_X2 U2352 ( .B1(n3249), .B2(n3359), .A(n214), .ZN(n1243) );
  OAI21_X2 U2353 ( .B1(n3247), .B2(n3358), .A(n211), .ZN(n1244) );
  OAI21_X2 U2354 ( .B1(n3245), .B2(n3358), .A(n210), .ZN(n1245) );
  OAI21_X2 U2355 ( .B1(n3243), .B2(n3358), .A(n209), .ZN(n1246) );
  OAI21_X2 U2356 ( .B1(n3241), .B2(n3358), .A(n208), .ZN(n1247) );
  OAI21_X2 U2357 ( .B1(n3239), .B2(n3358), .A(n207), .ZN(n1248) );
  OAI21_X2 U2358 ( .B1(n3237), .B2(n3358), .A(n206), .ZN(n1249) );
  OAI21_X2 U2359 ( .B1(n3235), .B2(n3358), .A(n205), .ZN(n1250) );
  OAI21_X2 U2360 ( .B1(n3233), .B2(n3358), .A(n235), .ZN(n1251) );
  OAI21_X2 U2361 ( .B1(n3231), .B2(n3358), .A(n234), .ZN(n1252) );
  OAI21_X2 U2362 ( .B1(n3229), .B2(n3358), .A(n233), .ZN(n1253) );
  OAI21_X2 U2363 ( .B1(n3227), .B2(n3359), .A(n232), .ZN(n1254) );
  OAI21_X2 U2364 ( .B1(n3225), .B2(n3359), .A(n231), .ZN(n1255) );
  OAI21_X2 U2365 ( .B1(n3223), .B2(n3359), .A(n230), .ZN(n1256) );
  OAI21_X2 U2366 ( .B1(n3221), .B2(n204), .A(n229), .ZN(n1257) );
  OAI21_X2 U2367 ( .B1(n3219), .B2(n3360), .A(n228), .ZN(n1258) );
  OAI21_X2 U2368 ( .B1(n3217), .B2(n204), .A(n227), .ZN(n1259) );
  OAI21_X2 U2369 ( .B1(n3215), .B2(n204), .A(n226), .ZN(n1260) );
  OAI21_X2 U2370 ( .B1(n3213), .B2(n3358), .A(n224), .ZN(n1261) );
  OAI21_X2 U2371 ( .B1(n3211), .B2(n3359), .A(n223), .ZN(n1262) );
  OAI21_X2 U2372 ( .B1(n3209), .B2(n204), .A(n222), .ZN(n1263) );
  OAI21_X2 U2373 ( .B1(n3207), .B2(n204), .A(n221), .ZN(n1264) );
  OAI21_X2 U2374 ( .B1(n3205), .B2(n3359), .A(n220), .ZN(n1265) );
  OAI21_X2 U2375 ( .B1(n3203), .B2(n3359), .A(n219), .ZN(n1266) );
  OAI21_X2 U2376 ( .B1(n3201), .B2(n3359), .A(n218), .ZN(n1267) );
  OAI21_X2 U2377 ( .B1(n3199), .B2(n3359), .A(n217), .ZN(n1268) );
  OAI21_X2 U2378 ( .B1(n3197), .B2(n3359), .A(n216), .ZN(n1269) );
  OAI21_X2 U2379 ( .B1(n3195), .B2(n3359), .A(n215), .ZN(n1270) );
  OAI21_X2 U2380 ( .B1(n3193), .B2(n3359), .A(n213), .ZN(n1271) );
  OAI21_X2 U2381 ( .B1(n3191), .B2(n3358), .A(n212), .ZN(n1272) );
  OAI21_X2 U2382 ( .B1(n3253), .B2(n3362), .A(n203), .ZN(n1273) );
  OAI21_X2 U2383 ( .B1(n3251), .B2(n3363), .A(n192), .ZN(n1274) );
  OAI21_X2 U2384 ( .B1(n3249), .B2(n3363), .A(n181), .ZN(n1275) );
  OAI21_X2 U2385 ( .B1(n3247), .B2(n3362), .A(n178), .ZN(n1276) );
  OAI21_X2 U2386 ( .B1(n3245), .B2(n3362), .A(n177), .ZN(n1277) );
  OAI21_X2 U2387 ( .B1(n3243), .B2(n3362), .A(n176), .ZN(n1278) );
  OAI21_X2 U2388 ( .B1(n3241), .B2(n3362), .A(n175), .ZN(n1279) );
  OAI21_X2 U2389 ( .B1(n3239), .B2(n3362), .A(n174), .ZN(n1280) );
  OAI21_X2 U2390 ( .B1(n3237), .B2(n3362), .A(n173), .ZN(n1281) );
  OAI21_X2 U2391 ( .B1(n3235), .B2(n3362), .A(n172), .ZN(n1282) );
  OAI21_X2 U2392 ( .B1(n3233), .B2(n3362), .A(n202), .ZN(n1283) );
  OAI21_X2 U2393 ( .B1(n3231), .B2(n3362), .A(n201), .ZN(n1284) );
  OAI21_X2 U2394 ( .B1(n3229), .B2(n3362), .A(n200), .ZN(n1285) );
  OAI21_X2 U2395 ( .B1(n3227), .B2(n3363), .A(n199), .ZN(n1286) );
  OAI21_X2 U2396 ( .B1(n3225), .B2(n3363), .A(n198), .ZN(n1287) );
  OAI21_X2 U2397 ( .B1(n3223), .B2(n3363), .A(n197), .ZN(n1288) );
  OAI21_X2 U2398 ( .B1(n3221), .B2(n171), .A(n196), .ZN(n1289) );
  OAI21_X2 U2399 ( .B1(n3219), .B2(n3364), .A(n195), .ZN(n1290) );
  OAI21_X2 U2400 ( .B1(n3217), .B2(n171), .A(n194), .ZN(n1291) );
  OAI21_X2 U2401 ( .B1(n3215), .B2(n171), .A(n193), .ZN(n1292) );
  OAI21_X2 U2402 ( .B1(n3213), .B2(n3362), .A(n191), .ZN(n1293) );
  OAI21_X2 U2403 ( .B1(n3211), .B2(n3363), .A(n190), .ZN(n1294) );
  OAI21_X2 U2404 ( .B1(n3209), .B2(n171), .A(n189), .ZN(n1295) );
  OAI21_X2 U2405 ( .B1(n3207), .B2(n171), .A(n188), .ZN(n1296) );
  OAI21_X2 U2406 ( .B1(n3205), .B2(n3363), .A(n187), .ZN(n1297) );
  OAI21_X2 U2407 ( .B1(n3203), .B2(n3363), .A(n186), .ZN(n1298) );
  OAI21_X2 U2408 ( .B1(n3201), .B2(n3363), .A(n185), .ZN(n1299) );
  OAI21_X2 U2409 ( .B1(n3199), .B2(n3363), .A(n184), .ZN(n1300) );
  OAI21_X2 U2410 ( .B1(n3197), .B2(n3363), .A(n183), .ZN(n1301) );
  OAI21_X2 U2411 ( .B1(n3195), .B2(n3363), .A(n182), .ZN(n1302) );
  OAI21_X2 U2412 ( .B1(n3193), .B2(n3363), .A(n180), .ZN(n1303) );
  OAI21_X2 U2413 ( .B1(n3191), .B2(n3362), .A(n179), .ZN(n1304) );
  OAI21_X2 U2414 ( .B1(n3252), .B2(n3367), .A(n169), .ZN(n1305) );
  OAI21_X2 U2415 ( .B1(n3250), .B2(n3367), .A(n158), .ZN(n1306) );
  OAI21_X2 U2416 ( .B1(n3248), .B2(n3368), .A(n147), .ZN(n1307) );
  OAI21_X2 U2417 ( .B1(n3246), .B2(n3367), .A(n144), .ZN(n1308) );
  OAI21_X2 U2418 ( .B1(n3244), .B2(n3367), .A(n143), .ZN(n1309) );
  OAI21_X2 U2419 ( .B1(n3242), .B2(n3367), .A(n142), .ZN(n1310) );
  OAI21_X2 U2420 ( .B1(n3240), .B2(n3367), .A(n141), .ZN(n1311) );
  OAI21_X2 U2421 ( .B1(n3238), .B2(n3367), .A(n140), .ZN(n1312) );
  OAI21_X2 U2422 ( .B1(n3236), .B2(n3367), .A(n139), .ZN(n1313) );
  OAI21_X2 U2423 ( .B1(n3234), .B2(n3367), .A(n138), .ZN(n1314) );
  OAI21_X2 U2424 ( .B1(n3232), .B2(n3367), .A(n168), .ZN(n1315) );
  OAI21_X2 U2425 ( .B1(n3230), .B2(n3367), .A(n167), .ZN(n1316) );
  OAI21_X2 U2426 ( .B1(n3228), .B2(n3367), .A(n166), .ZN(n1317) );
  OAI21_X2 U2427 ( .B1(n3226), .B2(n3368), .A(n165), .ZN(n1318) );
  OAI21_X2 U2428 ( .B1(n3224), .B2(n3368), .A(n164), .ZN(n1319) );
  OAI21_X2 U2429 ( .B1(n3222), .B2(n3368), .A(n163), .ZN(n1320) );
  OAI21_X2 U2430 ( .B1(n3220), .B2(n137), .A(n162), .ZN(n1321) );
  OAI21_X2 U2431 ( .B1(n3218), .B2(n3368), .A(n161), .ZN(n1322) );
  OAI21_X2 U2432 ( .B1(n3216), .B2(n137), .A(n160), .ZN(n1323) );
  OAI21_X2 U2433 ( .B1(n3214), .B2(n137), .A(n159), .ZN(n1324) );
  OAI21_X2 U2434 ( .B1(n3212), .B2(n3369), .A(n157), .ZN(n1325) );
  OAI21_X2 U2435 ( .B1(n3210), .B2(n3368), .A(n156), .ZN(n1326) );
  OAI21_X2 U2436 ( .B1(n3208), .B2(n137), .A(n155), .ZN(n1327) );
  OAI21_X2 U2437 ( .B1(n3206), .B2(n137), .A(n154), .ZN(n1328) );
  OAI21_X2 U2438 ( .B1(n3204), .B2(n3368), .A(n153), .ZN(n1329) );
  OAI21_X2 U2439 ( .B1(n3202), .B2(n3368), .A(n152), .ZN(n1330) );
  OAI21_X2 U2440 ( .B1(n3200), .B2(n3368), .A(n151), .ZN(n1331) );
  OAI21_X2 U2441 ( .B1(n3198), .B2(n3368), .A(n150), .ZN(n1332) );
  OAI21_X2 U2442 ( .B1(n3196), .B2(n3368), .A(n149), .ZN(n1333) );
  OAI21_X2 U2443 ( .B1(n3194), .B2(n3368), .A(n148), .ZN(n1334) );
  OAI21_X2 U2444 ( .B1(n3192), .B2(n3368), .A(n146), .ZN(n1335) );
  OAI21_X2 U2445 ( .B1(n3190), .B2(n3367), .A(n145), .ZN(n1336) );
  OAI21_X2 U2446 ( .B1(n3253), .B2(n3371), .A(n134), .ZN(n1337) );
  OAI21_X2 U2447 ( .B1(n3251), .B2(n3371), .A(n123), .ZN(n1338) );
  OAI21_X2 U2448 ( .B1(n3249), .B2(n3372), .A(n112), .ZN(n1339) );
  OAI21_X2 U2449 ( .B1(n3247), .B2(n3371), .A(n109), .ZN(n1340) );
  OAI21_X2 U2450 ( .B1(n3245), .B2(n3371), .A(n108), .ZN(n1341) );
  OAI21_X2 U2451 ( .B1(n3243), .B2(n3371), .A(n107), .ZN(n1342) );
  OAI21_X2 U2452 ( .B1(n3241), .B2(n3371), .A(n106), .ZN(n1343) );
  OAI21_X2 U2453 ( .B1(n3239), .B2(n3371), .A(n105), .ZN(n1344) );
  OAI21_X2 U2454 ( .B1(n3237), .B2(n3371), .A(n104), .ZN(n1345) );
  OAI21_X2 U2455 ( .B1(n3235), .B2(n3371), .A(n103), .ZN(n1346) );
  OAI21_X2 U2456 ( .B1(n3233), .B2(n3371), .A(n133), .ZN(n1347) );
  OAI21_X2 U2457 ( .B1(n3231), .B2(n3371), .A(n132), .ZN(n1348) );
  OAI21_X2 U2458 ( .B1(n3229), .B2(n3371), .A(n131), .ZN(n1349) );
  OAI21_X2 U2459 ( .B1(n3227), .B2(n3372), .A(n130), .ZN(n1350) );
  OAI21_X2 U2460 ( .B1(n3225), .B2(n3372), .A(n129), .ZN(n1351) );
  OAI21_X2 U2461 ( .B1(n3223), .B2(n3372), .A(n128), .ZN(n1352) );
  OAI21_X2 U2462 ( .B1(n3221), .B2(n102), .A(n127), .ZN(n1353) );
  OAI21_X2 U2463 ( .B1(n3219), .B2(n3372), .A(n126), .ZN(n1354) );
  OAI21_X2 U2464 ( .B1(n3217), .B2(n102), .A(n125), .ZN(n1355) );
  OAI21_X2 U2465 ( .B1(n3215), .B2(n102), .A(n124), .ZN(n1356) );
  OAI21_X2 U2466 ( .B1(n3213), .B2(n3373), .A(n122), .ZN(n1357) );
  OAI21_X2 U2467 ( .B1(n3211), .B2(n3372), .A(n121), .ZN(n1358) );
  OAI21_X2 U2468 ( .B1(n3209), .B2(n102), .A(n120), .ZN(n1359) );
  OAI21_X2 U2469 ( .B1(n3207), .B2(n102), .A(n119), .ZN(n1360) );
  OAI21_X2 U2470 ( .B1(n3205), .B2(n3372), .A(n118), .ZN(n1361) );
  OAI21_X2 U2471 ( .B1(n3203), .B2(n3372), .A(n117), .ZN(n1362) );
  OAI21_X2 U2472 ( .B1(n3201), .B2(n3372), .A(n116), .ZN(n1363) );
  OAI21_X2 U2473 ( .B1(n3199), .B2(n3372), .A(n115), .ZN(n1364) );
  OAI21_X2 U2474 ( .B1(n3197), .B2(n3372), .A(n114), .ZN(n1365) );
  OAI21_X2 U2475 ( .B1(n3195), .B2(n3372), .A(n113), .ZN(n1366) );
  OAI21_X2 U2476 ( .B1(n3193), .B2(n3372), .A(n111), .ZN(n1367) );
  OAI21_X2 U2477 ( .B1(n3191), .B2(n3371), .A(n110), .ZN(n1368) );
  OAI21_X2 U2478 ( .B1(n3253), .B2(n3375), .A(n100), .ZN(n1369) );
  OAI21_X2 U2479 ( .B1(n3251), .B2(n3375), .A(n89), .ZN(n1370) );
  OAI21_X2 U2480 ( .B1(n3249), .B2(n3376), .A(n78), .ZN(n1371) );
  OAI21_X2 U2481 ( .B1(n3247), .B2(n3375), .A(n75), .ZN(n1372) );
  OAI21_X2 U2482 ( .B1(n3245), .B2(n3375), .A(n74), .ZN(n1373) );
  OAI21_X2 U2483 ( .B1(n3243), .B2(n3375), .A(n73), .ZN(n1374) );
  OAI21_X2 U2484 ( .B1(n3241), .B2(n3375), .A(n72), .ZN(n1375) );
  OAI21_X2 U2485 ( .B1(n3239), .B2(n3375), .A(n71), .ZN(n1376) );
  OAI21_X2 U2486 ( .B1(n3237), .B2(n3375), .A(n70), .ZN(n1377) );
  OAI21_X2 U2487 ( .B1(n3235), .B2(n3375), .A(n69), .ZN(n1378) );
  OAI21_X2 U2488 ( .B1(n3233), .B2(n3375), .A(n99), .ZN(n1379) );
  OAI21_X2 U2489 ( .B1(n3231), .B2(n3375), .A(n98), .ZN(n1380) );
  OAI21_X2 U2490 ( .B1(n3229), .B2(n3375), .A(n97), .ZN(n1381) );
  OAI21_X2 U2491 ( .B1(n3227), .B2(n3376), .A(n96), .ZN(n1382) );
  OAI21_X2 U2492 ( .B1(n3225), .B2(n3376), .A(n95), .ZN(n1383) );
  OAI21_X2 U2493 ( .B1(n3223), .B2(n3376), .A(n94), .ZN(n1384) );
  OAI21_X2 U2494 ( .B1(n3221), .B2(n68), .A(n93), .ZN(n1385) );
  OAI21_X2 U2495 ( .B1(n3219), .B2(n3376), .A(n92), .ZN(n1386) );
  OAI21_X2 U2496 ( .B1(n3217), .B2(n68), .A(n91), .ZN(n1387) );
  OAI21_X2 U2497 ( .B1(n3215), .B2(n68), .A(n90), .ZN(n1388) );
  OAI21_X2 U2498 ( .B1(n3213), .B2(n3377), .A(n88), .ZN(n1389) );
  OAI21_X2 U2499 ( .B1(n3211), .B2(n3376), .A(n87), .ZN(n1390) );
  OAI21_X2 U2500 ( .B1(n3209), .B2(n68), .A(n86), .ZN(n1391) );
  OAI21_X2 U2501 ( .B1(n3207), .B2(n68), .A(n85), .ZN(n1392) );
  OAI21_X2 U2502 ( .B1(n3205), .B2(n3376), .A(n84), .ZN(n1393) );
  OAI21_X2 U2503 ( .B1(n3203), .B2(n3376), .A(n83), .ZN(n1394) );
  OAI21_X2 U2504 ( .B1(n3201), .B2(n3376), .A(n82), .ZN(n1395) );
  OAI21_X2 U2505 ( .B1(n3199), .B2(n3376), .A(n81), .ZN(n1396) );
  OAI21_X2 U2506 ( .B1(n3197), .B2(n3376), .A(n80), .ZN(n1397) );
  OAI21_X2 U2507 ( .B1(n3195), .B2(n3376), .A(n79), .ZN(n1398) );
  OAI21_X2 U2508 ( .B1(n3193), .B2(n3376), .A(n77), .ZN(n1399) );
  OAI21_X2 U2509 ( .B1(n3191), .B2(n3375), .A(n76), .ZN(n1400) );
  OAI21_X2 U2510 ( .B1(n3379), .B2(n3252), .A(n65), .ZN(n1401) );
  OAI21_X2 U2511 ( .B1(n3379), .B2(n3250), .A(n43), .ZN(n1402) );
  OAI21_X2 U2512 ( .B1(n3380), .B2(n3248), .A(n21), .ZN(n1403) );
  OAI21_X2 U2513 ( .B1(n3379), .B2(n3246), .A(n15), .ZN(n1404) );
  OAI21_X2 U2514 ( .B1(n3379), .B2(n3244), .A(n13), .ZN(n1405) );
  OAI21_X2 U2515 ( .B1(n3379), .B2(n3242), .A(n11), .ZN(n1406) );
  OAI21_X2 U2516 ( .B1(n3379), .B2(n3240), .A(n9), .ZN(n1407) );
  OAI21_X2 U2517 ( .B1(n3379), .B2(n3238), .A(n7), .ZN(n1408) );
  OAI21_X2 U2518 ( .B1(n3379), .B2(n3236), .A(n5), .ZN(n1409) );
  OAI21_X2 U2519 ( .B1(n3379), .B2(n3234), .A(n3), .ZN(n1410) );
  OAI21_X2 U2520 ( .B1(n3379), .B2(n3232), .A(n63), .ZN(n1411) );
  OAI21_X2 U2521 ( .B1(n3379), .B2(n3230), .A(n61), .ZN(n1412) );
  OAI21_X2 U2522 ( .B1(n3379), .B2(n3228), .A(n59), .ZN(n1413) );
  OAI21_X2 U2523 ( .B1(n3380), .B2(n3226), .A(n57), .ZN(n1414) );
  OAI21_X2 U2524 ( .B1(n3380), .B2(n3224), .A(n55), .ZN(n1415) );
  OAI21_X2 U2525 ( .B1(n3380), .B2(n3222), .A(n53), .ZN(n1416) );
  OAI21_X2 U2526 ( .B1(n1), .B2(n3220), .A(n51), .ZN(n1417) );
  OAI21_X2 U2527 ( .B1(n3380), .B2(n3218), .A(n49), .ZN(n1418) );
  OAI21_X2 U2528 ( .B1(n1), .B2(n3216), .A(n47), .ZN(n1419) );
  OAI21_X2 U2529 ( .B1(n1), .B2(n3214), .A(n45), .ZN(n1420) );
  OAI21_X2 U2530 ( .B1(n3381), .B2(n3212), .A(n41), .ZN(n1421) );
  OAI21_X2 U2531 ( .B1(n3380), .B2(n3210), .A(n39), .ZN(n1422) );
  OAI21_X2 U2532 ( .B1(n1), .B2(n3208), .A(n37), .ZN(n1423) );
  OAI21_X2 U2533 ( .B1(n1), .B2(n3206), .A(n35), .ZN(n1424) );
  OAI21_X2 U2534 ( .B1(n3380), .B2(n3204), .A(n33), .ZN(n1425) );
  OAI21_X2 U2535 ( .B1(n3380), .B2(n3202), .A(n31), .ZN(n1426) );
  OAI21_X2 U2536 ( .B1(n3380), .B2(n3200), .A(n29), .ZN(n1427) );
  OAI21_X2 U2537 ( .B1(n3380), .B2(n3198), .A(n27), .ZN(n1428) );
  OAI21_X2 U2538 ( .B1(n3380), .B2(n3196), .A(n25), .ZN(n1429) );
  OAI21_X2 U2539 ( .B1(n3380), .B2(n3194), .A(n23), .ZN(n1430) );
  OAI21_X2 U2540 ( .B1(n3380), .B2(n3192), .A(n19), .ZN(n1431) );
  OAI21_X2 U2541 ( .B1(n3379), .B2(n3190), .A(n17), .ZN(n1432) );
  OAI21_X2 U2542 ( .B1(n3252), .B2(n3259), .A(n1078), .ZN(n1433) );
  OAI21_X2 U2543 ( .B1(n3250), .B2(n3259), .A(n1067), .ZN(n1434) );
  OAI21_X2 U2544 ( .B1(n3248), .B2(n3260), .A(n1056), .ZN(n1435) );
  OAI21_X2 U2545 ( .B1(n3246), .B2(n3259), .A(n1053), .ZN(n1436) );
  OAI21_X2 U2546 ( .B1(n3244), .B2(n3259), .A(n1052), .ZN(n1437) );
  OAI21_X2 U2547 ( .B1(n3242), .B2(n3259), .A(n1051), .ZN(n1438) );
  OAI21_X2 U2548 ( .B1(n3240), .B2(n3259), .A(n1050), .ZN(n1439) );
  OAI21_X2 U2549 ( .B1(n3238), .B2(n3259), .A(n1049), .ZN(n1440) );
  OAI21_X2 U2550 ( .B1(n3236), .B2(n3259), .A(n1048), .ZN(n1441) );
  OAI21_X2 U2551 ( .B1(n3234), .B2(n3259), .A(n1047), .ZN(n1442) );
  OAI21_X2 U2552 ( .B1(n3232), .B2(n3259), .A(n1077), .ZN(n1443) );
  OAI21_X2 U2553 ( .B1(n3230), .B2(n3259), .A(n1076), .ZN(n1444) );
  OAI21_X2 U2554 ( .B1(n3228), .B2(n3259), .A(n1075), .ZN(n1445) );
  OAI21_X2 U2555 ( .B1(n3226), .B2(n3260), .A(n1074), .ZN(n1446) );
  OAI21_X2 U2556 ( .B1(n3224), .B2(n3260), .A(n1073), .ZN(n1447) );
  OAI21_X2 U2557 ( .B1(n3222), .B2(n3260), .A(n1072), .ZN(n1448) );
  OAI21_X2 U2558 ( .B1(n3220), .B2(n1046), .A(n1071), .ZN(n1449) );
  OAI21_X2 U2559 ( .B1(n3218), .B2(n3260), .A(n1070), .ZN(n1450) );
  OAI21_X2 U2560 ( .B1(n3216), .B2(n1046), .A(n1069), .ZN(n1451) );
  OAI21_X2 U2561 ( .B1(n3214), .B2(n1046), .A(n1068), .ZN(n1452) );
  OAI21_X2 U2562 ( .B1(n3212), .B2(n3261), .A(n1066), .ZN(n1453) );
  OAI21_X2 U2563 ( .B1(n3210), .B2(n3260), .A(n1065), .ZN(n1454) );
  OAI21_X2 U2564 ( .B1(n3208), .B2(n1046), .A(n1064), .ZN(n1455) );
  OAI21_X2 U2565 ( .B1(n3206), .B2(n1046), .A(n1063), .ZN(n1456) );
  OAI21_X2 U2566 ( .B1(n3204), .B2(n3260), .A(n1062), .ZN(n1457) );
  OAI21_X2 U2567 ( .B1(n3202), .B2(n3260), .A(n1061), .ZN(n1458) );
  OAI21_X2 U2568 ( .B1(n3200), .B2(n3260), .A(n1060), .ZN(n1459) );
  OAI21_X2 U2569 ( .B1(n3198), .B2(n3260), .A(n1059), .ZN(n1460) );
  OAI21_X2 U2570 ( .B1(n3196), .B2(n3260), .A(n1058), .ZN(n1461) );
  OAI21_X2 U2571 ( .B1(n3194), .B2(n3260), .A(n1057), .ZN(n1462) );
  OAI21_X2 U2572 ( .B1(n3192), .B2(n3260), .A(n1055), .ZN(n1463) );
  OAI21_X2 U2573 ( .B1(n3190), .B2(n3259), .A(n1054), .ZN(n1464) );
  OAI21_X2 U2574 ( .B1(n3252), .B2(n3263), .A(n1045), .ZN(n1465) );
  OAI21_X2 U2575 ( .B1(n3250), .B2(n3263), .A(n1034), .ZN(n1466) );
  OAI21_X2 U2576 ( .B1(n3248), .B2(n3264), .A(n1023), .ZN(n1467) );
  OAI21_X2 U2577 ( .B1(n3246), .B2(n3263), .A(n1020), .ZN(n1468) );
  OAI21_X2 U2578 ( .B1(n3244), .B2(n3263), .A(n1019), .ZN(n1469) );
  OAI21_X2 U2579 ( .B1(n3242), .B2(n3263), .A(n1018), .ZN(n1470) );
  OAI21_X2 U2580 ( .B1(n3240), .B2(n3263), .A(n1017), .ZN(n1471) );
  OAI21_X2 U2581 ( .B1(n3238), .B2(n3263), .A(n1016), .ZN(n1472) );
  OAI21_X2 U2582 ( .B1(n3236), .B2(n3263), .A(n1015), .ZN(n1473) );
  OAI21_X2 U2583 ( .B1(n3234), .B2(n3263), .A(n1014), .ZN(n1474) );
  OAI21_X2 U2584 ( .B1(n3232), .B2(n3263), .A(n1044), .ZN(n1475) );
  OAI21_X2 U2585 ( .B1(n3230), .B2(n3263), .A(n1043), .ZN(n1476) );
  OAI21_X2 U2586 ( .B1(n3228), .B2(n3263), .A(n1042), .ZN(n1477) );
  OAI21_X2 U2587 ( .B1(n3226), .B2(n3264), .A(n1041), .ZN(n1478) );
  OAI21_X2 U2588 ( .B1(n3224), .B2(n3264), .A(n1040), .ZN(n1479) );
  OAI21_X2 U2589 ( .B1(n3222), .B2(n3264), .A(n1039), .ZN(n1480) );
  OAI21_X2 U2590 ( .B1(n3220), .B2(n1013), .A(n1038), .ZN(n1481) );
  OAI21_X2 U2591 ( .B1(n3218), .B2(n3264), .A(n1037), .ZN(n1482) );
  OAI21_X2 U2592 ( .B1(n3216), .B2(n1013), .A(n1036), .ZN(n1483) );
  OAI21_X2 U2593 ( .B1(n3214), .B2(n1013), .A(n1035), .ZN(n1484) );
  OAI21_X2 U2594 ( .B1(n3212), .B2(n3265), .A(n1033), .ZN(n1485) );
  OAI21_X2 U2595 ( .B1(n3210), .B2(n3264), .A(n1032), .ZN(n1486) );
  OAI21_X2 U2596 ( .B1(n3208), .B2(n1013), .A(n1031), .ZN(n1487) );
  OAI21_X2 U2597 ( .B1(n3206), .B2(n1013), .A(n1030), .ZN(n1488) );
  OAI21_X2 U2598 ( .B1(n3204), .B2(n3264), .A(n1029), .ZN(n1489) );
  OAI21_X2 U2599 ( .B1(n3202), .B2(n3264), .A(n1028), .ZN(n1490) );
  OAI21_X2 U2600 ( .B1(n3200), .B2(n3264), .A(n1027), .ZN(n1491) );
  OAI21_X2 U2601 ( .B1(n3198), .B2(n3264), .A(n1026), .ZN(n1492) );
  OAI21_X2 U2602 ( .B1(n3196), .B2(n3264), .A(n1025), .ZN(n1493) );
  OAI21_X2 U2603 ( .B1(n3194), .B2(n3264), .A(n1024), .ZN(n1494) );
  OAI21_X2 U2604 ( .B1(n3192), .B2(n3264), .A(n1022), .ZN(n1495) );
  OAI21_X2 U2605 ( .B1(n3190), .B2(n3263), .A(n1021), .ZN(n1496) );
  OAI21_X2 U2606 ( .B1(n3252), .B2(n3266), .A(n1011), .ZN(n1497) );
  OAI21_X2 U2607 ( .B1(n3250), .B2(n3267), .A(n1000), .ZN(n1498) );
  OAI21_X2 U2608 ( .B1(n3248), .B2(n3267), .A(n989), .ZN(n1499) );
  OAI21_X2 U2609 ( .B1(n3246), .B2(n3266), .A(n986), .ZN(n1500) );
  OAI21_X2 U2610 ( .B1(n3244), .B2(n3266), .A(n985), .ZN(n1501) );
  OAI21_X2 U2611 ( .B1(n3242), .B2(n3266), .A(n984), .ZN(n1502) );
  OAI21_X2 U2612 ( .B1(n3240), .B2(n3266), .A(n983), .ZN(n1503) );
  OAI21_X2 U2613 ( .B1(n3238), .B2(n3266), .A(n982), .ZN(n1504) );
  OAI21_X2 U2614 ( .B1(n3236), .B2(n3266), .A(n981), .ZN(n1505) );
  OAI21_X2 U2615 ( .B1(n3234), .B2(n3266), .A(n980), .ZN(n1506) );
  OAI21_X2 U2616 ( .B1(n3232), .B2(n3266), .A(n1010), .ZN(n1507) );
  OAI21_X2 U2617 ( .B1(n3230), .B2(n3266), .A(n1009), .ZN(n1508) );
  OAI21_X2 U2618 ( .B1(n3228), .B2(n3266), .A(n1008), .ZN(n1509) );
  OAI21_X2 U2619 ( .B1(n3226), .B2(n3267), .A(n1007), .ZN(n1510) );
  OAI21_X2 U2620 ( .B1(n3224), .B2(n3267), .A(n1006), .ZN(n1511) );
  OAI21_X2 U2621 ( .B1(n3222), .B2(n3267), .A(n1005), .ZN(n1512) );
  OAI21_X2 U2622 ( .B1(n3220), .B2(n979), .A(n1004), .ZN(n1513) );
  OAI21_X2 U2623 ( .B1(n3218), .B2(n3268), .A(n1003), .ZN(n1514) );
  OAI21_X2 U2624 ( .B1(n3216), .B2(n979), .A(n1002), .ZN(n1515) );
  OAI21_X2 U2625 ( .B1(n3214), .B2(n979), .A(n1001), .ZN(n1516) );
  OAI21_X2 U2626 ( .B1(n3212), .B2(n3266), .A(n999), .ZN(n1517) );
  OAI21_X2 U2627 ( .B1(n3210), .B2(n3267), .A(n998), .ZN(n1518) );
  OAI21_X2 U2628 ( .B1(n3208), .B2(n979), .A(n997), .ZN(n1519) );
  OAI21_X2 U2629 ( .B1(n3206), .B2(n979), .A(n996), .ZN(n1520) );
  OAI21_X2 U2630 ( .B1(n3204), .B2(n3267), .A(n995), .ZN(n1521) );
  OAI21_X2 U2631 ( .B1(n3202), .B2(n3267), .A(n994), .ZN(n1522) );
  OAI21_X2 U2632 ( .B1(n3200), .B2(n3267), .A(n993), .ZN(n1523) );
  OAI21_X2 U2633 ( .B1(n3198), .B2(n3267), .A(n992), .ZN(n1524) );
  OAI21_X2 U2634 ( .B1(n3196), .B2(n3267), .A(n991), .ZN(n1525) );
  OAI21_X2 U2635 ( .B1(n3194), .B2(n3267), .A(n990), .ZN(n1526) );
  OAI21_X2 U2636 ( .B1(n3192), .B2(n3267), .A(n988), .ZN(n1527) );
  OAI21_X2 U2637 ( .B1(n3190), .B2(n3266), .A(n987), .ZN(n1528) );
  OAI21_X2 U2638 ( .B1(n3252), .B2(n3270), .A(n977), .ZN(n1529) );
  OAI21_X2 U2639 ( .B1(n3250), .B2(n3271), .A(n966), .ZN(n1530) );
  OAI21_X2 U2640 ( .B1(n3248), .B2(n3271), .A(n955), .ZN(n1531) );
  OAI21_X2 U2641 ( .B1(n3246), .B2(n3270), .A(n952), .ZN(n1532) );
  OAI21_X2 U2642 ( .B1(n3244), .B2(n3270), .A(n951), .ZN(n1533) );
  OAI21_X2 U2643 ( .B1(n3242), .B2(n3270), .A(n950), .ZN(n1534) );
  OAI21_X2 U2644 ( .B1(n3240), .B2(n3270), .A(n949), .ZN(n1535) );
  OAI21_X2 U2645 ( .B1(n3238), .B2(n3270), .A(n948), .ZN(n1536) );
  OAI21_X2 U2646 ( .B1(n3236), .B2(n3270), .A(n947), .ZN(n1537) );
  OAI21_X2 U2647 ( .B1(n3234), .B2(n3270), .A(n946), .ZN(n1538) );
  OAI21_X2 U2648 ( .B1(n3232), .B2(n3270), .A(n976), .ZN(n1539) );
  OAI21_X2 U2649 ( .B1(n3230), .B2(n3270), .A(n975), .ZN(n1540) );
  OAI21_X2 U2650 ( .B1(n3228), .B2(n3270), .A(n974), .ZN(n1541) );
  OAI21_X2 U2651 ( .B1(n3226), .B2(n3271), .A(n973), .ZN(n1542) );
  OAI21_X2 U2652 ( .B1(n3224), .B2(n3271), .A(n972), .ZN(n1543) );
  OAI21_X2 U2653 ( .B1(n3222), .B2(n3271), .A(n971), .ZN(n1544) );
  OAI21_X2 U2654 ( .B1(n3220), .B2(n945), .A(n970), .ZN(n1545) );
  OAI21_X2 U2655 ( .B1(n3218), .B2(n3272), .A(n969), .ZN(n1546) );
  OAI21_X2 U2656 ( .B1(n3216), .B2(n945), .A(n968), .ZN(n1547) );
  OAI21_X2 U2657 ( .B1(n3214), .B2(n945), .A(n967), .ZN(n1548) );
  OAI21_X2 U2658 ( .B1(n3212), .B2(n3270), .A(n965), .ZN(n1549) );
  OAI21_X2 U2659 ( .B1(n3210), .B2(n3271), .A(n964), .ZN(n1550) );
  OAI21_X2 U2660 ( .B1(n3208), .B2(n945), .A(n963), .ZN(n1551) );
  OAI21_X2 U2661 ( .B1(n3206), .B2(n945), .A(n962), .ZN(n1552) );
  OAI21_X2 U2662 ( .B1(n3204), .B2(n3271), .A(n961), .ZN(n1553) );
  OAI21_X2 U2663 ( .B1(n3202), .B2(n3271), .A(n960), .ZN(n1554) );
  OAI21_X2 U2664 ( .B1(n3200), .B2(n3271), .A(n959), .ZN(n1555) );
  OAI21_X2 U2665 ( .B1(n3198), .B2(n3271), .A(n958), .ZN(n1556) );
  OAI21_X2 U2666 ( .B1(n3196), .B2(n3271), .A(n957), .ZN(n1557) );
  OAI21_X2 U2667 ( .B1(n3194), .B2(n3271), .A(n956), .ZN(n1558) );
  OAI21_X2 U2668 ( .B1(n3192), .B2(n3271), .A(n954), .ZN(n1559) );
  OAI21_X2 U2669 ( .B1(n3190), .B2(n3270), .A(n953), .ZN(n1560) );
  OAI21_X2 U2670 ( .B1(n3252), .B2(n3275), .A(n944), .ZN(n1561) );
  OAI21_X2 U2671 ( .B1(n3250), .B2(n3275), .A(n933), .ZN(n1562) );
  OAI21_X2 U2672 ( .B1(n3248), .B2(n3276), .A(n922), .ZN(n1563) );
  OAI21_X2 U2673 ( .B1(n3246), .B2(n3275), .A(n919), .ZN(n1564) );
  OAI21_X2 U2674 ( .B1(n3244), .B2(n3275), .A(n918), .ZN(n1565) );
  OAI21_X2 U2675 ( .B1(n3242), .B2(n3275), .A(n917), .ZN(n1566) );
  OAI21_X2 U2676 ( .B1(n3240), .B2(n3275), .A(n916), .ZN(n1567) );
  OAI21_X2 U2677 ( .B1(n3238), .B2(n3275), .A(n915), .ZN(n1568) );
  OAI21_X2 U2678 ( .B1(n3236), .B2(n3275), .A(n914), .ZN(n1569) );
  OAI21_X2 U2679 ( .B1(n3234), .B2(n3275), .A(n913), .ZN(n1570) );
  OAI21_X2 U2680 ( .B1(n3232), .B2(n3275), .A(n943), .ZN(n1571) );
  OAI21_X2 U2681 ( .B1(n3230), .B2(n3275), .A(n942), .ZN(n1572) );
  OAI21_X2 U2682 ( .B1(n3228), .B2(n3275), .A(n941), .ZN(n1573) );
  OAI21_X2 U2683 ( .B1(n3226), .B2(n3276), .A(n940), .ZN(n1574) );
  OAI21_X2 U2684 ( .B1(n3224), .B2(n3276), .A(n939), .ZN(n1575) );
  OAI21_X2 U2685 ( .B1(n3222), .B2(n3276), .A(n938), .ZN(n1576) );
  OAI21_X2 U2686 ( .B1(n3220), .B2(n912), .A(n937), .ZN(n1577) );
  OAI21_X2 U2687 ( .B1(n3218), .B2(n3276), .A(n936), .ZN(n1578) );
  OAI21_X2 U2688 ( .B1(n3216), .B2(n912), .A(n935), .ZN(n1579) );
  OAI21_X2 U2689 ( .B1(n3214), .B2(n912), .A(n934), .ZN(n1580) );
  OAI21_X2 U2690 ( .B1(n3212), .B2(n3277), .A(n932), .ZN(n1581) );
  OAI21_X2 U2691 ( .B1(n3210), .B2(n3276), .A(n931), .ZN(n1582) );
  OAI21_X2 U2692 ( .B1(n3208), .B2(n912), .A(n930), .ZN(n1583) );
  OAI21_X2 U2693 ( .B1(n3206), .B2(n912), .A(n929), .ZN(n1584) );
  OAI21_X2 U2694 ( .B1(n3204), .B2(n3276), .A(n928), .ZN(n1585) );
  OAI21_X2 U2695 ( .B1(n3202), .B2(n3276), .A(n927), .ZN(n1586) );
  OAI21_X2 U2696 ( .B1(n3200), .B2(n3276), .A(n926), .ZN(n1587) );
  OAI21_X2 U2697 ( .B1(n3198), .B2(n3276), .A(n925), .ZN(n1588) );
  OAI21_X2 U2698 ( .B1(n3196), .B2(n3276), .A(n924), .ZN(n1589) );
  OAI21_X2 U2699 ( .B1(n3194), .B2(n3276), .A(n923), .ZN(n1590) );
  OAI21_X2 U2700 ( .B1(n3192), .B2(n3276), .A(n921), .ZN(n1591) );
  OAI21_X2 U2701 ( .B1(n3190), .B2(n3275), .A(n920), .ZN(n1592) );
  OAI21_X2 U2702 ( .B1(n3252), .B2(n3279), .A(n910), .ZN(n1593) );
  OAI21_X2 U2703 ( .B1(n3250), .B2(n3279), .A(n899), .ZN(n1594) );
  OAI21_X2 U2704 ( .B1(n3248), .B2(n3280), .A(n888), .ZN(n1595) );
  OAI21_X2 U2705 ( .B1(n3246), .B2(n3279), .A(n885), .ZN(n1596) );
  OAI21_X2 U2706 ( .B1(n3244), .B2(n3279), .A(n884), .ZN(n1597) );
  OAI21_X2 U2707 ( .B1(n3242), .B2(n3279), .A(n883), .ZN(n1598) );
  OAI21_X2 U2708 ( .B1(n3240), .B2(n3279), .A(n882), .ZN(n1599) );
  OAI21_X2 U2709 ( .B1(n3238), .B2(n3279), .A(n881), .ZN(n1600) );
  OAI21_X2 U2710 ( .B1(n3236), .B2(n3279), .A(n880), .ZN(n1601) );
  OAI21_X2 U2711 ( .B1(n3234), .B2(n3279), .A(n879), .ZN(n1602) );
  OAI21_X2 U2712 ( .B1(n3232), .B2(n3279), .A(n909), .ZN(n1603) );
  OAI21_X2 U2713 ( .B1(n3230), .B2(n3279), .A(n908), .ZN(n1604) );
  OAI21_X2 U2714 ( .B1(n3228), .B2(n3279), .A(n907), .ZN(n1605) );
  OAI21_X2 U2715 ( .B1(n3226), .B2(n3280), .A(n906), .ZN(n1606) );
  OAI21_X2 U2716 ( .B1(n3224), .B2(n3280), .A(n905), .ZN(n1607) );
  OAI21_X2 U2717 ( .B1(n3222), .B2(n3280), .A(n904), .ZN(n1608) );
  OAI21_X2 U2718 ( .B1(n3220), .B2(n878), .A(n903), .ZN(n1609) );
  OAI21_X2 U2719 ( .B1(n3218), .B2(n3280), .A(n902), .ZN(n1610) );
  OAI21_X2 U2720 ( .B1(n3216), .B2(n878), .A(n901), .ZN(n1611) );
  OAI21_X2 U2721 ( .B1(n3214), .B2(n878), .A(n900), .ZN(n1612) );
  OAI21_X2 U2722 ( .B1(n3212), .B2(n3281), .A(n898), .ZN(n1613) );
  OAI21_X2 U2723 ( .B1(n3210), .B2(n3280), .A(n897), .ZN(n1614) );
  OAI21_X2 U2724 ( .B1(n3208), .B2(n878), .A(n896), .ZN(n1615) );
  OAI21_X2 U2725 ( .B1(n3206), .B2(n878), .A(n895), .ZN(n1616) );
  OAI21_X2 U2726 ( .B1(n3204), .B2(n3280), .A(n894), .ZN(n1617) );
  OAI21_X2 U2727 ( .B1(n3202), .B2(n3280), .A(n893), .ZN(n1618) );
  OAI21_X2 U2728 ( .B1(n3200), .B2(n3280), .A(n892), .ZN(n1619) );
  OAI21_X2 U2729 ( .B1(n3198), .B2(n3280), .A(n891), .ZN(n1620) );
  OAI21_X2 U2730 ( .B1(n3196), .B2(n3280), .A(n890), .ZN(n1621) );
  OAI21_X2 U2731 ( .B1(n3194), .B2(n3280), .A(n889), .ZN(n1622) );
  OAI21_X2 U2732 ( .B1(n3192), .B2(n3280), .A(n887), .ZN(n1623) );
  OAI21_X2 U2733 ( .B1(n3190), .B2(n3279), .A(n886), .ZN(n1624) );
  OAI21_X2 U2734 ( .B1(n3252), .B2(n3282), .A(n874), .ZN(n1625) );
  OAI21_X2 U2735 ( .B1(n3250), .B2(n3283), .A(n863), .ZN(n1626) );
  OAI21_X2 U2736 ( .B1(n3248), .B2(n3283), .A(n852), .ZN(n1627) );
  OAI21_X2 U2737 ( .B1(n3246), .B2(n3282), .A(n849), .ZN(n1628) );
  OAI21_X2 U2738 ( .B1(n3244), .B2(n3282), .A(n848), .ZN(n1629) );
  OAI21_X2 U2739 ( .B1(n3242), .B2(n3282), .A(n847), .ZN(n1630) );
  OAI21_X2 U2740 ( .B1(n3240), .B2(n3282), .A(n846), .ZN(n1631) );
  OAI21_X2 U2741 ( .B1(n3238), .B2(n3282), .A(n845), .ZN(n1632) );
  OAI21_X2 U2742 ( .B1(n3236), .B2(n3282), .A(n844), .ZN(n1633) );
  OAI21_X2 U2743 ( .B1(n3234), .B2(n3282), .A(n843), .ZN(n1634) );
  OAI21_X2 U2744 ( .B1(n3232), .B2(n3282), .A(n873), .ZN(n1635) );
  OAI21_X2 U2745 ( .B1(n3230), .B2(n3282), .A(n872), .ZN(n1636) );
  OAI21_X2 U2746 ( .B1(n3228), .B2(n3282), .A(n871), .ZN(n1637) );
  OAI21_X2 U2747 ( .B1(n3226), .B2(n3283), .A(n870), .ZN(n1638) );
  OAI21_X2 U2748 ( .B1(n3224), .B2(n3283), .A(n869), .ZN(n1639) );
  OAI21_X2 U2749 ( .B1(n3222), .B2(n3283), .A(n868), .ZN(n1640) );
  OAI21_X2 U2750 ( .B1(n3220), .B2(n842), .A(n867), .ZN(n1641) );
  OAI21_X2 U2751 ( .B1(n3218), .B2(n3284), .A(n866), .ZN(n1642) );
  OAI21_X2 U2752 ( .B1(n3216), .B2(n842), .A(n865), .ZN(n1643) );
  OAI21_X2 U2753 ( .B1(n3214), .B2(n842), .A(n864), .ZN(n1644) );
  OAI21_X2 U2754 ( .B1(n3212), .B2(n3282), .A(n862), .ZN(n1645) );
  OAI21_X2 U2755 ( .B1(n3210), .B2(n3283), .A(n861), .ZN(n1646) );
  OAI21_X2 U2756 ( .B1(n3208), .B2(n842), .A(n860), .ZN(n1647) );
  OAI21_X2 U2757 ( .B1(n3206), .B2(n842), .A(n859), .ZN(n1648) );
  OAI21_X2 U2758 ( .B1(n3204), .B2(n3283), .A(n858), .ZN(n1649) );
  OAI21_X2 U2759 ( .B1(n3202), .B2(n3283), .A(n857), .ZN(n1650) );
  OAI21_X2 U2760 ( .B1(n3200), .B2(n3283), .A(n856), .ZN(n1651) );
  OAI21_X2 U2761 ( .B1(n3198), .B2(n3283), .A(n855), .ZN(n1652) );
  OAI21_X2 U2762 ( .B1(n3196), .B2(n3283), .A(n854), .ZN(n1653) );
  OAI21_X2 U2763 ( .B1(n3194), .B2(n3283), .A(n853), .ZN(n1654) );
  OAI21_X2 U2764 ( .B1(n3192), .B2(n3283), .A(n851), .ZN(n1655) );
  OAI21_X2 U2765 ( .B1(n3190), .B2(n3282), .A(n850), .ZN(n1656) );
  OAI21_X2 U2766 ( .B1(n3252), .B2(n3286), .A(n841), .ZN(n1657) );
  OAI21_X2 U2767 ( .B1(n3250), .B2(n3287), .A(n830), .ZN(n1658) );
  OAI21_X2 U2768 ( .B1(n3248), .B2(n3287), .A(n819), .ZN(n1659) );
  OAI21_X2 U2769 ( .B1(n3246), .B2(n3286), .A(n816), .ZN(n1660) );
  OAI21_X2 U2770 ( .B1(n3244), .B2(n3286), .A(n815), .ZN(n1661) );
  OAI21_X2 U2771 ( .B1(n3242), .B2(n3286), .A(n814), .ZN(n1662) );
  OAI21_X2 U2772 ( .B1(n3240), .B2(n3286), .A(n813), .ZN(n1663) );
  OAI21_X2 U2773 ( .B1(n3238), .B2(n3286), .A(n812), .ZN(n1664) );
  OAI21_X2 U2774 ( .B1(n3236), .B2(n3286), .A(n811), .ZN(n1665) );
  OAI21_X2 U2775 ( .B1(n3234), .B2(n3286), .A(n810), .ZN(n1666) );
  OAI21_X2 U2776 ( .B1(n3232), .B2(n3286), .A(n840), .ZN(n1667) );
  OAI21_X2 U2777 ( .B1(n3230), .B2(n3286), .A(n839), .ZN(n1668) );
  OAI21_X2 U2778 ( .B1(n3228), .B2(n3286), .A(n838), .ZN(n1669) );
  OAI21_X2 U2779 ( .B1(n3226), .B2(n3287), .A(n837), .ZN(n1670) );
  OAI21_X2 U2780 ( .B1(n3224), .B2(n3287), .A(n836), .ZN(n1671) );
  OAI21_X2 U2781 ( .B1(n3222), .B2(n3287), .A(n835), .ZN(n1672) );
  OAI21_X2 U2782 ( .B1(n3220), .B2(n809), .A(n834), .ZN(n1673) );
  OAI21_X2 U2783 ( .B1(n3218), .B2(n3288), .A(n833), .ZN(n1674) );
  OAI21_X2 U2784 ( .B1(n3216), .B2(n809), .A(n832), .ZN(n1675) );
  OAI21_X2 U2785 ( .B1(n3214), .B2(n809), .A(n831), .ZN(n1676) );
  OAI21_X2 U2786 ( .B1(n3212), .B2(n3286), .A(n829), .ZN(n1677) );
  OAI21_X2 U2787 ( .B1(n3210), .B2(n3287), .A(n828), .ZN(n1678) );
  OAI21_X2 U2788 ( .B1(n3208), .B2(n809), .A(n827), .ZN(n1679) );
  OAI21_X2 U2789 ( .B1(n3206), .B2(n809), .A(n826), .ZN(n1680) );
  OAI21_X2 U2790 ( .B1(n3204), .B2(n3287), .A(n825), .ZN(n1681) );
  OAI21_X2 U2791 ( .B1(n3202), .B2(n3287), .A(n824), .ZN(n1682) );
  OAI21_X2 U2792 ( .B1(n3200), .B2(n3287), .A(n823), .ZN(n1683) );
  OAI21_X2 U2793 ( .B1(n3198), .B2(n3287), .A(n822), .ZN(n1684) );
  OAI21_X2 U2794 ( .B1(n3196), .B2(n3287), .A(n821), .ZN(n1685) );
  OAI21_X2 U2795 ( .B1(n3194), .B2(n3287), .A(n820), .ZN(n1686) );
  OAI21_X2 U2796 ( .B1(n3192), .B2(n3287), .A(n818), .ZN(n1687) );
  OAI21_X2 U2797 ( .B1(n3190), .B2(n3286), .A(n817), .ZN(n1688) );
  OAI21_X2 U2798 ( .B1(n3252), .B2(n3291), .A(n808), .ZN(n1689) );
  OAI21_X2 U2799 ( .B1(n3250), .B2(n3291), .A(n797), .ZN(n1690) );
  OAI21_X2 U2800 ( .B1(n3248), .B2(n3292), .A(n786), .ZN(n1691) );
  OAI21_X2 U2801 ( .B1(n3246), .B2(n3291), .A(n783), .ZN(n1692) );
  OAI21_X2 U2802 ( .B1(n3244), .B2(n3291), .A(n782), .ZN(n1693) );
  OAI21_X2 U2803 ( .B1(n3242), .B2(n3291), .A(n781), .ZN(n1694) );
  OAI21_X2 U2804 ( .B1(n3240), .B2(n3291), .A(n780), .ZN(n1695) );
  OAI21_X2 U2805 ( .B1(n3238), .B2(n3291), .A(n779), .ZN(n1696) );
  OAI21_X2 U2806 ( .B1(n3236), .B2(n3291), .A(n778), .ZN(n1697) );
  OAI21_X2 U2807 ( .B1(n3234), .B2(n3291), .A(n777), .ZN(n1698) );
  OAI21_X2 U2808 ( .B1(n3232), .B2(n3291), .A(n807), .ZN(n1699) );
  OAI21_X2 U2809 ( .B1(n3230), .B2(n3291), .A(n806), .ZN(n1700) );
  OAI21_X2 U2810 ( .B1(n3228), .B2(n3291), .A(n805), .ZN(n1701) );
  OAI21_X2 U2811 ( .B1(n3226), .B2(n3292), .A(n804), .ZN(n1702) );
  OAI21_X2 U2812 ( .B1(n3224), .B2(n3292), .A(n803), .ZN(n1703) );
  OAI21_X2 U2813 ( .B1(n3222), .B2(n3292), .A(n802), .ZN(n1704) );
  OAI21_X2 U2814 ( .B1(n3220), .B2(n776), .A(n801), .ZN(n1705) );
  OAI21_X2 U2815 ( .B1(n3218), .B2(n3292), .A(n800), .ZN(n1706) );
  OAI21_X2 U2816 ( .B1(n3216), .B2(n776), .A(n799), .ZN(n1707) );
  OAI21_X2 U2817 ( .B1(n3214), .B2(n776), .A(n798), .ZN(n1708) );
  OAI21_X2 U2818 ( .B1(n3212), .B2(n3293), .A(n796), .ZN(n1709) );
  OAI21_X2 U2819 ( .B1(n3210), .B2(n3292), .A(n795), .ZN(n1710) );
  OAI21_X2 U2820 ( .B1(n3208), .B2(n776), .A(n794), .ZN(n1711) );
  OAI21_X2 U2821 ( .B1(n3206), .B2(n776), .A(n793), .ZN(n1712) );
  OAI21_X2 U2822 ( .B1(n3204), .B2(n3292), .A(n792), .ZN(n1713) );
  OAI21_X2 U2823 ( .B1(n3202), .B2(n3292), .A(n791), .ZN(n1714) );
  OAI21_X2 U2824 ( .B1(n3200), .B2(n3292), .A(n790), .ZN(n1715) );
  OAI21_X2 U2825 ( .B1(n3198), .B2(n3292), .A(n789), .ZN(n1716) );
  OAI21_X2 U2826 ( .B1(n3196), .B2(n3292), .A(n788), .ZN(n1717) );
  OAI21_X2 U2827 ( .B1(n3194), .B2(n3292), .A(n787), .ZN(n1718) );
  OAI21_X2 U2828 ( .B1(n3192), .B2(n3292), .A(n785), .ZN(n1719) );
  OAI21_X2 U2829 ( .B1(n3190), .B2(n3291), .A(n784), .ZN(n1720) );
  OAI21_X2 U2830 ( .B1(n3252), .B2(n3295), .A(n774), .ZN(n1721) );
  OAI21_X2 U2831 ( .B1(n3250), .B2(n3295), .A(n763), .ZN(n1722) );
  OAI21_X2 U2832 ( .B1(n3248), .B2(n3296), .A(n752), .ZN(n1723) );
  OAI21_X2 U2833 ( .B1(n3246), .B2(n3295), .A(n749), .ZN(n1724) );
  OAI21_X2 U2834 ( .B1(n3244), .B2(n3295), .A(n748), .ZN(n1725) );
  OAI21_X2 U2835 ( .B1(n3242), .B2(n3295), .A(n747), .ZN(n1726) );
  OAI21_X2 U2836 ( .B1(n3240), .B2(n3295), .A(n746), .ZN(n1727) );
  OAI21_X2 U2837 ( .B1(n3238), .B2(n3295), .A(n745), .ZN(n1728) );
  OAI21_X2 U2838 ( .B1(n3236), .B2(n3295), .A(n744), .ZN(n1729) );
  OAI21_X2 U2839 ( .B1(n3234), .B2(n3295), .A(n743), .ZN(n1730) );
  OAI21_X2 U2840 ( .B1(n3232), .B2(n3295), .A(n773), .ZN(n1731) );
  OAI21_X2 U2841 ( .B1(n3230), .B2(n3295), .A(n772), .ZN(n1732) );
  OAI21_X2 U2842 ( .B1(n3228), .B2(n3295), .A(n771), .ZN(n1733) );
  OAI21_X2 U2843 ( .B1(n3226), .B2(n3296), .A(n770), .ZN(n1734) );
  OAI21_X2 U2844 ( .B1(n3224), .B2(n3296), .A(n769), .ZN(n1735) );
  OAI21_X2 U2845 ( .B1(n3222), .B2(n3296), .A(n768), .ZN(n1736) );
  OAI21_X2 U2846 ( .B1(n3220), .B2(n742), .A(n767), .ZN(n1737) );
  OAI21_X2 U2847 ( .B1(n3218), .B2(n3296), .A(n766), .ZN(n1738) );
  OAI21_X2 U2848 ( .B1(n3216), .B2(n742), .A(n765), .ZN(n1739) );
  OAI21_X2 U2849 ( .B1(n3214), .B2(n742), .A(n764), .ZN(n1740) );
  OAI21_X2 U2850 ( .B1(n3212), .B2(n3297), .A(n762), .ZN(n1741) );
  OAI21_X2 U2851 ( .B1(n3210), .B2(n3296), .A(n761), .ZN(n1742) );
  OAI21_X2 U2852 ( .B1(n3208), .B2(n742), .A(n760), .ZN(n1743) );
  OAI21_X2 U2853 ( .B1(n3206), .B2(n742), .A(n759), .ZN(n1744) );
  OAI21_X2 U2854 ( .B1(n3204), .B2(n3296), .A(n758), .ZN(n1745) );
  OAI21_X2 U2855 ( .B1(n3202), .B2(n3296), .A(n757), .ZN(n1746) );
  OAI21_X2 U2856 ( .B1(n3200), .B2(n3296), .A(n756), .ZN(n1747) );
  OAI21_X2 U2857 ( .B1(n3198), .B2(n3296), .A(n755), .ZN(n1748) );
  OAI21_X2 U2858 ( .B1(n3196), .B2(n3296), .A(n754), .ZN(n1749) );
  OAI21_X2 U2859 ( .B1(n3194), .B2(n3296), .A(n753), .ZN(n1750) );
  OAI21_X2 U2860 ( .B1(n3192), .B2(n3296), .A(n751), .ZN(n1751) );
  OAI21_X2 U2861 ( .B1(n3190), .B2(n3295), .A(n750), .ZN(n1752) );
  OAI21_X2 U2862 ( .B1(n3253), .B2(n3302), .A(n707), .ZN(n1753) );
  OAI21_X2 U2863 ( .B1(n3251), .B2(n3303), .A(n696), .ZN(n1754) );
  OAI21_X2 U2864 ( .B1(n3249), .B2(n3303), .A(n685), .ZN(n1755) );
  OAI21_X2 U2865 ( .B1(n3247), .B2(n3302), .A(n682), .ZN(n1756) );
  OAI21_X2 U2866 ( .B1(n3245), .B2(n3302), .A(n681), .ZN(n1757) );
  OAI21_X2 U2867 ( .B1(n3243), .B2(n3302), .A(n680), .ZN(n1758) );
  OAI21_X2 U2868 ( .B1(n3241), .B2(n3302), .A(n679), .ZN(n1759) );
  OAI21_X2 U2869 ( .B1(n3239), .B2(n3302), .A(n678), .ZN(n1760) );
  OAI21_X2 U2870 ( .B1(n3237), .B2(n3302), .A(n677), .ZN(n1761) );
  OAI21_X2 U2871 ( .B1(n3235), .B2(n3302), .A(n676), .ZN(n1762) );
  OAI21_X2 U2872 ( .B1(n3233), .B2(n3302), .A(n706), .ZN(n1763) );
  OAI21_X2 U2873 ( .B1(n3231), .B2(n3302), .A(n705), .ZN(n1764) );
  OAI21_X2 U2874 ( .B1(n3229), .B2(n3302), .A(n704), .ZN(n1765) );
  OAI21_X2 U2875 ( .B1(n3227), .B2(n3303), .A(n703), .ZN(n1766) );
  OAI21_X2 U2876 ( .B1(n3225), .B2(n3303), .A(n702), .ZN(n1767) );
  OAI21_X2 U2877 ( .B1(n3223), .B2(n3303), .A(n701), .ZN(n1768) );
  OAI21_X2 U2878 ( .B1(n3221), .B2(n675), .A(n700), .ZN(n1769) );
  OAI21_X2 U2879 ( .B1(n3219), .B2(n3304), .A(n699), .ZN(n1770) );
  OAI21_X2 U2880 ( .B1(n3217), .B2(n675), .A(n698), .ZN(n1771) );
  OAI21_X2 U2881 ( .B1(n3215), .B2(n675), .A(n697), .ZN(n1772) );
  OAI21_X2 U2882 ( .B1(n3213), .B2(n3302), .A(n695), .ZN(n1773) );
  OAI21_X2 U2883 ( .B1(n3211), .B2(n3303), .A(n694), .ZN(n1774) );
  OAI21_X2 U2884 ( .B1(n3209), .B2(n675), .A(n693), .ZN(n1775) );
  OAI21_X2 U2885 ( .B1(n3207), .B2(n675), .A(n692), .ZN(n1776) );
  OAI21_X2 U2886 ( .B1(n3205), .B2(n3303), .A(n691), .ZN(n1777) );
  OAI21_X2 U2887 ( .B1(n3203), .B2(n3303), .A(n690), .ZN(n1778) );
  OAI21_X2 U2888 ( .B1(n3201), .B2(n3303), .A(n689), .ZN(n1779) );
  OAI21_X2 U2889 ( .B1(n3199), .B2(n3303), .A(n688), .ZN(n1780) );
  OAI21_X2 U2890 ( .B1(n3197), .B2(n3303), .A(n687), .ZN(n1781) );
  OAI21_X2 U2891 ( .B1(n3195), .B2(n3303), .A(n686), .ZN(n1782) );
  OAI21_X2 U2892 ( .B1(n3193), .B2(n3303), .A(n684), .ZN(n1783) );
  OAI21_X2 U2893 ( .B1(n3191), .B2(n3302), .A(n683), .ZN(n1784) );
  OAI21_X2 U2894 ( .B1(n3253), .B2(n3306), .A(n674), .ZN(n1785) );
  OAI21_X2 U2895 ( .B1(n3251), .B2(n3307), .A(n663), .ZN(n1786) );
  OAI21_X2 U2896 ( .B1(n3249), .B2(n3307), .A(n652), .ZN(n1787) );
  OAI21_X2 U2897 ( .B1(n3247), .B2(n3306), .A(n649), .ZN(n1788) );
  OAI21_X2 U2898 ( .B1(n3245), .B2(n3306), .A(n648), .ZN(n1789) );
  OAI21_X2 U2899 ( .B1(n3243), .B2(n3306), .A(n647), .ZN(n1790) );
  OAI21_X2 U2900 ( .B1(n3241), .B2(n3306), .A(n646), .ZN(n1791) );
  OAI21_X2 U2901 ( .B1(n3239), .B2(n3306), .A(n645), .ZN(n1792) );
  OAI21_X2 U2902 ( .B1(n3237), .B2(n3306), .A(n644), .ZN(n1793) );
  OAI21_X2 U2903 ( .B1(n3235), .B2(n3306), .A(n643), .ZN(n1794) );
  OAI21_X2 U2904 ( .B1(n3233), .B2(n3306), .A(n673), .ZN(n1795) );
  OAI21_X2 U2905 ( .B1(n3231), .B2(n3306), .A(n672), .ZN(n1796) );
  OAI21_X2 U2906 ( .B1(n3229), .B2(n3306), .A(n671), .ZN(n1797) );
  OAI21_X2 U2907 ( .B1(n3227), .B2(n3307), .A(n670), .ZN(n1798) );
  OAI21_X2 U2908 ( .B1(n3225), .B2(n3307), .A(n669), .ZN(n1799) );
  OAI21_X2 U2909 ( .B1(n3223), .B2(n3307), .A(n668), .ZN(n1800) );
  OAI21_X2 U2910 ( .B1(n3221), .B2(n642), .A(n667), .ZN(n1801) );
  OAI21_X2 U2911 ( .B1(n3219), .B2(n3308), .A(n666), .ZN(n1802) );
  OAI21_X2 U2912 ( .B1(n3217), .B2(n642), .A(n665), .ZN(n1803) );
  OAI21_X2 U2913 ( .B1(n3215), .B2(n642), .A(n664), .ZN(n1804) );
  OAI21_X2 U2914 ( .B1(n3213), .B2(n3306), .A(n662), .ZN(n1805) );
  OAI21_X2 U2915 ( .B1(n3211), .B2(n3307), .A(n661), .ZN(n1806) );
  OAI21_X2 U2916 ( .B1(n3209), .B2(n642), .A(n660), .ZN(n1807) );
  OAI21_X2 U2917 ( .B1(n3207), .B2(n642), .A(n659), .ZN(n1808) );
  OAI21_X2 U2918 ( .B1(n3205), .B2(n3307), .A(n658), .ZN(n1809) );
  OAI21_X2 U2919 ( .B1(n3203), .B2(n3307), .A(n657), .ZN(n1810) );
  OAI21_X2 U2920 ( .B1(n3201), .B2(n3307), .A(n656), .ZN(n1811) );
  OAI21_X2 U2921 ( .B1(n3199), .B2(n3307), .A(n655), .ZN(n1812) );
  OAI21_X2 U2922 ( .B1(n3197), .B2(n3307), .A(n654), .ZN(n1813) );
  OAI21_X2 U2923 ( .B1(n3195), .B2(n3307), .A(n653), .ZN(n1814) );
  OAI21_X2 U2924 ( .B1(n3193), .B2(n3307), .A(n651), .ZN(n1815) );
  OAI21_X2 U2925 ( .B1(n3191), .B2(n3306), .A(n650), .ZN(n1816) );
  OAI21_X2 U2926 ( .B1(n3253), .B2(n3311), .A(n641), .ZN(n1817) );
  OAI21_X2 U2927 ( .B1(n3251), .B2(n3311), .A(n630), .ZN(n1818) );
  OAI21_X2 U2928 ( .B1(n3249), .B2(n3312), .A(n619), .ZN(n1819) );
  OAI21_X2 U2929 ( .B1(n3247), .B2(n3311), .A(n616), .ZN(n1820) );
  OAI21_X2 U2930 ( .B1(n3245), .B2(n3311), .A(n615), .ZN(n1821) );
  OAI21_X2 U2931 ( .B1(n3243), .B2(n3311), .A(n614), .ZN(n1822) );
  OAI21_X2 U2932 ( .B1(n3241), .B2(n3311), .A(n613), .ZN(n1823) );
  OAI21_X2 U2933 ( .B1(n3239), .B2(n3311), .A(n612), .ZN(n1824) );
  OAI21_X2 U2934 ( .B1(n3237), .B2(n3311), .A(n611), .ZN(n1825) );
  OAI21_X2 U2935 ( .B1(n3235), .B2(n3311), .A(n610), .ZN(n1826) );
  OAI21_X2 U2936 ( .B1(n3233), .B2(n3311), .A(n640), .ZN(n1827) );
  OAI21_X2 U2937 ( .B1(n3231), .B2(n3311), .A(n639), .ZN(n1828) );
  OAI21_X2 U2938 ( .B1(n3229), .B2(n3311), .A(n638), .ZN(n1829) );
  OAI21_X2 U2939 ( .B1(n3227), .B2(n3312), .A(n637), .ZN(n1830) );
  OAI21_X2 U2940 ( .B1(n3225), .B2(n3312), .A(n636), .ZN(n1831) );
  OAI21_X2 U2941 ( .B1(n3223), .B2(n3312), .A(n635), .ZN(n1832) );
  OAI21_X2 U2942 ( .B1(n3221), .B2(n609), .A(n634), .ZN(n1833) );
  OAI21_X2 U2943 ( .B1(n3219), .B2(n3312), .A(n633), .ZN(n1834) );
  OAI21_X2 U2944 ( .B1(n3217), .B2(n609), .A(n632), .ZN(n1835) );
  OAI21_X2 U2945 ( .B1(n3215), .B2(n609), .A(n631), .ZN(n1836) );
  OAI21_X2 U2946 ( .B1(n3213), .B2(n3313), .A(n629), .ZN(n1837) );
  OAI21_X2 U2947 ( .B1(n3211), .B2(n3312), .A(n628), .ZN(n1838) );
  OAI21_X2 U2948 ( .B1(n3209), .B2(n609), .A(n627), .ZN(n1839) );
  OAI21_X2 U2949 ( .B1(n3207), .B2(n609), .A(n626), .ZN(n1840) );
  OAI21_X2 U2950 ( .B1(n3205), .B2(n3312), .A(n625), .ZN(n1841) );
  OAI21_X2 U2951 ( .B1(n3203), .B2(n3312), .A(n624), .ZN(n1842) );
  OAI21_X2 U2952 ( .B1(n3201), .B2(n3312), .A(n623), .ZN(n1843) );
  OAI21_X2 U2953 ( .B1(n3199), .B2(n3312), .A(n622), .ZN(n1844) );
  OAI21_X2 U2954 ( .B1(n3197), .B2(n3312), .A(n621), .ZN(n1845) );
  OAI21_X2 U2955 ( .B1(n3195), .B2(n3312), .A(n620), .ZN(n1846) );
  OAI21_X2 U2956 ( .B1(n3193), .B2(n3312), .A(n618), .ZN(n1847) );
  OAI21_X2 U2957 ( .B1(n3191), .B2(n3311), .A(n617), .ZN(n1848) );
  OAI21_X2 U2958 ( .B1(n3253), .B2(n3315), .A(n607), .ZN(n1849) );
  OAI21_X2 U2959 ( .B1(n3251), .B2(n3315), .A(n596), .ZN(n1850) );
  OAI21_X2 U2960 ( .B1(n3249), .B2(n3316), .A(n585), .ZN(n1851) );
  OAI21_X2 U2961 ( .B1(n3247), .B2(n3315), .A(n582), .ZN(n1852) );
  OAI21_X2 U2962 ( .B1(n3245), .B2(n3315), .A(n581), .ZN(n1853) );
  OAI21_X2 U2963 ( .B1(n3243), .B2(n3315), .A(n580), .ZN(n1854) );
  OAI21_X2 U2964 ( .B1(n3241), .B2(n3315), .A(n579), .ZN(n1855) );
  OAI21_X2 U2965 ( .B1(n3239), .B2(n3315), .A(n578), .ZN(n1856) );
  OAI21_X2 U2966 ( .B1(n3237), .B2(n3315), .A(n577), .ZN(n1857) );
  OAI21_X2 U2967 ( .B1(n3235), .B2(n3315), .A(n576), .ZN(n1858) );
  OAI21_X2 U2968 ( .B1(n3233), .B2(n3315), .A(n606), .ZN(n1859) );
  OAI21_X2 U2969 ( .B1(n3231), .B2(n3315), .A(n605), .ZN(n1860) );
  OAI21_X2 U2970 ( .B1(n3229), .B2(n3315), .A(n604), .ZN(n1861) );
  OAI21_X2 U2971 ( .B1(n3227), .B2(n3316), .A(n603), .ZN(n1862) );
  OAI21_X2 U2972 ( .B1(n3225), .B2(n3316), .A(n602), .ZN(n1863) );
  OAI21_X2 U2973 ( .B1(n3223), .B2(n3316), .A(n601), .ZN(n1864) );
  OAI21_X2 U2974 ( .B1(n3221), .B2(n575), .A(n600), .ZN(n1865) );
  OAI21_X2 U2975 ( .B1(n3219), .B2(n3316), .A(n599), .ZN(n1866) );
  OAI21_X2 U2976 ( .B1(n3217), .B2(n575), .A(n598), .ZN(n1867) );
  OAI21_X2 U2977 ( .B1(n3215), .B2(n575), .A(n597), .ZN(n1868) );
  OAI21_X2 U2978 ( .B1(n3213), .B2(n3317), .A(n595), .ZN(n1869) );
  OAI21_X2 U2979 ( .B1(n3211), .B2(n3316), .A(n594), .ZN(n1870) );
  OAI21_X2 U2980 ( .B1(n3209), .B2(n575), .A(n593), .ZN(n1871) );
  OAI21_X2 U2981 ( .B1(n3207), .B2(n575), .A(n592), .ZN(n1872) );
  OAI21_X2 U2982 ( .B1(n3205), .B2(n3316), .A(n591), .ZN(n1873) );
  OAI21_X2 U2983 ( .B1(n3203), .B2(n3316), .A(n590), .ZN(n1874) );
  OAI21_X2 U2984 ( .B1(n3201), .B2(n3316), .A(n589), .ZN(n1875) );
  OAI21_X2 U2985 ( .B1(n3199), .B2(n3316), .A(n588), .ZN(n1876) );
  OAI21_X2 U2986 ( .B1(n3197), .B2(n3316), .A(n587), .ZN(n1877) );
  OAI21_X2 U2987 ( .B1(n3195), .B2(n3316), .A(n586), .ZN(n1878) );
  OAI21_X2 U2988 ( .B1(n3193), .B2(n3316), .A(n584), .ZN(n1879) );
  OAI21_X2 U2989 ( .B1(n3191), .B2(n3315), .A(n583), .ZN(n1880) );
  OAI21_X2 U2990 ( .B1(n3253), .B2(n3318), .A(n573), .ZN(n1881) );
  OAI21_X2 U2991 ( .B1(n3251), .B2(n3319), .A(n562), .ZN(n1882) );
  OAI21_X2 U2992 ( .B1(n3249), .B2(n3319), .A(n551), .ZN(n1883) );
  OAI21_X2 U2993 ( .B1(n3247), .B2(n3318), .A(n548), .ZN(n1884) );
  OAI21_X2 U2994 ( .B1(n3245), .B2(n3318), .A(n547), .ZN(n1885) );
  OAI21_X2 U2995 ( .B1(n3243), .B2(n3318), .A(n546), .ZN(n1886) );
  OAI21_X2 U2996 ( .B1(n3241), .B2(n3318), .A(n545), .ZN(n1887) );
  OAI21_X2 U2997 ( .B1(n3239), .B2(n3318), .A(n544), .ZN(n1888) );
  OAI21_X2 U2998 ( .B1(n3237), .B2(n3318), .A(n543), .ZN(n1889) );
  OAI21_X2 U2999 ( .B1(n3235), .B2(n3318), .A(n542), .ZN(n1890) );
  OAI21_X2 U3000 ( .B1(n3233), .B2(n3318), .A(n572), .ZN(n1891) );
  OAI21_X2 U3001 ( .B1(n3231), .B2(n3318), .A(n571), .ZN(n1892) );
  OAI21_X2 U3002 ( .B1(n3229), .B2(n3318), .A(n570), .ZN(n1893) );
  OAI21_X2 U3003 ( .B1(n3227), .B2(n3319), .A(n569), .ZN(n1894) );
  OAI21_X2 U3004 ( .B1(n3225), .B2(n3319), .A(n568), .ZN(n1895) );
  OAI21_X2 U3005 ( .B1(n3223), .B2(n3319), .A(n567), .ZN(n1896) );
  OAI21_X2 U3006 ( .B1(n3221), .B2(n541), .A(n566), .ZN(n1897) );
  OAI21_X2 U3007 ( .B1(n3219), .B2(n3320), .A(n565), .ZN(n1898) );
  OAI21_X2 U3008 ( .B1(n3217), .B2(n541), .A(n564), .ZN(n1899) );
  OAI21_X2 U3009 ( .B1(n3215), .B2(n541), .A(n563), .ZN(n1900) );
  OAI21_X2 U3010 ( .B1(n3213), .B2(n3318), .A(n561), .ZN(n1901) );
  OAI21_X2 U3011 ( .B1(n3211), .B2(n3319), .A(n560), .ZN(n1902) );
  OAI21_X2 U3012 ( .B1(n3209), .B2(n541), .A(n559), .ZN(n1903) );
  OAI21_X2 U3013 ( .B1(n3207), .B2(n541), .A(n558), .ZN(n1904) );
  OAI21_X2 U3014 ( .B1(n3205), .B2(n3319), .A(n557), .ZN(n1905) );
  OAI21_X2 U3015 ( .B1(n3203), .B2(n3319), .A(n556), .ZN(n1906) );
  OAI21_X2 U3016 ( .B1(n3201), .B2(n3319), .A(n555), .ZN(n1907) );
  OAI21_X2 U3017 ( .B1(n3199), .B2(n3319), .A(n554), .ZN(n1908) );
  OAI21_X2 U3018 ( .B1(n3197), .B2(n3319), .A(n553), .ZN(n1909) );
  OAI21_X2 U3019 ( .B1(n3195), .B2(n3319), .A(n552), .ZN(n1910) );
  OAI21_X2 U3020 ( .B1(n3193), .B2(n3319), .A(n550), .ZN(n1911) );
  OAI21_X2 U3021 ( .B1(n3191), .B2(n3318), .A(n549), .ZN(n1912) );
  OAI21_X2 U3022 ( .B1(n3253), .B2(n3322), .A(n540), .ZN(n1913) );
  OAI21_X2 U3023 ( .B1(n3251), .B2(n3323), .A(n529), .ZN(n1914) );
  OAI21_X2 U3024 ( .B1(n3249), .B2(n3323), .A(n518), .ZN(n1915) );
  OAI21_X2 U3025 ( .B1(n3247), .B2(n3322), .A(n515), .ZN(n1916) );
  OAI21_X2 U3026 ( .B1(n3245), .B2(n3322), .A(n514), .ZN(n1917) );
  OAI21_X2 U3027 ( .B1(n3243), .B2(n3322), .A(n513), .ZN(n1918) );
  OAI21_X2 U3028 ( .B1(n3241), .B2(n3322), .A(n512), .ZN(n1919) );
  OAI21_X2 U3029 ( .B1(n3239), .B2(n3322), .A(n511), .ZN(n1920) );
  OAI21_X2 U3030 ( .B1(n3237), .B2(n3322), .A(n510), .ZN(n1921) );
  OAI21_X2 U3031 ( .B1(n3235), .B2(n3322), .A(n509), .ZN(n1922) );
  OAI21_X2 U3032 ( .B1(n3233), .B2(n3322), .A(n539), .ZN(n1923) );
  OAI21_X2 U3033 ( .B1(n3231), .B2(n3322), .A(n538), .ZN(n1924) );
  OAI21_X2 U3034 ( .B1(n3229), .B2(n3322), .A(n537), .ZN(n1925) );
  OAI21_X2 U3035 ( .B1(n3227), .B2(n3323), .A(n536), .ZN(n1926) );
  OAI21_X2 U3036 ( .B1(n3225), .B2(n3323), .A(n535), .ZN(n1927) );
  OAI21_X2 U3037 ( .B1(n3223), .B2(n3323), .A(n534), .ZN(n1928) );
  OAI21_X2 U3038 ( .B1(n3221), .B2(n508), .A(n533), .ZN(n1929) );
  OAI21_X2 U3039 ( .B1(n3219), .B2(n3324), .A(n532), .ZN(n1930) );
  OAI21_X2 U3040 ( .B1(n3217), .B2(n508), .A(n531), .ZN(n1931) );
  OAI21_X2 U3041 ( .B1(n3215), .B2(n508), .A(n530), .ZN(n1932) );
  OAI21_X2 U3042 ( .B1(n3213), .B2(n3322), .A(n528), .ZN(n1933) );
  OAI21_X2 U3043 ( .B1(n3211), .B2(n3323), .A(n527), .ZN(n1934) );
  OAI21_X2 U3044 ( .B1(n3209), .B2(n508), .A(n526), .ZN(n1935) );
  OAI21_X2 U3045 ( .B1(n3207), .B2(n508), .A(n525), .ZN(n1936) );
  OAI21_X2 U3046 ( .B1(n3205), .B2(n3323), .A(n524), .ZN(n1937) );
  OAI21_X2 U3047 ( .B1(n3203), .B2(n3323), .A(n523), .ZN(n1938) );
  OAI21_X2 U3048 ( .B1(n3201), .B2(n3323), .A(n522), .ZN(n1939) );
  OAI21_X2 U3049 ( .B1(n3199), .B2(n3323), .A(n521), .ZN(n1940) );
  OAI21_X2 U3050 ( .B1(n3197), .B2(n3323), .A(n520), .ZN(n1941) );
  OAI21_X2 U3051 ( .B1(n3195), .B2(n3323), .A(n519), .ZN(n1942) );
  OAI21_X2 U3052 ( .B1(n3193), .B2(n3323), .A(n517), .ZN(n1943) );
  OAI21_X2 U3053 ( .B1(n3191), .B2(n3322), .A(n516), .ZN(n1944) );
  OAI21_X2 U3054 ( .B1(n3253), .B2(n3327), .A(n507), .ZN(n1945) );
  OAI21_X2 U3055 ( .B1(n3251), .B2(n3327), .A(n496), .ZN(n1946) );
  OAI21_X2 U3056 ( .B1(n3249), .B2(n3328), .A(n485), .ZN(n1947) );
  OAI21_X2 U3057 ( .B1(n3247), .B2(n3327), .A(n482), .ZN(n1948) );
  OAI21_X2 U3058 ( .B1(n3245), .B2(n3327), .A(n481), .ZN(n1949) );
  OAI21_X2 U3059 ( .B1(n3243), .B2(n3327), .A(n480), .ZN(n1950) );
  OAI21_X2 U3060 ( .B1(n3241), .B2(n3327), .A(n479), .ZN(n1951) );
  OAI21_X2 U3061 ( .B1(n3239), .B2(n3327), .A(n478), .ZN(n1952) );
  OAI21_X2 U3062 ( .B1(n3237), .B2(n3327), .A(n477), .ZN(n1953) );
  OAI21_X2 U3063 ( .B1(n3235), .B2(n3327), .A(n476), .ZN(n1954) );
  OAI21_X2 U3064 ( .B1(n3233), .B2(n3327), .A(n506), .ZN(n1955) );
  OAI21_X2 U3065 ( .B1(n3231), .B2(n3327), .A(n505), .ZN(n1956) );
  OAI21_X2 U3066 ( .B1(n3229), .B2(n3327), .A(n504), .ZN(n1957) );
  OAI21_X2 U3067 ( .B1(n3227), .B2(n3328), .A(n503), .ZN(n1958) );
  OAI21_X2 U3068 ( .B1(n3225), .B2(n3328), .A(n502), .ZN(n1959) );
  OAI21_X2 U3069 ( .B1(n3223), .B2(n3328), .A(n501), .ZN(n1960) );
  OAI21_X2 U3070 ( .B1(n3221), .B2(n475), .A(n500), .ZN(n1961) );
  OAI21_X2 U3071 ( .B1(n3219), .B2(n3328), .A(n499), .ZN(n1962) );
  OAI21_X2 U3072 ( .B1(n3217), .B2(n475), .A(n498), .ZN(n1963) );
  OAI21_X2 U3073 ( .B1(n3215), .B2(n475), .A(n497), .ZN(n1964) );
  OAI21_X2 U3074 ( .B1(n3213), .B2(n3329), .A(n495), .ZN(n1965) );
  OAI21_X2 U3075 ( .B1(n3211), .B2(n3328), .A(n494), .ZN(n1966) );
  OAI21_X2 U3076 ( .B1(n3209), .B2(n475), .A(n493), .ZN(n1967) );
  OAI21_X2 U3077 ( .B1(n3207), .B2(n475), .A(n492), .ZN(n1968) );
  OAI21_X2 U3078 ( .B1(n3205), .B2(n3328), .A(n491), .ZN(n1969) );
  OAI21_X2 U3079 ( .B1(n3203), .B2(n3328), .A(n490), .ZN(n1970) );
  OAI21_X2 U3080 ( .B1(n3201), .B2(n3328), .A(n489), .ZN(n1971) );
  OAI21_X2 U3081 ( .B1(n3199), .B2(n3328), .A(n488), .ZN(n1972) );
  OAI21_X2 U3082 ( .B1(n3197), .B2(n3328), .A(n487), .ZN(n1973) );
  OAI21_X2 U3083 ( .B1(n3195), .B2(n3328), .A(n486), .ZN(n1974) );
  OAI21_X2 U3084 ( .B1(n3193), .B2(n3328), .A(n484), .ZN(n1975) );
  OAI21_X2 U3085 ( .B1(n3191), .B2(n3327), .A(n483), .ZN(n1976) );
  OAI21_X2 U3086 ( .B1(n3253), .B2(n3331), .A(n473), .ZN(n1977) );
  OAI21_X2 U3087 ( .B1(n3251), .B2(n3331), .A(n462), .ZN(n1978) );
  OAI21_X2 U3088 ( .B1(n3249), .B2(n3332), .A(n451), .ZN(n1979) );
  OAI21_X2 U3089 ( .B1(n3247), .B2(n3331), .A(n448), .ZN(n1980) );
  OAI21_X2 U3090 ( .B1(n3245), .B2(n3331), .A(n447), .ZN(n1981) );
  OAI21_X2 U3091 ( .B1(n3243), .B2(n3331), .A(n446), .ZN(n1982) );
  OAI21_X2 U3092 ( .B1(n3241), .B2(n3331), .A(n445), .ZN(n1983) );
  OAI21_X2 U3093 ( .B1(n3239), .B2(n3331), .A(n444), .ZN(n1984) );
  OAI21_X2 U3094 ( .B1(n3237), .B2(n3331), .A(n443), .ZN(n1985) );
  OAI21_X2 U3095 ( .B1(n3235), .B2(n3331), .A(n442), .ZN(n1986) );
  OAI21_X2 U3096 ( .B1(n3233), .B2(n3331), .A(n472), .ZN(n1987) );
  OAI21_X2 U3097 ( .B1(n3231), .B2(n3331), .A(n471), .ZN(n1988) );
  OAI21_X2 U3098 ( .B1(n3229), .B2(n3331), .A(n470), .ZN(n1989) );
  OAI21_X2 U3099 ( .B1(n3227), .B2(n3332), .A(n469), .ZN(n1990) );
  OAI21_X2 U3100 ( .B1(n3225), .B2(n3332), .A(n468), .ZN(n1991) );
  OAI21_X2 U3101 ( .B1(n3223), .B2(n3332), .A(n467), .ZN(n1992) );
  OAI21_X2 U3102 ( .B1(n3221), .B2(n441), .A(n466), .ZN(n1993) );
  OAI21_X2 U3103 ( .B1(n3219), .B2(n3332), .A(n465), .ZN(n1994) );
  OAI21_X2 U3104 ( .B1(n3217), .B2(n441), .A(n464), .ZN(n1995) );
  OAI21_X2 U3105 ( .B1(n3215), .B2(n441), .A(n463), .ZN(n1996) );
  OAI21_X2 U3106 ( .B1(n3213), .B2(n3333), .A(n461), .ZN(n1997) );
  OAI21_X2 U3107 ( .B1(n3211), .B2(n3332), .A(n460), .ZN(n1998) );
  OAI21_X2 U3108 ( .B1(n3209), .B2(n441), .A(n459), .ZN(n1999) );
  OAI21_X2 U3109 ( .B1(n3207), .B2(n441), .A(n458), .ZN(n2000) );
  OAI21_X2 U3110 ( .B1(n3205), .B2(n3332), .A(n457), .ZN(n2001) );
  OAI21_X2 U3111 ( .B1(n3203), .B2(n3332), .A(n456), .ZN(n2002) );
  OAI21_X2 U3112 ( .B1(n3201), .B2(n3332), .A(n455), .ZN(n2003) );
  OAI21_X2 U3113 ( .B1(n3199), .B2(n3332), .A(n454), .ZN(n2004) );
  OAI21_X2 U3114 ( .B1(n3197), .B2(n3332), .A(n453), .ZN(n2005) );
  OAI21_X2 U3115 ( .B1(n3195), .B2(n3332), .A(n452), .ZN(n2006) );
  OAI21_X2 U3116 ( .B1(n3193), .B2(n3332), .A(n450), .ZN(n2007) );
  OAI21_X2 U3117 ( .B1(n3191), .B2(n3331), .A(n449), .ZN(n2008) );
  OAI21_X2 U3118 ( .B1(n3253), .B2(n3334), .A(n438), .ZN(n2009) );
  OAI21_X2 U3119 ( .B1(n3251), .B2(n3335), .A(n427), .ZN(n2010) );
  OAI21_X2 U3120 ( .B1(n3249), .B2(n3335), .A(n416), .ZN(n2011) );
  OAI21_X2 U3121 ( .B1(n3247), .B2(n3334), .A(n413), .ZN(n2012) );
  OAI21_X2 U3122 ( .B1(n3245), .B2(n3334), .A(n412), .ZN(n2013) );
  OAI21_X2 U3123 ( .B1(n3243), .B2(n3334), .A(n411), .ZN(n2014) );
  OAI21_X2 U3124 ( .B1(n3241), .B2(n3334), .A(n410), .ZN(n2015) );
  OAI21_X2 U3125 ( .B1(n3239), .B2(n3334), .A(n409), .ZN(n2016) );
  OAI21_X2 U3126 ( .B1(n3237), .B2(n3334), .A(n408), .ZN(n2017) );
  OAI21_X2 U3127 ( .B1(n3235), .B2(n3334), .A(n407), .ZN(n2018) );
  OAI21_X2 U3128 ( .B1(n3233), .B2(n3334), .A(n437), .ZN(n2019) );
  OAI21_X2 U3129 ( .B1(n3231), .B2(n3334), .A(n436), .ZN(n2020) );
  OAI21_X2 U3130 ( .B1(n3229), .B2(n3334), .A(n435), .ZN(n2021) );
  OAI21_X2 U3131 ( .B1(n3227), .B2(n3335), .A(n434), .ZN(n2022) );
  OAI21_X2 U3132 ( .B1(n3225), .B2(n3335), .A(n433), .ZN(n2023) );
  OAI21_X2 U3133 ( .B1(n3223), .B2(n3335), .A(n432), .ZN(n2024) );
  OAI21_X2 U3134 ( .B1(n3221), .B2(n406), .A(n431), .ZN(n2025) );
  OAI21_X2 U3135 ( .B1(n3219), .B2(n3336), .A(n430), .ZN(n2026) );
  OAI21_X2 U3136 ( .B1(n3217), .B2(n406), .A(n429), .ZN(n2027) );
  OAI21_X2 U3137 ( .B1(n3215), .B2(n406), .A(n428), .ZN(n2028) );
  OAI21_X2 U3138 ( .B1(n3213), .B2(n3334), .A(n426), .ZN(n2029) );
  OAI21_X2 U3139 ( .B1(n3211), .B2(n3335), .A(n425), .ZN(n2030) );
  OAI21_X2 U3140 ( .B1(n3209), .B2(n406), .A(n424), .ZN(n2031) );
  OAI21_X2 U3141 ( .B1(n3207), .B2(n406), .A(n423), .ZN(n2032) );
  OAI21_X2 U3142 ( .B1(n3205), .B2(n3335), .A(n422), .ZN(n2033) );
  OAI21_X2 U3143 ( .B1(n3203), .B2(n3335), .A(n421), .ZN(n2034) );
  OAI21_X2 U3144 ( .B1(n3201), .B2(n3335), .A(n420), .ZN(n2035) );
  OAI21_X2 U3145 ( .B1(n3199), .B2(n3335), .A(n419), .ZN(n2036) );
  OAI21_X2 U3146 ( .B1(n3197), .B2(n3335), .A(n418), .ZN(n2037) );
  OAI21_X2 U3147 ( .B1(n3195), .B2(n3335), .A(n417), .ZN(n2038) );
  OAI21_X2 U3148 ( .B1(n3193), .B2(n3335), .A(n415), .ZN(n2039) );
  OAI21_X2 U3149 ( .B1(n3191), .B2(n3334), .A(n414), .ZN(n2040) );
  OAI21_X2 U3150 ( .B1(n3253), .B2(n3338), .A(n405), .ZN(n2041) );
  OAI21_X2 U3151 ( .B1(n3251), .B2(n3339), .A(n394), .ZN(n2042) );
  OAI21_X2 U3152 ( .B1(n3249), .B2(n3339), .A(n383), .ZN(n2043) );
  OAI21_X2 U3153 ( .B1(n3247), .B2(n3338), .A(n380), .ZN(n2044) );
  OAI21_X2 U3154 ( .B1(n3245), .B2(n3338), .A(n379), .ZN(n2045) );
  OAI21_X2 U3155 ( .B1(n3243), .B2(n3338), .A(n378), .ZN(n2046) );
  OAI21_X2 U3156 ( .B1(n3241), .B2(n3338), .A(n377), .ZN(n2047) );
  OAI21_X2 U3157 ( .B1(n3239), .B2(n3338), .A(n376), .ZN(n2048) );
  OAI21_X2 U3158 ( .B1(n3237), .B2(n3338), .A(n375), .ZN(n2049) );
  OAI21_X2 U3159 ( .B1(n3235), .B2(n3338), .A(n374), .ZN(n2050) );
  OAI21_X2 U3160 ( .B1(n3233), .B2(n3338), .A(n404), .ZN(n2051) );
  OAI21_X2 U3161 ( .B1(n3231), .B2(n3338), .A(n403), .ZN(n2052) );
  OAI21_X2 U3162 ( .B1(n3229), .B2(n3338), .A(n402), .ZN(n2053) );
  OAI21_X2 U3163 ( .B1(n3227), .B2(n3339), .A(n401), .ZN(n2054) );
  OAI21_X2 U3164 ( .B1(n3225), .B2(n3339), .A(n400), .ZN(n2055) );
  OAI21_X2 U3165 ( .B1(n3223), .B2(n3339), .A(n399), .ZN(n2056) );
  OAI21_X2 U3166 ( .B1(n3221), .B2(n373), .A(n398), .ZN(n2057) );
  OAI21_X2 U3167 ( .B1(n3219), .B2(n3340), .A(n397), .ZN(n2058) );
  OAI21_X2 U3168 ( .B1(n3217), .B2(n373), .A(n396), .ZN(n2059) );
  OAI21_X2 U3169 ( .B1(n3215), .B2(n373), .A(n395), .ZN(n2060) );
  OAI21_X2 U3170 ( .B1(n3213), .B2(n3338), .A(n393), .ZN(n2061) );
  OAI21_X2 U3171 ( .B1(n3211), .B2(n3339), .A(n392), .ZN(n2062) );
  OAI21_X2 U3172 ( .B1(n3209), .B2(n373), .A(n391), .ZN(n2063) );
  OAI21_X2 U3173 ( .B1(n3207), .B2(n373), .A(n390), .ZN(n2064) );
  OAI21_X2 U3174 ( .B1(n3205), .B2(n3339), .A(n389), .ZN(n2065) );
  OAI21_X2 U3175 ( .B1(n3203), .B2(n3339), .A(n388), .ZN(n2066) );
  OAI21_X2 U3176 ( .B1(n3201), .B2(n3339), .A(n387), .ZN(n2067) );
  OAI21_X2 U3177 ( .B1(n3199), .B2(n3339), .A(n386), .ZN(n2068) );
  OAI21_X2 U3178 ( .B1(n3197), .B2(n3339), .A(n385), .ZN(n2069) );
  OAI21_X2 U3179 ( .B1(n3195), .B2(n3339), .A(n384), .ZN(n2070) );
  OAI21_X2 U3180 ( .B1(n3193), .B2(n3339), .A(n382), .ZN(n2071) );
  OAI21_X2 U3181 ( .B1(n3191), .B2(n3338), .A(n381), .ZN(n2072) );
  OAI21_X2 U3182 ( .B1(n3253), .B2(n3347), .A(n339), .ZN(n2073) );
  OAI21_X2 U3183 ( .B1(n3251), .B2(n3347), .A(n328), .ZN(n2074) );
  OAI21_X2 U3184 ( .B1(n3249), .B2(n3348), .A(n317), .ZN(n2075) );
  OAI21_X2 U3185 ( .B1(n3247), .B2(n3347), .A(n314), .ZN(n2076) );
  OAI21_X2 U3186 ( .B1(n3245), .B2(n3347), .A(n313), .ZN(n2077) );
  OAI21_X2 U3187 ( .B1(n3243), .B2(n3347), .A(n312), .ZN(n2078) );
  OAI21_X2 U3188 ( .B1(n3241), .B2(n3347), .A(n311), .ZN(n2079) );
  OAI21_X2 U3189 ( .B1(n3239), .B2(n3347), .A(n310), .ZN(n2080) );
  OAI21_X2 U3190 ( .B1(n3237), .B2(n3347), .A(n309), .ZN(n2081) );
  OAI21_X2 U3191 ( .B1(n3235), .B2(n3347), .A(n308), .ZN(n2082) );
  OAI21_X2 U3192 ( .B1(n3233), .B2(n3347), .A(n338), .ZN(n2083) );
  OAI21_X2 U3193 ( .B1(n3231), .B2(n3347), .A(n337), .ZN(n2084) );
  OAI21_X2 U3194 ( .B1(n3229), .B2(n3347), .A(n336), .ZN(n2085) );
  OAI21_X2 U3195 ( .B1(n3227), .B2(n3348), .A(n335), .ZN(n2086) );
  OAI21_X2 U3196 ( .B1(n3225), .B2(n3348), .A(n334), .ZN(n2087) );
  OAI21_X2 U3197 ( .B1(n3223), .B2(n3348), .A(n333), .ZN(n2088) );
  OAI21_X2 U3198 ( .B1(n3221), .B2(n307), .A(n332), .ZN(n2089) );
  OAI21_X2 U3199 ( .B1(n3219), .B2(n3348), .A(n331), .ZN(n2090) );
  OAI21_X2 U3200 ( .B1(n3217), .B2(n307), .A(n330), .ZN(n2091) );
  OAI21_X2 U3201 ( .B1(n3215), .B2(n307), .A(n329), .ZN(n2092) );
  OAI21_X2 U3202 ( .B1(n3213), .B2(n3349), .A(n327), .ZN(n2093) );
  OAI21_X2 U3203 ( .B1(n3211), .B2(n3348), .A(n326), .ZN(n2094) );
  OAI21_X2 U3204 ( .B1(n3209), .B2(n307), .A(n325), .ZN(n2095) );
  OAI21_X2 U3205 ( .B1(n3207), .B2(n307), .A(n324), .ZN(n2096) );
  OAI21_X2 U3206 ( .B1(n3205), .B2(n3348), .A(n323), .ZN(n2097) );
  OAI21_X2 U3207 ( .B1(n3203), .B2(n3348), .A(n322), .ZN(n2098) );
  OAI21_X2 U3208 ( .B1(n3201), .B2(n3348), .A(n321), .ZN(n2099) );
  OAI21_X2 U3209 ( .B1(n3199), .B2(n3348), .A(n320), .ZN(n2100) );
  OAI21_X2 U3210 ( .B1(n3197), .B2(n3348), .A(n319), .ZN(n2101) );
  OAI21_X2 U3211 ( .B1(n3195), .B2(n3348), .A(n318), .ZN(n2102) );
  OAI21_X2 U3212 ( .B1(n3193), .B2(n3348), .A(n316), .ZN(n2103) );
  OAI21_X2 U3213 ( .B1(n3191), .B2(n3347), .A(n315), .ZN(n2104) );
  OAI21_X2 U3214 ( .B1(n3252), .B2(n3351), .A(n305), .ZN(n2105) );
  OAI21_X2 U3215 ( .B1(n3250), .B2(n3351), .A(n294), .ZN(n2106) );
  OAI21_X2 U3216 ( .B1(n3248), .B2(n3352), .A(n283), .ZN(n2107) );
  OAI21_X2 U3217 ( .B1(n3246), .B2(n3351), .A(n280), .ZN(n2108) );
  OAI21_X2 U3218 ( .B1(n3244), .B2(n3351), .A(n279), .ZN(n2109) );
  OAI21_X2 U3219 ( .B1(n3242), .B2(n3351), .A(n278), .ZN(n2110) );
  OAI21_X2 U3220 ( .B1(n3240), .B2(n3351), .A(n277), .ZN(n2111) );
  OAI21_X2 U3221 ( .B1(n3238), .B2(n3351), .A(n276), .ZN(n2112) );
  OAI21_X2 U3222 ( .B1(n3236), .B2(n3351), .A(n275), .ZN(n2113) );
  OAI21_X2 U3223 ( .B1(n3234), .B2(n3351), .A(n274), .ZN(n2114) );
  OAI21_X2 U3224 ( .B1(n3232), .B2(n3351), .A(n304), .ZN(n2115) );
  OAI21_X2 U3225 ( .B1(n3230), .B2(n3351), .A(n303), .ZN(n2116) );
  OAI21_X2 U3226 ( .B1(n3228), .B2(n3351), .A(n302), .ZN(n2117) );
  OAI21_X2 U3227 ( .B1(n3226), .B2(n3352), .A(n301), .ZN(n2118) );
  OAI21_X2 U3228 ( .B1(n3224), .B2(n3352), .A(n300), .ZN(n2119) );
  OAI21_X2 U3229 ( .B1(n3222), .B2(n3352), .A(n299), .ZN(n2120) );
  OAI21_X2 U3230 ( .B1(n3220), .B2(n273), .A(n298), .ZN(n2121) );
  OAI21_X2 U3231 ( .B1(n3218), .B2(n3352), .A(n297), .ZN(n2122) );
  OAI21_X2 U3232 ( .B1(n3216), .B2(n273), .A(n296), .ZN(n2123) );
  OAI21_X2 U3233 ( .B1(n3214), .B2(n273), .A(n295), .ZN(n2124) );
  OAI21_X2 U3234 ( .B1(n3212), .B2(n3353), .A(n293), .ZN(n2125) );
  OAI21_X2 U3235 ( .B1(n3210), .B2(n3352), .A(n292), .ZN(n2126) );
  OAI21_X2 U3236 ( .B1(n3208), .B2(n273), .A(n291), .ZN(n2127) );
  OAI21_X2 U3237 ( .B1(n3206), .B2(n273), .A(n290), .ZN(n2128) );
  OAI21_X2 U3238 ( .B1(n3204), .B2(n3352), .A(n289), .ZN(n2129) );
  OAI21_X2 U3239 ( .B1(n3202), .B2(n3352), .A(n288), .ZN(n2130) );
  OAI21_X2 U3240 ( .B1(n3200), .B2(n3352), .A(n287), .ZN(n2131) );
  OAI21_X2 U3241 ( .B1(n3198), .B2(n3352), .A(n286), .ZN(n2132) );
  OAI21_X2 U3242 ( .B1(n3196), .B2(n3352), .A(n285), .ZN(n2133) );
  OAI21_X2 U3243 ( .B1(n3194), .B2(n3352), .A(n284), .ZN(n2134) );
  OAI21_X2 U3244 ( .B1(n3192), .B2(n3352), .A(n282), .ZN(n2135) );
  OAI21_X2 U3245 ( .B1(n3190), .B2(n3351), .A(n281), .ZN(n2136) );
  INV_X4 U3246 ( .A(n3184), .ZN(n3172) );
  INV_X4 U3247 ( .A(n3174), .ZN(n3176) );
  INV_X4 U3248 ( .A(n3174), .ZN(n3175) );
  INV_X4 U3249 ( .A(N11), .ZN(n3173) );
  INV_X4 U3250 ( .A(n3173), .ZN(n3177) );
  INV_X4 U3251 ( .A(n3185), .ZN(n3189) );
  INV_X4 U3252 ( .A(n3185), .ZN(n3188) );
  INV_X4 U3253 ( .A(N11), .ZN(n3183) );
  BUF_X4 U3254 ( .A(N9), .Z(n3152) );
  INV_X4 U3255 ( .A(n3174), .ZN(n3180) );
  INV_X4 U3256 ( .A(n3174), .ZN(n3179) );
  INV_X4 U3257 ( .A(n3173), .ZN(n3178) );
  INV_X4 U3258 ( .A(n1046), .ZN(n3258) );
  INV_X4 U3259 ( .A(n1013), .ZN(n3262) );
  INV_X4 U3260 ( .A(n137), .ZN(n3366) );
  INV_X4 U3261 ( .A(n102), .ZN(n3370) );
  INV_X4 U3262 ( .A(n68), .ZN(n3374) );
  INV_X4 U3263 ( .A(n1), .ZN(n3378) );
  INV_X4 U3264 ( .A(n912), .ZN(n3274) );
  INV_X4 U3265 ( .A(n878), .ZN(n3278) );
  INV_X4 U3266 ( .A(n776), .ZN(n3290) );
  INV_X4 U3267 ( .A(n742), .ZN(n3294) );
  INV_X4 U3268 ( .A(n609), .ZN(n3310) );
  INV_X4 U3269 ( .A(n575), .ZN(n3314) );
  INV_X4 U3270 ( .A(n475), .ZN(n3326) );
  INV_X4 U3271 ( .A(n441), .ZN(n3330) );
  INV_X4 U3272 ( .A(n340), .ZN(n3342) );
  INV_X4 U3273 ( .A(n307), .ZN(n3346) );
  INV_X4 U3274 ( .A(n273), .ZN(n3350) );
  INV_X4 U3275 ( .A(n239), .ZN(n3354) );
  INV_X4 U3276 ( .A(N12), .ZN(n3185) );
  INV_X4 U3277 ( .A(n3185), .ZN(n3187) );
  INV_X4 U3278 ( .A(n3185), .ZN(n3186) );
  INV_X4 U3279 ( .A(N11), .ZN(n3174) );
  INV_X4 U3280 ( .A(n3183), .ZN(n3184) );
  INV_X4 U3281 ( .A(n1079), .ZN(n3257) );
  INV_X4 U3282 ( .A(n3257), .ZN(n3254) );
  INV_X4 U3283 ( .A(n3257), .ZN(n3255) );
  INV_X4 U3284 ( .A(n3257), .ZN(n3256) );
  INV_X4 U3285 ( .A(n3258), .ZN(n3259) );
  INV_X4 U3286 ( .A(n3258), .ZN(n3260) );
  INV_X4 U3287 ( .A(n3258), .ZN(n3261) );
  INV_X4 U3288 ( .A(n3262), .ZN(n3263) );
  INV_X4 U3289 ( .A(n3262), .ZN(n3264) );
  INV_X4 U3290 ( .A(n3262), .ZN(n3265) );
  INV_X4 U3291 ( .A(n979), .ZN(n3269) );
  INV_X4 U3292 ( .A(n3269), .ZN(n3266) );
  INV_X4 U3293 ( .A(n3269), .ZN(n3267) );
  INV_X4 U3294 ( .A(n3269), .ZN(n3268) );
  INV_X4 U3295 ( .A(n945), .ZN(n3273) );
  INV_X4 U3296 ( .A(n3273), .ZN(n3270) );
  INV_X4 U3297 ( .A(n3273), .ZN(n3271) );
  INV_X4 U3298 ( .A(n3273), .ZN(n3272) );
  INV_X4 U3299 ( .A(n3274), .ZN(n3275) );
  INV_X4 U3300 ( .A(n3274), .ZN(n3276) );
  INV_X4 U3301 ( .A(n3274), .ZN(n3277) );
  INV_X4 U3302 ( .A(n3278), .ZN(n3279) );
  INV_X4 U3303 ( .A(n3278), .ZN(n3280) );
  INV_X4 U3304 ( .A(n3278), .ZN(n3281) );
  INV_X4 U3305 ( .A(n842), .ZN(n3285) );
  INV_X4 U3306 ( .A(n3285), .ZN(n3282) );
  INV_X4 U3307 ( .A(n3285), .ZN(n3283) );
  INV_X4 U3308 ( .A(n3285), .ZN(n3284) );
  INV_X4 U3309 ( .A(n809), .ZN(n3289) );
  INV_X4 U3310 ( .A(n3289), .ZN(n3286) );
  INV_X4 U3311 ( .A(n3289), .ZN(n3287) );
  INV_X4 U3312 ( .A(n3289), .ZN(n3288) );
  INV_X4 U3313 ( .A(n3290), .ZN(n3291) );
  INV_X4 U3314 ( .A(n3290), .ZN(n3292) );
  INV_X4 U3315 ( .A(n3290), .ZN(n3293) );
  INV_X4 U3316 ( .A(n3294), .ZN(n3295) );
  INV_X4 U3317 ( .A(n3294), .ZN(n3296) );
  INV_X4 U3318 ( .A(n3294), .ZN(n3297) );
  INV_X4 U3319 ( .A(n709), .ZN(n3301) );
  INV_X4 U3320 ( .A(n3301), .ZN(n3298) );
  INV_X4 U3321 ( .A(n3301), .ZN(n3299) );
  INV_X4 U3322 ( .A(n3301), .ZN(n3300) );
  INV_X4 U3323 ( .A(n675), .ZN(n3305) );
  INV_X4 U3324 ( .A(n3305), .ZN(n3302) );
  INV_X4 U3325 ( .A(n3305), .ZN(n3303) );
  INV_X4 U3326 ( .A(n3305), .ZN(n3304) );
  INV_X4 U3327 ( .A(n642), .ZN(n3309) );
  INV_X4 U3328 ( .A(n3309), .ZN(n3306) );
  INV_X4 U3329 ( .A(n3309), .ZN(n3307) );
  INV_X4 U3330 ( .A(n3309), .ZN(n3308) );
  INV_X4 U3331 ( .A(n3310), .ZN(n3311) );
  INV_X4 U3332 ( .A(n3310), .ZN(n3312) );
  INV_X4 U3333 ( .A(n3310), .ZN(n3313) );
  INV_X4 U3334 ( .A(n3314), .ZN(n3315) );
  INV_X4 U3335 ( .A(n3314), .ZN(n3316) );
  INV_X4 U3336 ( .A(n3314), .ZN(n3317) );
  INV_X4 U3337 ( .A(n541), .ZN(n3321) );
  INV_X4 U3338 ( .A(n3321), .ZN(n3318) );
  INV_X4 U3339 ( .A(n3321), .ZN(n3319) );
  INV_X4 U3340 ( .A(n3321), .ZN(n3320) );
  INV_X4 U3341 ( .A(n508), .ZN(n3325) );
  INV_X4 U3342 ( .A(n3325), .ZN(n3322) );
  INV_X4 U3343 ( .A(n3325), .ZN(n3323) );
  INV_X4 U3344 ( .A(n3325), .ZN(n3324) );
  INV_X4 U3345 ( .A(n3326), .ZN(n3327) );
  INV_X4 U3346 ( .A(n3326), .ZN(n3328) );
  INV_X4 U3347 ( .A(n3326), .ZN(n3329) );
  INV_X4 U3348 ( .A(n3330), .ZN(n3331) );
  INV_X4 U3349 ( .A(n3330), .ZN(n3332) );
  INV_X4 U3350 ( .A(n3330), .ZN(n3333) );
  INV_X4 U3351 ( .A(n406), .ZN(n3337) );
  INV_X4 U3352 ( .A(n3337), .ZN(n3334) );
  INV_X4 U3353 ( .A(n3337), .ZN(n3335) );
  INV_X4 U3354 ( .A(n3337), .ZN(n3336) );
  INV_X4 U3355 ( .A(n373), .ZN(n3341) );
  INV_X4 U3356 ( .A(n3341), .ZN(n3338) );
  INV_X4 U3357 ( .A(n3341), .ZN(n3339) );
  INV_X4 U3358 ( .A(n3341), .ZN(n3340) );
  INV_X4 U3359 ( .A(n3342), .ZN(n3343) );
  INV_X4 U3360 ( .A(n3342), .ZN(n3344) );
  INV_X4 U3361 ( .A(n3342), .ZN(n3345) );
  INV_X4 U3362 ( .A(n3346), .ZN(n3347) );
  INV_X4 U3363 ( .A(n3346), .ZN(n3348) );
  INV_X4 U3364 ( .A(n3346), .ZN(n3349) );
  INV_X4 U3365 ( .A(n3350), .ZN(n3351) );
  INV_X4 U3366 ( .A(n3350), .ZN(n3352) );
  INV_X4 U3367 ( .A(n3350), .ZN(n3353) );
  INV_X4 U3368 ( .A(n3354), .ZN(n3355) );
  INV_X4 U3369 ( .A(n3354), .ZN(n3356) );
  INV_X4 U3370 ( .A(n3354), .ZN(n3357) );
  INV_X4 U3371 ( .A(n204), .ZN(n3361) );
  INV_X4 U3372 ( .A(n3361), .ZN(n3358) );
  INV_X4 U3373 ( .A(n3361), .ZN(n3359) );
  INV_X4 U3374 ( .A(n3361), .ZN(n3360) );
  INV_X4 U3375 ( .A(n171), .ZN(n3365) );
  INV_X4 U3376 ( .A(n3365), .ZN(n3362) );
  INV_X4 U3377 ( .A(n3365), .ZN(n3363) );
  INV_X4 U3378 ( .A(n3365), .ZN(n3364) );
  INV_X4 U3379 ( .A(n3366), .ZN(n3367) );
  INV_X4 U3380 ( .A(n3366), .ZN(n3368) );
  INV_X4 U3381 ( .A(n3366), .ZN(n3369) );
  INV_X4 U3382 ( .A(n3370), .ZN(n3371) );
  INV_X4 U3383 ( .A(n3370), .ZN(n3372) );
  INV_X4 U3384 ( .A(n3370), .ZN(n3373) );
  INV_X4 U3385 ( .A(n3374), .ZN(n3375) );
  INV_X4 U3386 ( .A(n3374), .ZN(n3376) );
  INV_X4 U3387 ( .A(n3374), .ZN(n3377) );
  INV_X4 U3388 ( .A(n3378), .ZN(n3379) );
  INV_X4 U3389 ( .A(n3378), .ZN(n3380) );
  INV_X4 U3390 ( .A(n3378), .ZN(n3381) );
  INV_X4 U3391 ( .A(wData[0]), .ZN(n3252) );
  INV_X4 U3392 ( .A(wData[0]), .ZN(n3253) );
  INV_X4 U3393 ( .A(wData[10]), .ZN(n3232) );
  INV_X4 U3394 ( .A(wData[10]), .ZN(n3233) );
  INV_X4 U3395 ( .A(wData[11]), .ZN(n3230) );
  INV_X4 U3396 ( .A(wData[11]), .ZN(n3231) );
  INV_X4 U3397 ( .A(wData[12]), .ZN(n3228) );
  INV_X4 U3398 ( .A(wData[12]), .ZN(n3229) );
  INV_X4 U3399 ( .A(wData[13]), .ZN(n3226) );
  INV_X4 U3400 ( .A(wData[13]), .ZN(n3227) );
  INV_X4 U3401 ( .A(wData[14]), .ZN(n3224) );
  INV_X4 U3402 ( .A(wData[14]), .ZN(n3225) );
  INV_X4 U3403 ( .A(wData[15]), .ZN(n3222) );
  INV_X4 U3404 ( .A(wData[15]), .ZN(n3223) );
  INV_X4 U3405 ( .A(wData[16]), .ZN(n3220) );
  INV_X4 U3406 ( .A(wData[16]), .ZN(n3221) );
  INV_X4 U3407 ( .A(wData[17]), .ZN(n3218) );
  INV_X4 U3408 ( .A(wData[17]), .ZN(n3219) );
  INV_X4 U3409 ( .A(wData[18]), .ZN(n3216) );
  INV_X4 U3410 ( .A(wData[18]), .ZN(n3217) );
  INV_X4 U3411 ( .A(wData[19]), .ZN(n3214) );
  INV_X4 U3412 ( .A(wData[19]), .ZN(n3215) );
  INV_X4 U3413 ( .A(wData[1]), .ZN(n3250) );
  INV_X4 U3414 ( .A(wData[1]), .ZN(n3251) );
  INV_X4 U3415 ( .A(wData[20]), .ZN(n3212) );
  INV_X4 U3416 ( .A(wData[20]), .ZN(n3213) );
  INV_X4 U3417 ( .A(wData[21]), .ZN(n3210) );
  INV_X4 U3418 ( .A(wData[21]), .ZN(n3211) );
  INV_X4 U3419 ( .A(wData[22]), .ZN(n3208) );
  INV_X4 U3420 ( .A(wData[22]), .ZN(n3209) );
  INV_X4 U3421 ( .A(wData[23]), .ZN(n3206) );
  INV_X4 U3422 ( .A(wData[23]), .ZN(n3207) );
  INV_X4 U3423 ( .A(wData[24]), .ZN(n3204) );
  INV_X4 U3424 ( .A(wData[24]), .ZN(n3205) );
  INV_X4 U3425 ( .A(wData[25]), .ZN(n3202) );
  INV_X4 U3426 ( .A(wData[25]), .ZN(n3203) );
  INV_X4 U3427 ( .A(wData[26]), .ZN(n3200) );
  INV_X4 U3428 ( .A(wData[26]), .ZN(n3201) );
  INV_X4 U3429 ( .A(wData[27]), .ZN(n3198) );
  INV_X4 U3430 ( .A(wData[27]), .ZN(n3199) );
  INV_X4 U3431 ( .A(wData[28]), .ZN(n3196) );
  INV_X4 U3432 ( .A(wData[28]), .ZN(n3197) );
  INV_X4 U3433 ( .A(wData[29]), .ZN(n3194) );
  INV_X4 U3434 ( .A(wData[29]), .ZN(n3195) );
  INV_X4 U3435 ( .A(wData[2]), .ZN(n3248) );
  INV_X4 U3436 ( .A(wData[2]), .ZN(n3249) );
  INV_X4 U3437 ( .A(wData[30]), .ZN(n3192) );
  INV_X4 U3438 ( .A(wData[30]), .ZN(n3193) );
  INV_X4 U3439 ( .A(wData[31]), .ZN(n3190) );
  INV_X4 U3440 ( .A(wData[31]), .ZN(n3191) );
  INV_X4 U3441 ( .A(wData[3]), .ZN(n3246) );
  INV_X4 U3442 ( .A(wData[3]), .ZN(n3247) );
  INV_X4 U3443 ( .A(wData[4]), .ZN(n3244) );
  INV_X4 U3444 ( .A(wData[4]), .ZN(n3245) );
  INV_X4 U3445 ( .A(wData[5]), .ZN(n3242) );
  INV_X4 U3446 ( .A(wData[5]), .ZN(n3243) );
  INV_X4 U3447 ( .A(wData[6]), .ZN(n3240) );
  INV_X4 U3448 ( .A(wData[6]), .ZN(n3241) );
  INV_X4 U3449 ( .A(wData[7]), .ZN(n3238) );
  INV_X4 U3450 ( .A(wData[7]), .ZN(n3239) );
  INV_X4 U3451 ( .A(wData[8]), .ZN(n3236) );
  INV_X4 U3452 ( .A(wData[8]), .ZN(n3237) );
  INV_X4 U3453 ( .A(wData[9]), .ZN(n3234) );
  INV_X4 U3454 ( .A(wData[9]), .ZN(n3235) );
  MUX2_X2 U3455 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n3107), .Z(n2137) );
  MUX2_X2 U3456 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n3107), .Z(n2138) );
  MUX2_X2 U3457 ( .A(n2138), .B(n2137), .S(N10), .Z(n2139) );
  MUX2_X2 U3458 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n3107), .Z(n2140) );
  MUX2_X2 U3459 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n3107), .Z(n2141) );
  MUX2_X2 U3460 ( .A(n2141), .B(n2140), .S(N10), .Z(n2142) );
  MUX2_X2 U3461 ( .A(n2142), .B(n2139), .S(n3184), .Z(n2143) );
  MUX2_X2 U3462 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n3107), .Z(n2144) );
  MUX2_X2 U3463 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n3107), .Z(n2145) );
  MUX2_X2 U3464 ( .A(n2145), .B(n2144), .S(N10), .Z(n2146) );
  MUX2_X2 U3465 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n3108), .Z(n2147) );
  MUX2_X2 U3466 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n3108), .Z(n2148) );
  MUX2_X2 U3467 ( .A(n2148), .B(n2147), .S(n3154), .Z(n2149) );
  MUX2_X2 U3468 ( .A(n2149), .B(n2146), .S(n3184), .Z(n2150) );
  MUX2_X2 U3469 ( .A(n2150), .B(n2143), .S(n3187), .Z(n2151) );
  MUX2_X2 U3470 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n3108), .Z(n2152) );
  MUX2_X2 U3471 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n3108), .Z(n2153) );
  MUX2_X2 U3472 ( .A(n2153), .B(n2152), .S(n3154), .Z(n2154) );
  MUX2_X2 U3473 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n3108), .Z(n2155) );
  MUX2_X2 U3474 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n3108), .Z(n2156) );
  MUX2_X2 U3475 ( .A(n2156), .B(n2155), .S(n3154), .Z(n2157) );
  MUX2_X2 U3476 ( .A(n2157), .B(n2154), .S(n3184), .Z(n2158) );
  MUX2_X2 U3477 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n3108), .Z(n2159) );
  MUX2_X2 U3478 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n3108), .Z(n2160) );
  MUX2_X2 U3479 ( .A(n2160), .B(n2159), .S(n3154), .Z(n2161) );
  MUX2_X2 U3480 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n3108), .Z(n2162) );
  MUX2_X2 U3481 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n3108), .Z(n2163) );
  MUX2_X2 U3482 ( .A(n2163), .B(n2162), .S(n3154), .Z(n2164) );
  MUX2_X2 U3483 ( .A(n2164), .B(n2161), .S(n3184), .Z(n2165) );
  MUX2_X2 U3484 ( .A(n2165), .B(n2158), .S(n3186), .Z(n2166) );
  MUX2_X2 U3485 ( .A(n2166), .B(n2151), .S(N13), .Z(rData[0]) );
  MUX2_X2 U3486 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n3108), .Z(n2167) );
  MUX2_X2 U3487 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n3109), .Z(n2168) );
  MUX2_X2 U3488 ( .A(n2168), .B(n2167), .S(n3154), .Z(n2169) );
  MUX2_X2 U3489 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n3109), .Z(n2170) );
  MUX2_X2 U3490 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n3109), .Z(n2171) );
  MUX2_X2 U3491 ( .A(n2171), .B(n2170), .S(n3154), .Z(n2172) );
  MUX2_X2 U3492 ( .A(n2172), .B(n2169), .S(n3184), .Z(n2173) );
  MUX2_X2 U3493 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n3109), .Z(n2174) );
  MUX2_X2 U3494 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n3109), .Z(n2175) );
  MUX2_X2 U3495 ( .A(n2175), .B(n2174), .S(n3154), .Z(n2176) );
  MUX2_X2 U3496 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n3109), .Z(n2177) );
  MUX2_X2 U3497 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n3109), .Z(n2178) );
  MUX2_X2 U3498 ( .A(n2178), .B(n2177), .S(n3154), .Z(n2179) );
  MUX2_X2 U3499 ( .A(n2179), .B(n2176), .S(n3184), .Z(n2180) );
  MUX2_X2 U3500 ( .A(n2180), .B(n2173), .S(n3186), .Z(n2181) );
  MUX2_X2 U3501 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n3109), .Z(n2182) );
  MUX2_X2 U3502 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n3109), .Z(n2183) );
  MUX2_X2 U3503 ( .A(n2183), .B(n2182), .S(n3154), .Z(n2184) );
  MUX2_X2 U3504 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n3109), .Z(n2185) );
  MUX2_X2 U3505 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n3109), .Z(n2186) );
  MUX2_X2 U3506 ( .A(n2186), .B(n2185), .S(n3154), .Z(n2187) );
  MUX2_X2 U3507 ( .A(n2187), .B(n2184), .S(n3184), .Z(n2188) );
  MUX2_X2 U3508 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n3110), .Z(n2189) );
  MUX2_X2 U3509 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n3110), .Z(n2190) );
  MUX2_X2 U3510 ( .A(n2190), .B(n2189), .S(n3155), .Z(n2191) );
  MUX2_X2 U3511 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n3110), .Z(n2192) );
  MUX2_X2 U3512 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n3110), .Z(n2193) );
  MUX2_X2 U3513 ( .A(n2193), .B(n2192), .S(n3155), .Z(n2194) );
  MUX2_X2 U3514 ( .A(n2194), .B(n2191), .S(n3175), .Z(n2195) );
  MUX2_X2 U3515 ( .A(n2195), .B(n2188), .S(N12), .Z(n2196) );
  MUX2_X2 U3516 ( .A(n2196), .B(n2181), .S(N13), .Z(rData[1]) );
  MUX2_X2 U3517 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n3110), .Z(n2197) );
  MUX2_X2 U3518 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n3110), .Z(n2198) );
  MUX2_X2 U3519 ( .A(n2198), .B(n2197), .S(n3155), .Z(n2199) );
  MUX2_X2 U3520 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n3110), .Z(n2200) );
  MUX2_X2 U3521 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n3110), .Z(n2201) );
  MUX2_X2 U3522 ( .A(n2201), .B(n2200), .S(n3155), .Z(n2202) );
  MUX2_X2 U3523 ( .A(n2202), .B(n2199), .S(n3175), .Z(n2203) );
  MUX2_X2 U3524 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n3110), .Z(n2204) );
  MUX2_X2 U3525 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n3110), .Z(n2205) );
  MUX2_X2 U3526 ( .A(n2205), .B(n2204), .S(n3155), .Z(n2206) );
  MUX2_X2 U3527 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n3110), .Z(n2207) );
  MUX2_X2 U3528 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n3111), .Z(n2208) );
  MUX2_X2 U3529 ( .A(n2208), .B(n2207), .S(n3155), .Z(n2209) );
  MUX2_X2 U3530 ( .A(n2209), .B(n2206), .S(n3175), .Z(n2210) );
  MUX2_X2 U3531 ( .A(n2210), .B(n2203), .S(n3187), .Z(n2211) );
  MUX2_X2 U3532 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n3111), .Z(n2212) );
  MUX2_X2 U3533 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n3111), .Z(n2213) );
  MUX2_X2 U3534 ( .A(n2213), .B(n2212), .S(n3155), .Z(n2214) );
  MUX2_X2 U3535 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n3111), .Z(n2215) );
  MUX2_X2 U3536 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n3111), .Z(n2216) );
  MUX2_X2 U3537 ( .A(n2216), .B(n2215), .S(n3155), .Z(n2217) );
  MUX2_X2 U3538 ( .A(n2217), .B(n2214), .S(n3175), .Z(n2218) );
  MUX2_X2 U3539 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n3111), .Z(n2219) );
  MUX2_X2 U3540 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n3111), .Z(n2220) );
  MUX2_X2 U3541 ( .A(n2220), .B(n2219), .S(n3155), .Z(n2221) );
  MUX2_X2 U3542 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n3111), .Z(n2222) );
  MUX2_X2 U3543 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n3111), .Z(n2223) );
  MUX2_X2 U3544 ( .A(n2223), .B(n2222), .S(n3155), .Z(n2224) );
  MUX2_X2 U3545 ( .A(n2224), .B(n2221), .S(n3175), .Z(n2225) );
  MUX2_X2 U3546 ( .A(n2225), .B(n2218), .S(N12), .Z(n2226) );
  MUX2_X2 U3547 ( .A(n2226), .B(n2211), .S(N13), .Z(rData[2]) );
  MUX2_X2 U3548 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n3111), .Z(n2227) );
  MUX2_X2 U3549 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n3111), .Z(n2228) );
  MUX2_X2 U3550 ( .A(n2228), .B(n2227), .S(n3155), .Z(n2229) );
  MUX2_X2 U3551 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n3112), .Z(n2230) );
  MUX2_X2 U3552 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n3112), .Z(n2231) );
  MUX2_X2 U3553 ( .A(n2231), .B(n2230), .S(n3156), .Z(n2232) );
  MUX2_X2 U3554 ( .A(n2232), .B(n2229), .S(n3175), .Z(n2233) );
  MUX2_X2 U3555 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n3112), .Z(n2234) );
  MUX2_X2 U3556 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n3112), .Z(n2235) );
  MUX2_X2 U3557 ( .A(n2235), .B(n2234), .S(n3156), .Z(n2236) );
  MUX2_X2 U3558 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n3112), .Z(n2237) );
  MUX2_X2 U3559 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n3112), .Z(n2238) );
  MUX2_X2 U3560 ( .A(n2238), .B(n2237), .S(n3156), .Z(n2239) );
  MUX2_X2 U3561 ( .A(n2239), .B(n2236), .S(n3175), .Z(n2240) );
  MUX2_X2 U3562 ( .A(n2240), .B(n2233), .S(n3186), .Z(n2241) );
  MUX2_X2 U3563 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n3112), .Z(n2242) );
  MUX2_X2 U3564 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n3112), .Z(n2243) );
  MUX2_X2 U3565 ( .A(n2243), .B(n2242), .S(n3156), .Z(n2244) );
  MUX2_X2 U3566 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n3112), .Z(n2245) );
  MUX2_X2 U3567 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n3112), .Z(n2246) );
  MUX2_X2 U3568 ( .A(n2246), .B(n2245), .S(n3156), .Z(n2247) );
  MUX2_X2 U3569 ( .A(n2247), .B(n2244), .S(n3175), .Z(n2248) );
  MUX2_X2 U3570 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n3112), .Z(n2249) );
  MUX2_X2 U3571 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n3113), .Z(n2250) );
  MUX2_X2 U3572 ( .A(n2250), .B(n2249), .S(n3156), .Z(n2251) );
  MUX2_X2 U3573 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n3113), .Z(n2252) );
  MUX2_X2 U3574 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n3113), .Z(n2253) );
  MUX2_X2 U3575 ( .A(n2253), .B(n2252), .S(n3156), .Z(n2254) );
  MUX2_X2 U3576 ( .A(n2254), .B(n2251), .S(n3175), .Z(n2255) );
  MUX2_X2 U3577 ( .A(n2255), .B(n2248), .S(N12), .Z(n2256) );
  MUX2_X2 U3578 ( .A(n2256), .B(n2241), .S(N13), .Z(rData[3]) );
  MUX2_X2 U3579 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n3113), .Z(n2257) );
  MUX2_X2 U3580 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n3113), .Z(n2258) );
  MUX2_X2 U3581 ( .A(n2258), .B(n2257), .S(n3156), .Z(n2259) );
  MUX2_X2 U3582 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n3113), .Z(n2260) );
  MUX2_X2 U3583 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n3113), .Z(n2261) );
  MUX2_X2 U3584 ( .A(n2261), .B(n2260), .S(n3156), .Z(n2262) );
  MUX2_X2 U3585 ( .A(n2262), .B(n2259), .S(n3175), .Z(n2263) );
  MUX2_X2 U3586 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n3113), .Z(n2264) );
  MUX2_X2 U3587 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n3113), .Z(n2265) );
  MUX2_X2 U3588 ( .A(n2265), .B(n2264), .S(n3156), .Z(n2266) );
  MUX2_X2 U3589 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n3113), .Z(n2267) );
  MUX2_X2 U3590 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n3113), .Z(n2268) );
  MUX2_X2 U3591 ( .A(n2268), .B(n2267), .S(n3156), .Z(n2269) );
  MUX2_X2 U3592 ( .A(n2269), .B(n2266), .S(n3175), .Z(n2270) );
  MUX2_X2 U3593 ( .A(n2270), .B(n2263), .S(n3187), .Z(n2271) );
  MUX2_X2 U3594 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n3114), .Z(n2272) );
  MUX2_X2 U3595 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n3114), .Z(n2273) );
  MUX2_X2 U3596 ( .A(n2273), .B(n2272), .S(n3157), .Z(n2274) );
  MUX2_X2 U3597 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n3114), .Z(n2275) );
  MUX2_X2 U3598 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n3114), .Z(n2276) );
  MUX2_X2 U3599 ( .A(n2276), .B(n2275), .S(n3157), .Z(n2277) );
  MUX2_X2 U3600 ( .A(n2277), .B(n2274), .S(n3176), .Z(n2278) );
  MUX2_X2 U3601 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n3114), .Z(n2279) );
  MUX2_X2 U3602 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n3114), .Z(n2280) );
  MUX2_X2 U3603 ( .A(n2280), .B(n2279), .S(n3157), .Z(n2281) );
  MUX2_X2 U3604 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n3114), .Z(n2282) );
  MUX2_X2 U3605 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n3114), .Z(n2283) );
  MUX2_X2 U3606 ( .A(n2283), .B(n2282), .S(n3157), .Z(n2284) );
  MUX2_X2 U3607 ( .A(n2284), .B(n2281), .S(n3176), .Z(n2285) );
  MUX2_X2 U3608 ( .A(n2285), .B(n2278), .S(n3186), .Z(n2286) );
  MUX2_X2 U3609 ( .A(n2286), .B(n2271), .S(N13), .Z(rData[4]) );
  MUX2_X2 U3610 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n3114), .Z(n2287) );
  MUX2_X2 U3611 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n3114), .Z(n2288) );
  MUX2_X2 U3612 ( .A(n2288), .B(n2287), .S(n3157), .Z(n2289) );
  MUX2_X2 U3613 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n3114), .Z(n2290) );
  MUX2_X2 U3614 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n3115), .Z(n2291) );
  MUX2_X2 U3615 ( .A(n2291), .B(n2290), .S(n3157), .Z(n2292) );
  MUX2_X2 U3616 ( .A(n2292), .B(n2289), .S(n3176), .Z(n2293) );
  MUX2_X2 U3617 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n3115), .Z(n2294) );
  MUX2_X2 U3618 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n3115), .Z(n2295) );
  MUX2_X2 U3619 ( .A(n2295), .B(n2294), .S(n3157), .Z(n2296) );
  MUX2_X2 U3620 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n3115), .Z(n2297) );
  MUX2_X2 U3621 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n3115), .Z(n2298) );
  MUX2_X2 U3622 ( .A(n2298), .B(n2297), .S(n3157), .Z(n2299) );
  MUX2_X2 U3623 ( .A(n2299), .B(n2296), .S(n3176), .Z(n2300) );
  MUX2_X2 U3624 ( .A(n2300), .B(n2293), .S(n3186), .Z(n2301) );
  MUX2_X2 U3625 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n3115), .Z(n2302) );
  MUX2_X2 U3626 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n3115), .Z(n2303) );
  MUX2_X2 U3627 ( .A(n2303), .B(n2302), .S(n3157), .Z(n2304) );
  MUX2_X2 U3628 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n3115), .Z(n2305) );
  MUX2_X2 U3629 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n3115), .Z(n2306) );
  MUX2_X2 U3630 ( .A(n2306), .B(n2305), .S(n3157), .Z(n2307) );
  MUX2_X2 U3631 ( .A(n2307), .B(n2304), .S(n3176), .Z(n2308) );
  MUX2_X2 U3632 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n3115), .Z(n2309) );
  MUX2_X2 U3633 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n3115), .Z(n2310) );
  MUX2_X2 U3634 ( .A(n2310), .B(n2309), .S(n3157), .Z(n2311) );
  MUX2_X2 U3635 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n3116), .Z(n2312) );
  MUX2_X2 U3636 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n3116), .Z(n2313) );
  MUX2_X2 U3637 ( .A(n2313), .B(n2312), .S(n3158), .Z(n2314) );
  MUX2_X2 U3638 ( .A(n2314), .B(n2311), .S(n3176), .Z(n2315) );
  MUX2_X2 U3639 ( .A(n2315), .B(n2308), .S(n3186), .Z(n2316) );
  MUX2_X2 U3640 ( .A(n2316), .B(n2301), .S(N13), .Z(rData[5]) );
  MUX2_X2 U3641 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n3116), .Z(n2317) );
  MUX2_X2 U3642 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n3116), .Z(n2318) );
  MUX2_X2 U3643 ( .A(n2318), .B(n2317), .S(n3158), .Z(n2319) );
  MUX2_X2 U3644 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n3116), .Z(n2320) );
  MUX2_X2 U3645 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n3116), .Z(n2321) );
  MUX2_X2 U3646 ( .A(n2321), .B(n2320), .S(n3158), .Z(n2322) );
  MUX2_X2 U3647 ( .A(n2322), .B(n2319), .S(n3176), .Z(n2323) );
  MUX2_X2 U3648 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n3116), .Z(n2324) );
  MUX2_X2 U3649 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n3116), .Z(n2325) );
  MUX2_X2 U3650 ( .A(n2325), .B(n2324), .S(n3158), .Z(n2326) );
  MUX2_X2 U3651 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n3116), .Z(n2327) );
  MUX2_X2 U3652 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n3116), .Z(n2328) );
  MUX2_X2 U3653 ( .A(n2328), .B(n2327), .S(n3158), .Z(n2329) );
  MUX2_X2 U3654 ( .A(n2329), .B(n2326), .S(n3176), .Z(n2330) );
  MUX2_X2 U3655 ( .A(n2330), .B(n2323), .S(n3186), .Z(n2331) );
  MUX2_X2 U3656 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n3116), .Z(n2332) );
  MUX2_X2 U3657 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n3117), .Z(n2333) );
  MUX2_X2 U3658 ( .A(n2333), .B(n2332), .S(n3158), .Z(n2334) );
  MUX2_X2 U3659 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n3117), .Z(n2335) );
  MUX2_X2 U3660 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n3117), .Z(n2336) );
  MUX2_X2 U3661 ( .A(n2336), .B(n2335), .S(n3158), .Z(n2337) );
  MUX2_X2 U3662 ( .A(n2337), .B(n2334), .S(n3176), .Z(n2338) );
  MUX2_X2 U3663 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n3117), .Z(n2339) );
  MUX2_X2 U3664 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n3117), .Z(n2340) );
  MUX2_X2 U3665 ( .A(n2340), .B(n2339), .S(n3158), .Z(n2341) );
  MUX2_X2 U3666 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n3117), .Z(n2342) );
  MUX2_X2 U3667 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n3117), .Z(n2343) );
  MUX2_X2 U3668 ( .A(n2343), .B(n2342), .S(n3158), .Z(n2344) );
  MUX2_X2 U3669 ( .A(n2344), .B(n2341), .S(n3176), .Z(n2345) );
  MUX2_X2 U3670 ( .A(n2345), .B(n2338), .S(n3186), .Z(n2346) );
  MUX2_X2 U3671 ( .A(n2346), .B(n2331), .S(N13), .Z(rData[6]) );
  MUX2_X2 U3672 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n3117), .Z(n2347) );
  MUX2_X2 U3673 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n3117), .Z(n2348) );
  MUX2_X2 U3674 ( .A(n2348), .B(n2347), .S(n3158), .Z(n2349) );
  MUX2_X2 U3675 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n3117), .Z(n2350) );
  MUX2_X2 U3676 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n3117), .Z(n2351) );
  MUX2_X2 U3677 ( .A(n2351), .B(n2350), .S(n3158), .Z(n2352) );
  MUX2_X2 U3678 ( .A(n2352), .B(n2349), .S(n3176), .Z(n2353) );
  MUX2_X2 U3679 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n3118), .Z(n2354) );
  MUX2_X2 U3680 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n3118), .Z(n2355) );
  MUX2_X2 U3681 ( .A(n2355), .B(n2354), .S(n3159), .Z(n2356) );
  MUX2_X2 U3682 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n3118), .Z(n2357) );
  MUX2_X2 U3683 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n3118), .Z(n2358) );
  MUX2_X2 U3684 ( .A(n2358), .B(n2357), .S(n3159), .Z(n2359) );
  MUX2_X2 U3685 ( .A(n2359), .B(n2356), .S(n3177), .Z(n2360) );
  MUX2_X2 U3686 ( .A(n2360), .B(n2353), .S(n3186), .Z(n2361) );
  MUX2_X2 U3687 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n3118), .Z(n2362) );
  MUX2_X2 U3688 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n3118), .Z(n2363) );
  MUX2_X2 U3689 ( .A(n2363), .B(n2362), .S(n3159), .Z(n2364) );
  MUX2_X2 U3690 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n3118), .Z(n2365) );
  MUX2_X2 U3691 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n3118), .Z(n2366) );
  MUX2_X2 U3692 ( .A(n2366), .B(n2365), .S(n3159), .Z(n2367) );
  MUX2_X2 U3693 ( .A(n2367), .B(n2364), .S(n3177), .Z(n2368) );
  MUX2_X2 U3694 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n3118), .Z(n2369) );
  MUX2_X2 U3695 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n3118), .Z(n2370) );
  MUX2_X2 U3696 ( .A(n2370), .B(n2369), .S(n3159), .Z(n2371) );
  MUX2_X2 U3697 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n3118), .Z(n2372) );
  MUX2_X2 U3698 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n3119), .Z(n2373) );
  MUX2_X2 U3699 ( .A(n2373), .B(n2372), .S(n3159), .Z(n2374) );
  MUX2_X2 U3700 ( .A(n2374), .B(n2371), .S(n3177), .Z(n2375) );
  MUX2_X2 U3701 ( .A(n2375), .B(n2368), .S(n3186), .Z(n2376) );
  MUX2_X2 U3702 ( .A(n2376), .B(n2361), .S(N13), .Z(rData[7]) );
  MUX2_X2 U3703 ( .A(\mem[30][8] ), .B(\mem[31][8] ), .S(n3119), .Z(n2377) );
  MUX2_X2 U3704 ( .A(\mem[28][8] ), .B(\mem[29][8] ), .S(n3119), .Z(n2378) );
  MUX2_X2 U3705 ( .A(n2378), .B(n2377), .S(n3159), .Z(n2379) );
  MUX2_X2 U3706 ( .A(\mem[26][8] ), .B(\mem[27][8] ), .S(n3119), .Z(n2380) );
  MUX2_X2 U3707 ( .A(\mem[24][8] ), .B(\mem[25][8] ), .S(n3119), .Z(n2381) );
  MUX2_X2 U3708 ( .A(n2381), .B(n2380), .S(n3159), .Z(n2382) );
  MUX2_X2 U3709 ( .A(n2382), .B(n2379), .S(n3177), .Z(n2383) );
  MUX2_X2 U3710 ( .A(\mem[22][8] ), .B(\mem[23][8] ), .S(n3119), .Z(n2384) );
  MUX2_X2 U3711 ( .A(\mem[20][8] ), .B(\mem[21][8] ), .S(n3119), .Z(n2385) );
  MUX2_X2 U3712 ( .A(n2385), .B(n2384), .S(n3159), .Z(n2386) );
  MUX2_X2 U3713 ( .A(\mem[18][8] ), .B(\mem[19][8] ), .S(n3119), .Z(n2387) );
  MUX2_X2 U3714 ( .A(\mem[16][8] ), .B(\mem[17][8] ), .S(n3119), .Z(n2388) );
  MUX2_X2 U3715 ( .A(n2388), .B(n2387), .S(n3159), .Z(n2389) );
  MUX2_X2 U3716 ( .A(n2389), .B(n2386), .S(n3177), .Z(n2390) );
  MUX2_X2 U3717 ( .A(n2390), .B(n2383), .S(n3186), .Z(n2391) );
  MUX2_X2 U3718 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n3119), .Z(n2392) );
  MUX2_X2 U3719 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n3119), .Z(n2393) );
  MUX2_X2 U3720 ( .A(n2393), .B(n2392), .S(n3159), .Z(n2394) );
  MUX2_X2 U3721 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n3120), .Z(n2395) );
  MUX2_X2 U3722 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(n3120), .Z(n2396) );
  MUX2_X2 U3723 ( .A(n2396), .B(n2395), .S(n3160), .Z(n2397) );
  MUX2_X2 U3724 ( .A(n2397), .B(n2394), .S(n3177), .Z(n2398) );
  MUX2_X2 U3725 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n3120), .Z(n2399) );
  MUX2_X2 U3726 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n3120), .Z(n2400) );
  MUX2_X2 U3727 ( .A(n2400), .B(n2399), .S(n3160), .Z(n2401) );
  MUX2_X2 U3728 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n3120), .Z(n2402) );
  MUX2_X2 U3729 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n3120), .Z(n2403) );
  MUX2_X2 U3730 ( .A(n2403), .B(n2402), .S(n3160), .Z(n2404) );
  MUX2_X2 U3731 ( .A(n2404), .B(n2401), .S(n3177), .Z(n2405) );
  MUX2_X2 U3732 ( .A(n2405), .B(n2398), .S(n3186), .Z(n2406) );
  MUX2_X2 U3733 ( .A(n2406), .B(n2391), .S(N13), .Z(rData[8]) );
  MUX2_X2 U3734 ( .A(\mem[30][9] ), .B(\mem[31][9] ), .S(n3120), .Z(n2407) );
  MUX2_X2 U3735 ( .A(\mem[28][9] ), .B(\mem[29][9] ), .S(n3120), .Z(n2408) );
  MUX2_X2 U3736 ( .A(n2408), .B(n2407), .S(n3160), .Z(n2409) );
  MUX2_X2 U3737 ( .A(\mem[26][9] ), .B(\mem[27][9] ), .S(n3120), .Z(n2410) );
  MUX2_X2 U3738 ( .A(\mem[24][9] ), .B(\mem[25][9] ), .S(n3120), .Z(n2411) );
  MUX2_X2 U3739 ( .A(n2411), .B(n2410), .S(n3160), .Z(n2412) );
  MUX2_X2 U3740 ( .A(n2412), .B(n2409), .S(n3177), .Z(n2413) );
  MUX2_X2 U3741 ( .A(\mem[22][9] ), .B(\mem[23][9] ), .S(n3120), .Z(n2414) );
  MUX2_X2 U3742 ( .A(\mem[20][9] ), .B(\mem[21][9] ), .S(n3121), .Z(n2415) );
  MUX2_X2 U3743 ( .A(n2415), .B(n2414), .S(n3160), .Z(n2416) );
  MUX2_X2 U3744 ( .A(\mem[18][9] ), .B(\mem[19][9] ), .S(n3121), .Z(n2417) );
  MUX2_X2 U3745 ( .A(\mem[16][9] ), .B(\mem[17][9] ), .S(n3121), .Z(n2418) );
  MUX2_X2 U3746 ( .A(n2418), .B(n2417), .S(n3160), .Z(n2419) );
  MUX2_X2 U3747 ( .A(n2419), .B(n2416), .S(n3177), .Z(n2420) );
  MUX2_X2 U3748 ( .A(n2420), .B(n2413), .S(n3186), .Z(n2421) );
  MUX2_X2 U3749 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n3121), .Z(n2422) );
  MUX2_X2 U3750 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n3121), .Z(n2423) );
  MUX2_X2 U3751 ( .A(n2423), .B(n2422), .S(n3160), .Z(n2424) );
  MUX2_X2 U3752 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n3121), .Z(n2425) );
  MUX2_X2 U3753 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n3121), .Z(n2426) );
  MUX2_X2 U3754 ( .A(n2426), .B(n2425), .S(n3160), .Z(n2427) );
  MUX2_X2 U3755 ( .A(n2427), .B(n2424), .S(n3177), .Z(n2428) );
  MUX2_X2 U3756 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n3121), .Z(n2429) );
  MUX2_X2 U3757 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n3121), .Z(n2430) );
  MUX2_X2 U3758 ( .A(n2430), .B(n2429), .S(n3160), .Z(n2431) );
  MUX2_X2 U3759 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n3121), .Z(n2432) );
  MUX2_X2 U3760 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n3121), .Z(n2433) );
  MUX2_X2 U3761 ( .A(n2433), .B(n2432), .S(n3160), .Z(n2434) );
  MUX2_X2 U3762 ( .A(n2434), .B(n2431), .S(n3177), .Z(n2435) );
  MUX2_X2 U3763 ( .A(n2435), .B(n2428), .S(n3186), .Z(n2436) );
  MUX2_X2 U3764 ( .A(n2436), .B(n2421), .S(N13), .Z(rData[9]) );
  MUX2_X2 U3765 ( .A(\mem[30][10] ), .B(\mem[31][10] ), .S(n3122), .Z(n2437)
         );
  MUX2_X2 U3766 ( .A(\mem[28][10] ), .B(\mem[29][10] ), .S(n3122), .Z(n2438)
         );
  MUX2_X2 U3767 ( .A(n2438), .B(n2437), .S(n3161), .Z(n2439) );
  MUX2_X2 U3768 ( .A(\mem[26][10] ), .B(\mem[27][10] ), .S(n3122), .Z(n2440)
         );
  MUX2_X2 U3769 ( .A(\mem[24][10] ), .B(\mem[25][10] ), .S(n3122), .Z(n2441)
         );
  MUX2_X2 U3770 ( .A(n2441), .B(n2440), .S(n3161), .Z(n2442) );
  MUX2_X2 U3771 ( .A(n2442), .B(n2439), .S(n3177), .Z(n2443) );
  MUX2_X2 U3772 ( .A(\mem[22][10] ), .B(\mem[23][10] ), .S(n3122), .Z(n2444)
         );
  MUX2_X2 U3773 ( .A(\mem[20][10] ), .B(\mem[21][10] ), .S(n3122), .Z(n2445)
         );
  MUX2_X2 U3774 ( .A(n2445), .B(n2444), .S(n3161), .Z(n2446) );
  MUX2_X2 U3775 ( .A(\mem[18][10] ), .B(\mem[19][10] ), .S(n3122), .Z(n2447)
         );
  MUX2_X2 U3776 ( .A(\mem[16][10] ), .B(\mem[17][10] ), .S(n3122), .Z(n2448)
         );
  MUX2_X2 U3777 ( .A(n2448), .B(n2447), .S(n3161), .Z(n2449) );
  MUX2_X2 U3778 ( .A(n2449), .B(n2446), .S(n3177), .Z(n2450) );
  MUX2_X2 U3779 ( .A(n2450), .B(n2443), .S(n3187), .Z(n2451) );
  MUX2_X2 U3780 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(n3122), .Z(n2452)
         );
  MUX2_X2 U3781 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(n3122), .Z(n2453)
         );
  MUX2_X2 U3782 ( .A(n2453), .B(n2452), .S(n3161), .Z(n2454) );
  MUX2_X2 U3783 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(n3122), .Z(n2455)
         );
  MUX2_X2 U3784 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(n3123), .Z(n2456) );
  MUX2_X2 U3785 ( .A(n2456), .B(n2455), .S(n3161), .Z(n2457) );
  MUX2_X2 U3786 ( .A(n2457), .B(n2454), .S(n3177), .Z(n2458) );
  MUX2_X2 U3787 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n3123), .Z(n2459) );
  MUX2_X2 U3788 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n3123), .Z(n2460) );
  MUX2_X2 U3789 ( .A(n2460), .B(n2459), .S(n3161), .Z(n2461) );
  MUX2_X2 U3790 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n3123), .Z(n2462) );
  MUX2_X2 U3791 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n3123), .Z(n2463) );
  MUX2_X2 U3792 ( .A(n2463), .B(n2462), .S(n3161), .Z(n2464) );
  MUX2_X2 U3793 ( .A(n2464), .B(n2461), .S(n3177), .Z(n2465) );
  MUX2_X2 U3794 ( .A(n2465), .B(n2458), .S(n3187), .Z(n2466) );
  MUX2_X2 U3795 ( .A(n2466), .B(n2451), .S(N13), .Z(rData[10]) );
  MUX2_X2 U3796 ( .A(\mem[30][11] ), .B(\mem[31][11] ), .S(n3123), .Z(n2467)
         );
  MUX2_X2 U3797 ( .A(\mem[28][11] ), .B(\mem[29][11] ), .S(n3123), .Z(n2468)
         );
  MUX2_X2 U3798 ( .A(n2468), .B(n2467), .S(n3161), .Z(n2469) );
  MUX2_X2 U3799 ( .A(\mem[26][11] ), .B(\mem[27][11] ), .S(n3123), .Z(n2470)
         );
  MUX2_X2 U3800 ( .A(\mem[24][11] ), .B(\mem[25][11] ), .S(n3123), .Z(n2471)
         );
  MUX2_X2 U3801 ( .A(n2471), .B(n2470), .S(n3161), .Z(n2472) );
  MUX2_X2 U3802 ( .A(n2472), .B(n2469), .S(n3177), .Z(n2473) );
  MUX2_X2 U3803 ( .A(\mem[22][11] ), .B(\mem[23][11] ), .S(n3123), .Z(n2474)
         );
  MUX2_X2 U3804 ( .A(\mem[20][11] ), .B(\mem[21][11] ), .S(n3123), .Z(n2475)
         );
  MUX2_X2 U3805 ( .A(n2475), .B(n2474), .S(n3161), .Z(n2476) );
  MUX2_X2 U3806 ( .A(\mem[18][11] ), .B(\mem[19][11] ), .S(n3124), .Z(n2477)
         );
  MUX2_X2 U3807 ( .A(\mem[16][11] ), .B(\mem[17][11] ), .S(n3124), .Z(n2478)
         );
  MUX2_X2 U3808 ( .A(n2478), .B(n2477), .S(n3162), .Z(n2479) );
  MUX2_X2 U3809 ( .A(n2479), .B(n2476), .S(n3177), .Z(n2480) );
  MUX2_X2 U3810 ( .A(n2480), .B(n2473), .S(n3187), .Z(n2481) );
  MUX2_X2 U3811 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n3124), .Z(n2482)
         );
  MUX2_X2 U3812 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n3124), .Z(n2483)
         );
  MUX2_X2 U3813 ( .A(n2483), .B(n2482), .S(n3162), .Z(n2484) );
  MUX2_X2 U3814 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n3124), .Z(n2485)
         );
  MUX2_X2 U3815 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(n3124), .Z(n2486) );
  MUX2_X2 U3816 ( .A(n2486), .B(n2485), .S(n3162), .Z(n2487) );
  MUX2_X2 U3817 ( .A(n2487), .B(n2484), .S(n3177), .Z(n2488) );
  MUX2_X2 U3818 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n3124), .Z(n2489) );
  MUX2_X2 U3819 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n3124), .Z(n2490) );
  MUX2_X2 U3820 ( .A(n2490), .B(n2489), .S(n3162), .Z(n2491) );
  MUX2_X2 U3821 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n3124), .Z(n2492) );
  MUX2_X2 U3822 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n3124), .Z(n2493) );
  MUX2_X2 U3823 ( .A(n2493), .B(n2492), .S(n3162), .Z(n2494) );
  MUX2_X2 U3824 ( .A(n2494), .B(n2491), .S(n3177), .Z(n2495) );
  MUX2_X2 U3825 ( .A(n2495), .B(n2488), .S(n3187), .Z(n2496) );
  MUX2_X2 U3826 ( .A(n2496), .B(n2481), .S(N13), .Z(rData[11]) );
  MUX2_X2 U3827 ( .A(\mem[30][12] ), .B(\mem[31][12] ), .S(n3124), .Z(n2497)
         );
  MUX2_X2 U3828 ( .A(\mem[28][12] ), .B(\mem[29][12] ), .S(n3125), .Z(n2498)
         );
  MUX2_X2 U3829 ( .A(n2498), .B(n2497), .S(n3162), .Z(n2499) );
  MUX2_X2 U3830 ( .A(\mem[26][12] ), .B(\mem[27][12] ), .S(n3125), .Z(n2500)
         );
  MUX2_X2 U3831 ( .A(\mem[24][12] ), .B(\mem[25][12] ), .S(n3125), .Z(n2501)
         );
  MUX2_X2 U3832 ( .A(n2501), .B(n2500), .S(n3162), .Z(n2502) );
  MUX2_X2 U3833 ( .A(n2502), .B(n2499), .S(n3177), .Z(n2503) );
  MUX2_X2 U3834 ( .A(\mem[22][12] ), .B(\mem[23][12] ), .S(n3125), .Z(n2504)
         );
  MUX2_X2 U3835 ( .A(\mem[20][12] ), .B(\mem[21][12] ), .S(n3125), .Z(n2505)
         );
  MUX2_X2 U3836 ( .A(n2505), .B(n2504), .S(n3162), .Z(n2506) );
  MUX2_X2 U3837 ( .A(\mem[18][12] ), .B(\mem[19][12] ), .S(n3125), .Z(n2507)
         );
  MUX2_X2 U3838 ( .A(\mem[16][12] ), .B(\mem[17][12] ), .S(n3125), .Z(n2508)
         );
  MUX2_X2 U3839 ( .A(n2508), .B(n2507), .S(n3162), .Z(n2509) );
  MUX2_X2 U3840 ( .A(n2509), .B(n2506), .S(n3177), .Z(n2510) );
  MUX2_X2 U3841 ( .A(n2510), .B(n2503), .S(n3187), .Z(n2511) );
  MUX2_X2 U3842 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n3125), .Z(n2512)
         );
  MUX2_X2 U3843 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n3125), .Z(n2513)
         );
  MUX2_X2 U3844 ( .A(n2513), .B(n2512), .S(n3162), .Z(n2514) );
  MUX2_X2 U3845 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n3125), .Z(n2515)
         );
  MUX2_X2 U3846 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n3125), .Z(n2516) );
  MUX2_X2 U3847 ( .A(n2516), .B(n2515), .S(n3162), .Z(n2517) );
  MUX2_X2 U3848 ( .A(n2517), .B(n2514), .S(n3177), .Z(n2518) );
  MUX2_X2 U3849 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n3126), .Z(n2519) );
  MUX2_X2 U3850 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n3126), .Z(n2520) );
  MUX2_X2 U3851 ( .A(n2520), .B(n2519), .S(n3163), .Z(n2521) );
  MUX2_X2 U3852 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n3126), .Z(n2522) );
  MUX2_X2 U3853 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n3126), .Z(n2523) );
  MUX2_X2 U3854 ( .A(n2523), .B(n2522), .S(n3163), .Z(n2524) );
  MUX2_X2 U3855 ( .A(n2524), .B(n2521), .S(n3178), .Z(n2525) );
  MUX2_X2 U3856 ( .A(n2525), .B(n2518), .S(n3187), .Z(n2526) );
  MUX2_X2 U3857 ( .A(n2526), .B(n2511), .S(N13), .Z(rData[12]) );
  MUX2_X2 U3858 ( .A(\mem[30][13] ), .B(\mem[31][13] ), .S(n3126), .Z(n2527)
         );
  MUX2_X2 U3859 ( .A(\mem[28][13] ), .B(\mem[29][13] ), .S(n3126), .Z(n2528)
         );
  MUX2_X2 U3860 ( .A(n2528), .B(n2527), .S(n3163), .Z(n2529) );
  MUX2_X2 U3861 ( .A(\mem[26][13] ), .B(\mem[27][13] ), .S(n3126), .Z(n2530)
         );
  MUX2_X2 U3862 ( .A(\mem[24][13] ), .B(\mem[25][13] ), .S(n3126), .Z(n2531)
         );
  MUX2_X2 U3863 ( .A(n2531), .B(n2530), .S(n3163), .Z(n2532) );
  MUX2_X2 U3864 ( .A(n2532), .B(n2529), .S(n3178), .Z(n2533) );
  MUX2_X2 U3865 ( .A(\mem[22][13] ), .B(\mem[23][13] ), .S(n3126), .Z(n2534)
         );
  MUX2_X2 U3866 ( .A(\mem[20][13] ), .B(\mem[21][13] ), .S(n3126), .Z(n2535)
         );
  MUX2_X2 U3867 ( .A(n2535), .B(n2534), .S(n3163), .Z(n2536) );
  MUX2_X2 U3868 ( .A(\mem[18][13] ), .B(\mem[19][13] ), .S(n3126), .Z(n2537)
         );
  MUX2_X2 U3869 ( .A(\mem[16][13] ), .B(\mem[17][13] ), .S(n3127), .Z(n2538)
         );
  MUX2_X2 U3870 ( .A(n2538), .B(n2537), .S(n3163), .Z(n2539) );
  MUX2_X2 U3871 ( .A(n2539), .B(n2536), .S(n3178), .Z(n2540) );
  MUX2_X2 U3872 ( .A(n2540), .B(n2533), .S(n3187), .Z(n2541) );
  MUX2_X2 U3873 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n3127), .Z(n2542)
         );
  MUX2_X2 U3874 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(n3127), .Z(n2543)
         );
  MUX2_X2 U3875 ( .A(n2543), .B(n2542), .S(n3163), .Z(n2544) );
  MUX2_X2 U3876 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(n3127), .Z(n2545)
         );
  MUX2_X2 U3877 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(n3127), .Z(n2546) );
  MUX2_X2 U3878 ( .A(n2546), .B(n2545), .S(n3163), .Z(n2547) );
  MUX2_X2 U3879 ( .A(n2547), .B(n2544), .S(n3178), .Z(n2548) );
  MUX2_X2 U3880 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n3127), .Z(n2549) );
  MUX2_X2 U3881 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n3127), .Z(n2550) );
  MUX2_X2 U3882 ( .A(n2550), .B(n2549), .S(n3163), .Z(n2551) );
  MUX2_X2 U3883 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n3127), .Z(n2552) );
  MUX2_X2 U3884 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n3127), .Z(n2553) );
  MUX2_X2 U3885 ( .A(n2553), .B(n2552), .S(n3163), .Z(n2554) );
  MUX2_X2 U3886 ( .A(n2554), .B(n2551), .S(n3178), .Z(n2555) );
  MUX2_X2 U3887 ( .A(n2555), .B(n2548), .S(n3187), .Z(n2556) );
  MUX2_X2 U3888 ( .A(n2556), .B(n2541), .S(N13), .Z(rData[13]) );
  MUX2_X2 U3889 ( .A(\mem[30][14] ), .B(\mem[31][14] ), .S(n3127), .Z(n2557)
         );
  MUX2_X2 U3890 ( .A(\mem[28][14] ), .B(\mem[29][14] ), .S(n3127), .Z(n2558)
         );
  MUX2_X2 U3891 ( .A(n2558), .B(n2557), .S(n3163), .Z(n2559) );
  MUX2_X2 U3892 ( .A(\mem[26][14] ), .B(\mem[27][14] ), .S(n3128), .Z(n2560)
         );
  MUX2_X2 U3893 ( .A(\mem[24][14] ), .B(\mem[25][14] ), .S(n3128), .Z(n2561)
         );
  MUX2_X2 U3894 ( .A(n2561), .B(n2560), .S(n3164), .Z(n2562) );
  MUX2_X2 U3895 ( .A(n2562), .B(n2559), .S(n3178), .Z(n2563) );
  MUX2_X2 U3896 ( .A(\mem[22][14] ), .B(\mem[23][14] ), .S(n3128), .Z(n2564)
         );
  MUX2_X2 U3897 ( .A(\mem[20][14] ), .B(\mem[21][14] ), .S(n3128), .Z(n2565)
         );
  MUX2_X2 U3898 ( .A(n2565), .B(n2564), .S(n3164), .Z(n2566) );
  MUX2_X2 U3899 ( .A(\mem[18][14] ), .B(\mem[19][14] ), .S(n3128), .Z(n2567)
         );
  MUX2_X2 U3900 ( .A(\mem[16][14] ), .B(\mem[17][14] ), .S(n3128), .Z(n2568)
         );
  MUX2_X2 U3901 ( .A(n2568), .B(n2567), .S(n3164), .Z(n2569) );
  MUX2_X2 U3902 ( .A(n2569), .B(n2566), .S(n3178), .Z(n2570) );
  MUX2_X2 U3903 ( .A(n2570), .B(n2563), .S(n3187), .Z(n2571) );
  MUX2_X2 U3904 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n3128), .Z(n2572)
         );
  MUX2_X2 U3905 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n3128), .Z(n2573)
         );
  MUX2_X2 U3906 ( .A(n2573), .B(n2572), .S(n3164), .Z(n2574) );
  MUX2_X2 U3907 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n3128), .Z(n2575)
         );
  MUX2_X2 U3908 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n3128), .Z(n2576) );
  MUX2_X2 U3909 ( .A(n2576), .B(n2575), .S(n3164), .Z(n2577) );
  MUX2_X2 U3910 ( .A(n2577), .B(n2574), .S(n3178), .Z(n2578) );
  MUX2_X2 U3911 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n3128), .Z(n2579) );
  MUX2_X2 U3912 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n3129), .Z(n2580) );
  MUX2_X2 U3913 ( .A(n2580), .B(n2579), .S(n3164), .Z(n2581) );
  MUX2_X2 U3914 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n3129), .Z(n2582) );
  MUX2_X2 U3915 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n3129), .Z(n2583) );
  MUX2_X2 U3916 ( .A(n2583), .B(n2582), .S(n3164), .Z(n2584) );
  MUX2_X2 U3917 ( .A(n2584), .B(n2581), .S(n3178), .Z(n2585) );
  MUX2_X2 U3918 ( .A(n2585), .B(n2578), .S(n3187), .Z(n2586) );
  MUX2_X2 U3919 ( .A(n2586), .B(n2571), .S(N13), .Z(rData[14]) );
  MUX2_X2 U3920 ( .A(\mem[30][15] ), .B(\mem[31][15] ), .S(n3129), .Z(n2587)
         );
  MUX2_X2 U3921 ( .A(\mem[28][15] ), .B(\mem[29][15] ), .S(n3129), .Z(n2588)
         );
  MUX2_X2 U3922 ( .A(n2588), .B(n2587), .S(n3164), .Z(n2589) );
  MUX2_X2 U3923 ( .A(\mem[26][15] ), .B(\mem[27][15] ), .S(n3129), .Z(n2590)
         );
  MUX2_X2 U3924 ( .A(\mem[24][15] ), .B(\mem[25][15] ), .S(n3129), .Z(n2591)
         );
  MUX2_X2 U3925 ( .A(n2591), .B(n2590), .S(n3164), .Z(n2592) );
  MUX2_X2 U3926 ( .A(n2592), .B(n2589), .S(n3178), .Z(n2593) );
  MUX2_X2 U3927 ( .A(\mem[22][15] ), .B(\mem[23][15] ), .S(n3129), .Z(n2594)
         );
  MUX2_X2 U3928 ( .A(\mem[20][15] ), .B(\mem[21][15] ), .S(n3129), .Z(n2595)
         );
  MUX2_X2 U3929 ( .A(n2595), .B(n2594), .S(n3164), .Z(n2596) );
  MUX2_X2 U3930 ( .A(\mem[18][15] ), .B(\mem[19][15] ), .S(n3129), .Z(n2597)
         );
  MUX2_X2 U3931 ( .A(\mem[16][15] ), .B(\mem[17][15] ), .S(n3129), .Z(n2598)
         );
  MUX2_X2 U3932 ( .A(n2598), .B(n2597), .S(n3164), .Z(n2599) );
  MUX2_X2 U3933 ( .A(n2599), .B(n2596), .S(n3178), .Z(n2600) );
  MUX2_X2 U3934 ( .A(n2600), .B(n2593), .S(n3187), .Z(n2601) );
  MUX2_X2 U3935 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n3130), .Z(n2602)
         );
  MUX2_X2 U3936 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n3130), .Z(n2603)
         );
  MUX2_X2 U3937 ( .A(n2603), .B(n2602), .S(n3165), .Z(n2604) );
  MUX2_X2 U3938 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n3130), .Z(n2605)
         );
  MUX2_X2 U3939 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n3130), .Z(n2606) );
  MUX2_X2 U3940 ( .A(n2606), .B(n2605), .S(n3165), .Z(n2607) );
  MUX2_X2 U3941 ( .A(n2607), .B(n2604), .S(n3179), .Z(n2608) );
  MUX2_X2 U3942 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n3130), .Z(n2609) );
  MUX2_X2 U3943 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n3130), .Z(n2610) );
  MUX2_X2 U3944 ( .A(n2610), .B(n2609), .S(n3165), .Z(n2611) );
  MUX2_X2 U3945 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n3130), .Z(n2612) );
  MUX2_X2 U3946 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n3130), .Z(n2613) );
  MUX2_X2 U3947 ( .A(n2613), .B(n2612), .S(n3165), .Z(n2614) );
  MUX2_X2 U3948 ( .A(n2614), .B(n2611), .S(n3179), .Z(n2615) );
  MUX2_X2 U3949 ( .A(n2615), .B(n2608), .S(n3188), .Z(n2616) );
  MUX2_X2 U3950 ( .A(n2616), .B(n2601), .S(N13), .Z(rData[15]) );
  MUX2_X2 U3951 ( .A(\mem[30][16] ), .B(\mem[31][16] ), .S(n3130), .Z(n2617)
         );
  MUX2_X2 U3952 ( .A(\mem[28][16] ), .B(\mem[29][16] ), .S(n3130), .Z(n2618)
         );
  MUX2_X2 U3953 ( .A(n2618), .B(n2617), .S(n3165), .Z(n2619) );
  MUX2_X2 U3954 ( .A(\mem[26][16] ), .B(\mem[27][16] ), .S(n3130), .Z(n2620)
         );
  MUX2_X2 U3955 ( .A(\mem[24][16] ), .B(\mem[25][16] ), .S(n3131), .Z(n2621)
         );
  MUX2_X2 U3956 ( .A(n2621), .B(n2620), .S(n3165), .Z(n2622) );
  MUX2_X2 U3957 ( .A(n2622), .B(n2619), .S(n3179), .Z(n2623) );
  MUX2_X2 U3958 ( .A(\mem[22][16] ), .B(\mem[23][16] ), .S(n3131), .Z(n2624)
         );
  MUX2_X2 U3959 ( .A(\mem[20][16] ), .B(\mem[21][16] ), .S(n3131), .Z(n2625)
         );
  MUX2_X2 U3960 ( .A(n2625), .B(n2624), .S(n3165), .Z(n2626) );
  MUX2_X2 U3961 ( .A(\mem[18][16] ), .B(\mem[19][16] ), .S(n3131), .Z(n2627)
         );
  MUX2_X2 U3962 ( .A(\mem[16][16] ), .B(\mem[17][16] ), .S(n3131), .Z(n2628)
         );
  MUX2_X2 U3963 ( .A(n2628), .B(n2627), .S(n3165), .Z(n2629) );
  MUX2_X2 U3964 ( .A(n2629), .B(n2626), .S(n3179), .Z(n2630) );
  MUX2_X2 U3965 ( .A(n2630), .B(n2623), .S(n3188), .Z(n2631) );
  MUX2_X2 U3966 ( .A(\mem[14][16] ), .B(\mem[15][16] ), .S(n3131), .Z(n2632)
         );
  MUX2_X2 U3967 ( .A(\mem[12][16] ), .B(\mem[13][16] ), .S(n3131), .Z(n2633)
         );
  MUX2_X2 U3968 ( .A(n2633), .B(n2632), .S(n3165), .Z(n2634) );
  MUX2_X2 U3969 ( .A(\mem[10][16] ), .B(\mem[11][16] ), .S(n3131), .Z(n2635)
         );
  MUX2_X2 U3970 ( .A(\mem[8][16] ), .B(\mem[9][16] ), .S(n3131), .Z(n2636) );
  MUX2_X2 U3971 ( .A(n2636), .B(n2635), .S(n3165), .Z(n2637) );
  MUX2_X2 U3972 ( .A(n2637), .B(n2634), .S(n3179), .Z(n2638) );
  MUX2_X2 U3973 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n3131), .Z(n2639) );
  MUX2_X2 U3974 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n3131), .Z(n2640) );
  MUX2_X2 U3975 ( .A(n2640), .B(n2639), .S(n3165), .Z(n2641) );
  MUX2_X2 U3976 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n3132), .Z(n2642) );
  MUX2_X2 U3977 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n3132), .Z(n2643) );
  MUX2_X2 U3978 ( .A(n2643), .B(n2642), .S(n3166), .Z(n2644) );
  MUX2_X2 U3979 ( .A(n2644), .B(n2641), .S(n3179), .Z(n2645) );
  MUX2_X2 U3980 ( .A(n2645), .B(n2638), .S(n3188), .Z(n2646) );
  MUX2_X2 U3981 ( .A(n2646), .B(n2631), .S(N13), .Z(rData[16]) );
  MUX2_X2 U3982 ( .A(\mem[30][17] ), .B(\mem[31][17] ), .S(n3132), .Z(n2647)
         );
  MUX2_X2 U3983 ( .A(\mem[28][17] ), .B(\mem[29][17] ), .S(n3132), .Z(n2648)
         );
  MUX2_X2 U3984 ( .A(n2648), .B(n2647), .S(n3166), .Z(n2649) );
  MUX2_X2 U3985 ( .A(\mem[26][17] ), .B(\mem[27][17] ), .S(n3132), .Z(n2650)
         );
  MUX2_X2 U3986 ( .A(\mem[24][17] ), .B(\mem[25][17] ), .S(n3132), .Z(n2651)
         );
  MUX2_X2 U3987 ( .A(n2651), .B(n2650), .S(n3166), .Z(n2652) );
  MUX2_X2 U3988 ( .A(n2652), .B(n2649), .S(n3179), .Z(n2653) );
  MUX2_X2 U3989 ( .A(\mem[22][17] ), .B(\mem[23][17] ), .S(n3132), .Z(n2654)
         );
  MUX2_X2 U3990 ( .A(\mem[20][17] ), .B(\mem[21][17] ), .S(n3132), .Z(n2655)
         );
  MUX2_X2 U3991 ( .A(n2655), .B(n2654), .S(n3166), .Z(n2656) );
  MUX2_X2 U3992 ( .A(\mem[18][17] ), .B(\mem[19][17] ), .S(n3132), .Z(n2657)
         );
  MUX2_X2 U3993 ( .A(\mem[16][17] ), .B(\mem[17][17] ), .S(n3132), .Z(n2658)
         );
  MUX2_X2 U3994 ( .A(n2658), .B(n2657), .S(n3166), .Z(n2659) );
  MUX2_X2 U3995 ( .A(n2659), .B(n2656), .S(n3179), .Z(n2660) );
  MUX2_X2 U3996 ( .A(n2660), .B(n2653), .S(n3188), .Z(n2661) );
  MUX2_X2 U3997 ( .A(\mem[14][17] ), .B(\mem[15][17] ), .S(n3132), .Z(n2662)
         );
  MUX2_X2 U3998 ( .A(\mem[12][17] ), .B(\mem[13][17] ), .S(n3133), .Z(n2663)
         );
  MUX2_X2 U3999 ( .A(n2663), .B(n2662), .S(n3166), .Z(n2664) );
  MUX2_X2 U4000 ( .A(\mem[10][17] ), .B(\mem[11][17] ), .S(n3133), .Z(n2665)
         );
  MUX2_X2 U4001 ( .A(\mem[8][17] ), .B(\mem[9][17] ), .S(n3133), .Z(n2666) );
  MUX2_X2 U4002 ( .A(n2666), .B(n2665), .S(n3166), .Z(n2667) );
  MUX2_X2 U4003 ( .A(n2667), .B(n2664), .S(n3179), .Z(n2668) );
  MUX2_X2 U4004 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n3133), .Z(n2669) );
  MUX2_X2 U4005 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n3133), .Z(n2670) );
  MUX2_X2 U4006 ( .A(n2670), .B(n2669), .S(n3166), .Z(n2671) );
  MUX2_X2 U4007 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n3133), .Z(n2672) );
  MUX2_X2 U4008 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n3133), .Z(n2673) );
  MUX2_X2 U4009 ( .A(n2673), .B(n2672), .S(n3166), .Z(n2674) );
  MUX2_X2 U4010 ( .A(n2674), .B(n2671), .S(n3179), .Z(n2675) );
  MUX2_X2 U4011 ( .A(n2675), .B(n2668), .S(n3188), .Z(n2676) );
  MUX2_X2 U4012 ( .A(n2676), .B(n2661), .S(N13), .Z(rData[17]) );
  MUX2_X2 U4013 ( .A(\mem[30][18] ), .B(\mem[31][18] ), .S(n3133), .Z(n2677)
         );
  MUX2_X2 U4014 ( .A(\mem[28][18] ), .B(\mem[29][18] ), .S(n3133), .Z(n2678)
         );
  MUX2_X2 U4015 ( .A(n2678), .B(n2677), .S(n3166), .Z(n2679) );
  MUX2_X2 U4016 ( .A(\mem[26][18] ), .B(\mem[27][18] ), .S(n3133), .Z(n2680)
         );
  MUX2_X2 U4017 ( .A(\mem[24][18] ), .B(\mem[25][18] ), .S(n3133), .Z(n2681)
         );
  MUX2_X2 U4018 ( .A(n2681), .B(n2680), .S(n3166), .Z(n2682) );
  MUX2_X2 U4019 ( .A(n2682), .B(n2679), .S(n3179), .Z(n2683) );
  MUX2_X2 U4020 ( .A(\mem[22][18] ), .B(\mem[23][18] ), .S(n3134), .Z(n2684)
         );
  MUX2_X2 U4021 ( .A(\mem[20][18] ), .B(\mem[21][18] ), .S(n3134), .Z(n2685)
         );
  MUX2_X2 U4022 ( .A(n2685), .B(n2684), .S(n3167), .Z(n2686) );
  MUX2_X2 U4023 ( .A(\mem[18][18] ), .B(\mem[19][18] ), .S(n3134), .Z(n2687)
         );
  MUX2_X2 U4024 ( .A(\mem[16][18] ), .B(\mem[17][18] ), .S(n3134), .Z(n2688)
         );
  MUX2_X2 U4025 ( .A(n2688), .B(n2687), .S(n3167), .Z(n2689) );
  MUX2_X2 U4026 ( .A(n2689), .B(n2686), .S(n3180), .Z(n2690) );
  MUX2_X2 U4027 ( .A(n2690), .B(n2683), .S(n3188), .Z(n2691) );
  MUX2_X2 U4028 ( .A(\mem[14][18] ), .B(\mem[15][18] ), .S(n3134), .Z(n2692)
         );
  MUX2_X2 U4029 ( .A(\mem[12][18] ), .B(\mem[13][18] ), .S(n3134), .Z(n2693)
         );
  MUX2_X2 U4030 ( .A(n2693), .B(n2692), .S(n3167), .Z(n2694) );
  MUX2_X2 U4031 ( .A(\mem[10][18] ), .B(\mem[11][18] ), .S(n3134), .Z(n2695)
         );
  MUX2_X2 U4032 ( .A(\mem[8][18] ), .B(\mem[9][18] ), .S(n3134), .Z(n2696) );
  MUX2_X2 U4033 ( .A(n2696), .B(n2695), .S(n3167), .Z(n2697) );
  MUX2_X2 U4034 ( .A(n2697), .B(n2694), .S(n3180), .Z(n2698) );
  MUX2_X2 U4035 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n3134), .Z(n2699) );
  MUX2_X2 U4036 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n3134), .Z(n2700) );
  MUX2_X2 U4037 ( .A(n2700), .B(n2699), .S(n3167), .Z(n2701) );
  MUX2_X2 U4038 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n3134), .Z(n2702) );
  MUX2_X2 U4039 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n3135), .Z(n2703) );
  MUX2_X2 U4040 ( .A(n2703), .B(n2702), .S(n3167), .Z(n2704) );
  MUX2_X2 U4041 ( .A(n2704), .B(n2701), .S(n3180), .Z(n2705) );
  MUX2_X2 U4042 ( .A(n2705), .B(n2698), .S(n3188), .Z(n2706) );
  MUX2_X2 U4043 ( .A(n2706), .B(n2691), .S(N13), .Z(rData[18]) );
  MUX2_X2 U4044 ( .A(\mem[30][19] ), .B(\mem[31][19] ), .S(n3135), .Z(n2707)
         );
  MUX2_X2 U4045 ( .A(\mem[28][19] ), .B(\mem[29][19] ), .S(n3135), .Z(n2708)
         );
  MUX2_X2 U4046 ( .A(n2708), .B(n2707), .S(n3167), .Z(n2709) );
  MUX2_X2 U4047 ( .A(\mem[26][19] ), .B(\mem[27][19] ), .S(n3135), .Z(n2710)
         );
  MUX2_X2 U4048 ( .A(\mem[24][19] ), .B(\mem[25][19] ), .S(n3135), .Z(n2711)
         );
  MUX2_X2 U4049 ( .A(n2711), .B(n2710), .S(n3167), .Z(n2712) );
  MUX2_X2 U4050 ( .A(n2712), .B(n2709), .S(n3180), .Z(n2713) );
  MUX2_X2 U4051 ( .A(\mem[22][19] ), .B(\mem[23][19] ), .S(n3135), .Z(n2714)
         );
  MUX2_X2 U4052 ( .A(\mem[20][19] ), .B(\mem[21][19] ), .S(n3135), .Z(n2715)
         );
  MUX2_X2 U4053 ( .A(n2715), .B(n2714), .S(n3167), .Z(n2716) );
  MUX2_X2 U4054 ( .A(\mem[18][19] ), .B(\mem[19][19] ), .S(n3135), .Z(n2717)
         );
  MUX2_X2 U4055 ( .A(\mem[16][19] ), .B(\mem[17][19] ), .S(n3135), .Z(n2718)
         );
  MUX2_X2 U4056 ( .A(n2718), .B(n2717), .S(n3167), .Z(n2719) );
  MUX2_X2 U4057 ( .A(n2719), .B(n2716), .S(n3180), .Z(n2720) );
  MUX2_X2 U4058 ( .A(n2720), .B(n2713), .S(n3188), .Z(n2721) );
  MUX2_X2 U4059 ( .A(\mem[14][19] ), .B(\mem[15][19] ), .S(n3135), .Z(n2722)
         );
  MUX2_X2 U4060 ( .A(\mem[12][19] ), .B(\mem[13][19] ), .S(n3135), .Z(n2723)
         );
  MUX2_X2 U4061 ( .A(n2723), .B(n2722), .S(n3167), .Z(n2724) );
  MUX2_X2 U4062 ( .A(\mem[10][19] ), .B(\mem[11][19] ), .S(n3136), .Z(n2725)
         );
  MUX2_X2 U4063 ( .A(\mem[8][19] ), .B(\mem[9][19] ), .S(n3136), .Z(n2726) );
  MUX2_X2 U4064 ( .A(n2726), .B(n2725), .S(n3168), .Z(n2727) );
  MUX2_X2 U4065 ( .A(n2727), .B(n2724), .S(n3180), .Z(n2728) );
  MUX2_X2 U4066 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n3136), .Z(n2729) );
  MUX2_X2 U4067 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n3136), .Z(n2730) );
  MUX2_X2 U4068 ( .A(n2730), .B(n2729), .S(n3168), .Z(n2731) );
  MUX2_X2 U4069 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n3136), .Z(n2732) );
  MUX2_X2 U4070 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n3136), .Z(n2733) );
  MUX2_X2 U4071 ( .A(n2733), .B(n2732), .S(n3168), .Z(n2734) );
  MUX2_X2 U4072 ( .A(n2734), .B(n2731), .S(n3180), .Z(n2735) );
  MUX2_X2 U4073 ( .A(n2735), .B(n2728), .S(n3188), .Z(n2736) );
  MUX2_X2 U4074 ( .A(n2736), .B(n2721), .S(N13), .Z(rData[19]) );
  MUX2_X2 U4075 ( .A(\mem[30][20] ), .B(\mem[31][20] ), .S(n3136), .Z(n2737)
         );
  MUX2_X2 U4076 ( .A(\mem[28][20] ), .B(\mem[29][20] ), .S(n3136), .Z(n2738)
         );
  MUX2_X2 U4077 ( .A(n2738), .B(n2737), .S(n3168), .Z(n2739) );
  MUX2_X2 U4078 ( .A(\mem[26][20] ), .B(\mem[27][20] ), .S(n3136), .Z(n2740)
         );
  MUX2_X2 U4079 ( .A(\mem[24][20] ), .B(\mem[25][20] ), .S(n3136), .Z(n2741)
         );
  MUX2_X2 U4080 ( .A(n2741), .B(n2740), .S(n3168), .Z(n2742) );
  MUX2_X2 U4081 ( .A(n2742), .B(n2739), .S(n3180), .Z(n2743) );
  MUX2_X2 U4082 ( .A(\mem[22][20] ), .B(\mem[23][20] ), .S(n3136), .Z(n2744)
         );
  MUX2_X2 U4083 ( .A(\mem[20][20] ), .B(\mem[21][20] ), .S(n3137), .Z(n2745)
         );
  MUX2_X2 U4084 ( .A(n2745), .B(n2744), .S(n3168), .Z(n2746) );
  MUX2_X2 U4085 ( .A(\mem[18][20] ), .B(\mem[19][20] ), .S(n3137), .Z(n2747)
         );
  MUX2_X2 U4086 ( .A(\mem[16][20] ), .B(\mem[17][20] ), .S(n3137), .Z(n2748)
         );
  MUX2_X2 U4087 ( .A(n2748), .B(n2747), .S(n3168), .Z(n2749) );
  MUX2_X2 U4088 ( .A(n2749), .B(n2746), .S(n3180), .Z(n2750) );
  MUX2_X2 U4089 ( .A(n2750), .B(n2743), .S(n3188), .Z(n2751) );
  MUX2_X2 U4090 ( .A(\mem[14][20] ), .B(\mem[15][20] ), .S(n3137), .Z(n2752)
         );
  MUX2_X2 U4091 ( .A(\mem[12][20] ), .B(\mem[13][20] ), .S(n3137), .Z(n2753)
         );
  MUX2_X2 U4092 ( .A(n2753), .B(n2752), .S(n3168), .Z(n2754) );
  MUX2_X2 U4093 ( .A(\mem[10][20] ), .B(\mem[11][20] ), .S(n3137), .Z(n2755)
         );
  MUX2_X2 U4094 ( .A(\mem[8][20] ), .B(\mem[9][20] ), .S(n3137), .Z(n2756) );
  MUX2_X2 U4095 ( .A(n2756), .B(n2755), .S(n3168), .Z(n2757) );
  MUX2_X2 U4096 ( .A(n2757), .B(n2754), .S(n3180), .Z(n2758) );
  MUX2_X2 U4097 ( .A(\mem[6][20] ), .B(\mem[7][20] ), .S(n3137), .Z(n2759) );
  MUX2_X2 U4098 ( .A(\mem[4][20] ), .B(\mem[5][20] ), .S(n3137), .Z(n2760) );
  MUX2_X2 U4099 ( .A(n2760), .B(n2759), .S(n3168), .Z(n2761) );
  MUX2_X2 U4100 ( .A(\mem[2][20] ), .B(\mem[3][20] ), .S(n3137), .Z(n2762) );
  MUX2_X2 U4101 ( .A(\mem[0][20] ), .B(\mem[1][20] ), .S(n3137), .Z(n2763) );
  MUX2_X2 U4102 ( .A(n2763), .B(n2762), .S(n3168), .Z(n2764) );
  MUX2_X2 U4103 ( .A(n2764), .B(n2761), .S(n3180), .Z(n2765) );
  MUX2_X2 U4104 ( .A(n2765), .B(n2758), .S(n3188), .Z(n2766) );
  MUX2_X2 U4105 ( .A(n2766), .B(n2751), .S(N13), .Z(rData[20]) );
  MUX2_X2 U4106 ( .A(\mem[30][21] ), .B(\mem[31][21] ), .S(n3138), .Z(n2767)
         );
  MUX2_X2 U4107 ( .A(\mem[28][21] ), .B(\mem[29][21] ), .S(n3138), .Z(n2768)
         );
  MUX2_X2 U4108 ( .A(n2768), .B(n2767), .S(n3169), .Z(n2769) );
  MUX2_X2 U4109 ( .A(\mem[26][21] ), .B(\mem[27][21] ), .S(n3138), .Z(n2770)
         );
  MUX2_X2 U4110 ( .A(\mem[24][21] ), .B(\mem[25][21] ), .S(n3138), .Z(n2771)
         );
  MUX2_X2 U4111 ( .A(n2771), .B(n2770), .S(n3169), .Z(n2772) );
  MUX2_X2 U4112 ( .A(n2772), .B(n2769), .S(n3180), .Z(n2773) );
  MUX2_X2 U4113 ( .A(\mem[22][21] ), .B(\mem[23][21] ), .S(n3138), .Z(n2774)
         );
  MUX2_X2 U4114 ( .A(\mem[20][21] ), .B(\mem[21][21] ), .S(n3138), .Z(n2775)
         );
  MUX2_X2 U4115 ( .A(n2775), .B(n2774), .S(n3169), .Z(n2776) );
  MUX2_X2 U4116 ( .A(\mem[18][21] ), .B(\mem[19][21] ), .S(n3138), .Z(n2777)
         );
  MUX2_X2 U4117 ( .A(\mem[16][21] ), .B(\mem[17][21] ), .S(n3138), .Z(n2778)
         );
  MUX2_X2 U4118 ( .A(n2778), .B(n2777), .S(n3169), .Z(n2779) );
  MUX2_X2 U4119 ( .A(n2779), .B(n2776), .S(n3180), .Z(n2780) );
  MUX2_X2 U4120 ( .A(n2780), .B(n2773), .S(n3189), .Z(n2781) );
  MUX2_X2 U4121 ( .A(\mem[14][21] ), .B(\mem[15][21] ), .S(n3138), .Z(n2782)
         );
  MUX2_X2 U4122 ( .A(\mem[12][21] ), .B(\mem[13][21] ), .S(n3138), .Z(n2783)
         );
  MUX2_X2 U4123 ( .A(n2783), .B(n2782), .S(n3169), .Z(n2784) );
  MUX2_X2 U4124 ( .A(\mem[10][21] ), .B(\mem[11][21] ), .S(n3138), .Z(n2785)
         );
  MUX2_X2 U4125 ( .A(\mem[8][21] ), .B(\mem[9][21] ), .S(n3139), .Z(n2786) );
  MUX2_X2 U4126 ( .A(n2786), .B(n2785), .S(n3169), .Z(n2787) );
  MUX2_X2 U4127 ( .A(n2787), .B(n2784), .S(n3179), .Z(n2788) );
  MUX2_X2 U4128 ( .A(\mem[6][21] ), .B(\mem[7][21] ), .S(n3139), .Z(n2789) );
  MUX2_X2 U4129 ( .A(\mem[4][21] ), .B(\mem[5][21] ), .S(n3139), .Z(n2790) );
  MUX2_X2 U4130 ( .A(n2790), .B(n2789), .S(n3169), .Z(n2791) );
  MUX2_X2 U4131 ( .A(\mem[2][21] ), .B(\mem[3][21] ), .S(n3139), .Z(n2792) );
  MUX2_X2 U4132 ( .A(\mem[0][21] ), .B(\mem[1][21] ), .S(n3139), .Z(n2793) );
  MUX2_X2 U4133 ( .A(n2793), .B(n2792), .S(n3169), .Z(n2794) );
  MUX2_X2 U4134 ( .A(n2794), .B(n2791), .S(n3177), .Z(n2795) );
  MUX2_X2 U4135 ( .A(n2795), .B(n2788), .S(n3189), .Z(n2796) );
  MUX2_X2 U4136 ( .A(n2796), .B(n2781), .S(N13), .Z(rData[21]) );
  MUX2_X2 U4137 ( .A(\mem[30][22] ), .B(\mem[31][22] ), .S(n3139), .Z(n2797)
         );
  MUX2_X2 U4138 ( .A(\mem[28][22] ), .B(\mem[29][22] ), .S(n3139), .Z(n2798)
         );
  MUX2_X2 U4139 ( .A(n2798), .B(n2797), .S(n3169), .Z(n2799) );
  MUX2_X2 U4140 ( .A(\mem[26][22] ), .B(\mem[27][22] ), .S(n3139), .Z(n2800)
         );
  MUX2_X2 U4141 ( .A(\mem[24][22] ), .B(\mem[25][22] ), .S(n3139), .Z(n2801)
         );
  MUX2_X2 U4142 ( .A(n2801), .B(n2800), .S(n3169), .Z(n2802) );
  MUX2_X2 U4143 ( .A(n2802), .B(n2799), .S(n3179), .Z(n2803) );
  MUX2_X2 U4144 ( .A(\mem[22][22] ), .B(\mem[23][22] ), .S(n3139), .Z(n2804)
         );
  MUX2_X2 U4145 ( .A(\mem[20][22] ), .B(\mem[21][22] ), .S(n3139), .Z(n2805)
         );
  MUX2_X2 U4146 ( .A(n2805), .B(n2804), .S(n3169), .Z(n2806) );
  MUX2_X2 U4147 ( .A(\mem[18][22] ), .B(\mem[19][22] ), .S(n3140), .Z(n2807)
         );
  MUX2_X2 U4148 ( .A(\mem[16][22] ), .B(\mem[17][22] ), .S(n3140), .Z(n2808)
         );
  MUX2_X2 U4149 ( .A(n2808), .B(n2807), .S(n3170), .Z(n2809) );
  MUX2_X2 U4150 ( .A(n2809), .B(n2806), .S(n3179), .Z(n2810) );
  MUX2_X2 U4151 ( .A(n2810), .B(n2803), .S(n3189), .Z(n2811) );
  MUX2_X2 U4152 ( .A(\mem[14][22] ), .B(\mem[15][22] ), .S(n3140), .Z(n2812)
         );
  MUX2_X2 U4153 ( .A(\mem[12][22] ), .B(\mem[13][22] ), .S(n3140), .Z(n2813)
         );
  MUX2_X2 U4154 ( .A(n2813), .B(n2812), .S(n3170), .Z(n2814) );
  MUX2_X2 U4155 ( .A(\mem[10][22] ), .B(\mem[11][22] ), .S(n3140), .Z(n2815)
         );
  MUX2_X2 U4156 ( .A(\mem[8][22] ), .B(\mem[9][22] ), .S(n3140), .Z(n2816) );
  MUX2_X2 U4157 ( .A(n2816), .B(n2815), .S(n3170), .Z(n2817) );
  MUX2_X2 U4158 ( .A(n2817), .B(n2814), .S(n3180), .Z(n2818) );
  MUX2_X2 U4159 ( .A(\mem[6][22] ), .B(\mem[7][22] ), .S(n3140), .Z(n2819) );
  MUX2_X2 U4160 ( .A(\mem[4][22] ), .B(\mem[5][22] ), .S(n3140), .Z(n2820) );
  MUX2_X2 U4161 ( .A(n2820), .B(n2819), .S(n3170), .Z(n2821) );
  MUX2_X2 U4162 ( .A(\mem[2][22] ), .B(\mem[3][22] ), .S(n3140), .Z(n2822) );
  MUX2_X2 U4163 ( .A(\mem[0][22] ), .B(\mem[1][22] ), .S(n3140), .Z(n2823) );
  MUX2_X2 U4164 ( .A(n2823), .B(n2822), .S(n3170), .Z(n2824) );
  MUX2_X2 U4165 ( .A(n2824), .B(n2821), .S(n3177), .Z(n2825) );
  MUX2_X2 U4166 ( .A(n2825), .B(n2818), .S(n3189), .Z(n2826) );
  MUX2_X2 U4167 ( .A(n2826), .B(n2811), .S(N13), .Z(rData[22]) );
  MUX2_X2 U4168 ( .A(\mem[30][23] ), .B(\mem[31][23] ), .S(n3140), .Z(n2827)
         );
  MUX2_X2 U4169 ( .A(\mem[28][23] ), .B(\mem[29][23] ), .S(n3141), .Z(n2828)
         );
  MUX2_X2 U4170 ( .A(n2828), .B(n2827), .S(n3170), .Z(n2829) );
  MUX2_X2 U4171 ( .A(\mem[26][23] ), .B(\mem[27][23] ), .S(n3141), .Z(n2830)
         );
  MUX2_X2 U4172 ( .A(\mem[24][23] ), .B(\mem[25][23] ), .S(n3141), .Z(n2831)
         );
  MUX2_X2 U4173 ( .A(n2831), .B(n2830), .S(n3170), .Z(n2832) );
  MUX2_X2 U4174 ( .A(n2832), .B(n2829), .S(n3180), .Z(n2833) );
  MUX2_X2 U4175 ( .A(\mem[22][23] ), .B(\mem[23][23] ), .S(n3141), .Z(n2834)
         );
  MUX2_X2 U4176 ( .A(\mem[20][23] ), .B(\mem[21][23] ), .S(n3141), .Z(n2835)
         );
  MUX2_X2 U4177 ( .A(n2835), .B(n2834), .S(n3170), .Z(n2836) );
  MUX2_X2 U4178 ( .A(\mem[18][23] ), .B(\mem[19][23] ), .S(n3141), .Z(n2837)
         );
  MUX2_X2 U4179 ( .A(\mem[16][23] ), .B(\mem[17][23] ), .S(n3141), .Z(n2838)
         );
  MUX2_X2 U4180 ( .A(n2838), .B(n2837), .S(n3170), .Z(n2839) );
  MUX2_X2 U4181 ( .A(n2839), .B(n2836), .S(n3178), .Z(n2840) );
  MUX2_X2 U4182 ( .A(n2840), .B(n2833), .S(n3189), .Z(n2841) );
  MUX2_X2 U4183 ( .A(\mem[14][23] ), .B(\mem[15][23] ), .S(n3141), .Z(n2842)
         );
  MUX2_X2 U4184 ( .A(\mem[12][23] ), .B(\mem[13][23] ), .S(n3141), .Z(n2843)
         );
  MUX2_X2 U4185 ( .A(n2843), .B(n2842), .S(n3170), .Z(n2844) );
  MUX2_X2 U4186 ( .A(\mem[10][23] ), .B(\mem[11][23] ), .S(n3141), .Z(n2845)
         );
  MUX2_X2 U4187 ( .A(\mem[8][23] ), .B(\mem[9][23] ), .S(n3141), .Z(n2846) );
  MUX2_X2 U4188 ( .A(n2846), .B(n2845), .S(n3170), .Z(n2847) );
  MUX2_X2 U4189 ( .A(n2847), .B(n2844), .S(n3179), .Z(n2848) );
  MUX2_X2 U4190 ( .A(\mem[6][23] ), .B(\mem[7][23] ), .S(n3142), .Z(n2849) );
  MUX2_X2 U4191 ( .A(\mem[4][23] ), .B(\mem[5][23] ), .S(n3142), .Z(n2850) );
  MUX2_X2 U4192 ( .A(n2850), .B(n2849), .S(n3171), .Z(n2851) );
  MUX2_X2 U4193 ( .A(\mem[2][23] ), .B(\mem[3][23] ), .S(n3142), .Z(n2852) );
  MUX2_X2 U4194 ( .A(\mem[0][23] ), .B(\mem[1][23] ), .S(n3142), .Z(n2853) );
  MUX2_X2 U4195 ( .A(n2853), .B(n2852), .S(n3171), .Z(n2854) );
  MUX2_X2 U4196 ( .A(n2854), .B(n2851), .S(n3181), .Z(n2855) );
  MUX2_X2 U4197 ( .A(n2855), .B(n2848), .S(n3189), .Z(n2856) );
  MUX2_X2 U4198 ( .A(n2856), .B(n2841), .S(N13), .Z(rData[23]) );
  MUX2_X2 U4199 ( .A(\mem[30][24] ), .B(\mem[31][24] ), .S(n3142), .Z(n2857)
         );
  MUX2_X2 U4200 ( .A(\mem[28][24] ), .B(\mem[29][24] ), .S(n3142), .Z(n2858)
         );
  MUX2_X2 U4201 ( .A(n2858), .B(n2857), .S(n3171), .Z(n2859) );
  MUX2_X2 U4202 ( .A(\mem[26][24] ), .B(\mem[27][24] ), .S(n3142), .Z(n2860)
         );
  MUX2_X2 U4203 ( .A(\mem[24][24] ), .B(\mem[25][24] ), .S(n3142), .Z(n2861)
         );
  MUX2_X2 U4204 ( .A(n2861), .B(n2860), .S(n3171), .Z(n2862) );
  MUX2_X2 U4205 ( .A(n2862), .B(n2859), .S(n3181), .Z(n2863) );
  MUX2_X2 U4206 ( .A(\mem[22][24] ), .B(\mem[23][24] ), .S(n3142), .Z(n2864)
         );
  MUX2_X2 U4207 ( .A(\mem[20][24] ), .B(\mem[21][24] ), .S(n3142), .Z(n2865)
         );
  MUX2_X2 U4208 ( .A(n2865), .B(n2864), .S(n3171), .Z(n2866) );
  MUX2_X2 U4209 ( .A(\mem[18][24] ), .B(\mem[19][24] ), .S(n3142), .Z(n2867)
         );
  MUX2_X2 U4210 ( .A(\mem[16][24] ), .B(\mem[17][24] ), .S(n3143), .Z(n2868)
         );
  MUX2_X2 U4211 ( .A(n2868), .B(n2867), .S(n3171), .Z(n2869) );
  MUX2_X2 U4212 ( .A(n2869), .B(n2866), .S(n3181), .Z(n2870) );
  MUX2_X2 U4213 ( .A(n2870), .B(n2863), .S(n3189), .Z(n2871) );
  MUX2_X2 U4214 ( .A(\mem[14][24] ), .B(\mem[15][24] ), .S(n3143), .Z(n2872)
         );
  MUX2_X2 U4215 ( .A(\mem[12][24] ), .B(\mem[13][24] ), .S(n3143), .Z(n2873)
         );
  MUX2_X2 U4216 ( .A(n2873), .B(n2872), .S(n3171), .Z(n2874) );
  MUX2_X2 U4217 ( .A(\mem[10][24] ), .B(\mem[11][24] ), .S(n3143), .Z(n2875)
         );
  MUX2_X2 U4218 ( .A(\mem[8][24] ), .B(\mem[9][24] ), .S(n3143), .Z(n2876) );
  MUX2_X2 U4219 ( .A(n2876), .B(n2875), .S(n3171), .Z(n2877) );
  MUX2_X2 U4220 ( .A(n2877), .B(n2874), .S(n3181), .Z(n2878) );
  MUX2_X2 U4221 ( .A(\mem[6][24] ), .B(\mem[7][24] ), .S(n3143), .Z(n2879) );
  MUX2_X2 U4222 ( .A(\mem[4][24] ), .B(\mem[5][24] ), .S(n3143), .Z(n2880) );
  MUX2_X2 U4223 ( .A(n2880), .B(n2879), .S(n3171), .Z(n2881) );
  MUX2_X2 U4224 ( .A(\mem[2][24] ), .B(\mem[3][24] ), .S(n3143), .Z(n2882) );
  MUX2_X2 U4225 ( .A(\mem[0][24] ), .B(\mem[1][24] ), .S(n3143), .Z(n2883) );
  MUX2_X2 U4226 ( .A(n2883), .B(n2882), .S(n3171), .Z(n2884) );
  MUX2_X2 U4227 ( .A(n2884), .B(n2881), .S(n3181), .Z(n2885) );
  MUX2_X2 U4228 ( .A(n2885), .B(n2878), .S(n3189), .Z(n2886) );
  MUX2_X2 U4229 ( .A(n2886), .B(n2871), .S(N13), .Z(rData[24]) );
  MUX2_X2 U4230 ( .A(\mem[30][25] ), .B(\mem[31][25] ), .S(n3143), .Z(n2887)
         );
  MUX2_X2 U4231 ( .A(\mem[28][25] ), .B(\mem[29][25] ), .S(n3143), .Z(n2888)
         );
  MUX2_X2 U4232 ( .A(n2888), .B(n2887), .S(n3171), .Z(n2889) );
  MUX2_X2 U4233 ( .A(\mem[26][25] ), .B(\mem[27][25] ), .S(n3144), .Z(n2890)
         );
  MUX2_X2 U4234 ( .A(\mem[24][25] ), .B(\mem[25][25] ), .S(n3144), .Z(n2891)
         );
  MUX2_X2 U4235 ( .A(n2891), .B(n2890), .S(N10), .Z(n2892) );
  MUX2_X2 U4236 ( .A(n2892), .B(n2889), .S(n3181), .Z(n2893) );
  MUX2_X2 U4237 ( .A(\mem[22][25] ), .B(\mem[23][25] ), .S(n3144), .Z(n2894)
         );
  MUX2_X2 U4238 ( .A(\mem[20][25] ), .B(\mem[21][25] ), .S(n3144), .Z(n2895)
         );
  MUX2_X2 U4239 ( .A(n2895), .B(n2894), .S(N10), .Z(n2896) );
  MUX2_X2 U4240 ( .A(\mem[18][25] ), .B(\mem[19][25] ), .S(n3144), .Z(n2897)
         );
  MUX2_X2 U4241 ( .A(\mem[16][25] ), .B(\mem[17][25] ), .S(n3144), .Z(n2898)
         );
  MUX2_X2 U4242 ( .A(n2898), .B(n2897), .S(N10), .Z(n2899) );
  MUX2_X2 U4243 ( .A(n2899), .B(n2896), .S(n3181), .Z(n2900) );
  MUX2_X2 U4244 ( .A(n2900), .B(n2893), .S(n3189), .Z(n2901) );
  MUX2_X2 U4245 ( .A(\mem[14][25] ), .B(\mem[15][25] ), .S(n3144), .Z(n2902)
         );
  MUX2_X2 U4246 ( .A(\mem[12][25] ), .B(\mem[13][25] ), .S(n3144), .Z(n2903)
         );
  MUX2_X2 U4247 ( .A(n2903), .B(n2902), .S(N10), .Z(n2904) );
  MUX2_X2 U4248 ( .A(\mem[10][25] ), .B(\mem[11][25] ), .S(n3144), .Z(n2905)
         );
  MUX2_X2 U4249 ( .A(\mem[8][25] ), .B(\mem[9][25] ), .S(n3144), .Z(n2906) );
  MUX2_X2 U4250 ( .A(n2906), .B(n2905), .S(N10), .Z(n2907) );
  MUX2_X2 U4251 ( .A(n2907), .B(n2904), .S(n3181), .Z(n2908) );
  MUX2_X2 U4252 ( .A(\mem[6][25] ), .B(\mem[7][25] ), .S(n3144), .Z(n2909) );
  MUX2_X2 U4253 ( .A(\mem[4][25] ), .B(\mem[5][25] ), .S(n3145), .Z(n2910) );
  MUX2_X2 U4254 ( .A(n2910), .B(n2909), .S(N10), .Z(n2911) );
  MUX2_X2 U4255 ( .A(\mem[2][25] ), .B(\mem[3][25] ), .S(n3145), .Z(n2912) );
  MUX2_X2 U4256 ( .A(\mem[0][25] ), .B(\mem[1][25] ), .S(n3145), .Z(n2913) );
  MUX2_X2 U4257 ( .A(n2913), .B(n2912), .S(N10), .Z(n2914) );
  MUX2_X2 U4258 ( .A(n2914), .B(n2911), .S(n3181), .Z(n2915) );
  MUX2_X2 U4259 ( .A(n2915), .B(n2908), .S(n3189), .Z(n2916) );
  MUX2_X2 U4260 ( .A(n2916), .B(n2901), .S(N13), .Z(rData[25]) );
  MUX2_X2 U4261 ( .A(\mem[30][26] ), .B(\mem[31][26] ), .S(n3145), .Z(n2917)
         );
  MUX2_X2 U4262 ( .A(\mem[28][26] ), .B(\mem[29][26] ), .S(n3145), .Z(n2918)
         );
  MUX2_X2 U4263 ( .A(n2918), .B(n2917), .S(N10), .Z(n2919) );
  MUX2_X2 U4264 ( .A(\mem[26][26] ), .B(\mem[27][26] ), .S(n3145), .Z(n2920)
         );
  MUX2_X2 U4265 ( .A(\mem[24][26] ), .B(\mem[25][26] ), .S(n3145), .Z(n2921)
         );
  MUX2_X2 U4266 ( .A(n2921), .B(n2920), .S(N10), .Z(n2922) );
  MUX2_X2 U4267 ( .A(n2922), .B(n2919), .S(n3181), .Z(n2923) );
  MUX2_X2 U4268 ( .A(\mem[22][26] ), .B(\mem[23][26] ), .S(n3145), .Z(n2924)
         );
  MUX2_X2 U4269 ( .A(\mem[20][26] ), .B(\mem[21][26] ), .S(n3145), .Z(n2925)
         );
  MUX2_X2 U4270 ( .A(n2925), .B(n2924), .S(N10), .Z(n2926) );
  MUX2_X2 U4271 ( .A(\mem[18][26] ), .B(\mem[19][26] ), .S(n3145), .Z(n2927)
         );
  MUX2_X2 U4272 ( .A(\mem[16][26] ), .B(\mem[17][26] ), .S(n3145), .Z(n2928)
         );
  MUX2_X2 U4273 ( .A(n2928), .B(n2927), .S(N10), .Z(n2929) );
  MUX2_X2 U4274 ( .A(n2929), .B(n2926), .S(n3181), .Z(n2930) );
  MUX2_X2 U4275 ( .A(n2930), .B(n2923), .S(n3189), .Z(n2931) );
  MUX2_X2 U4276 ( .A(\mem[14][26] ), .B(\mem[15][26] ), .S(n3146), .Z(n2932)
         );
  MUX2_X2 U4277 ( .A(\mem[12][26] ), .B(\mem[13][26] ), .S(n3146), .Z(n2933)
         );
  MUX2_X2 U4278 ( .A(n2933), .B(n2932), .S(N10), .Z(n2934) );
  MUX2_X2 U4279 ( .A(\mem[10][26] ), .B(\mem[11][26] ), .S(n3146), .Z(n2935)
         );
  MUX2_X2 U4280 ( .A(\mem[8][26] ), .B(\mem[9][26] ), .S(n3146), .Z(n2936) );
  MUX2_X2 U4281 ( .A(n2936), .B(n2935), .S(N10), .Z(n2937) );
  MUX2_X2 U4282 ( .A(n2937), .B(n2934), .S(n3182), .Z(n2938) );
  MUX2_X2 U4283 ( .A(\mem[6][26] ), .B(\mem[7][26] ), .S(n3146), .Z(n2939) );
  MUX2_X2 U4284 ( .A(\mem[4][26] ), .B(\mem[5][26] ), .S(n3146), .Z(n2940) );
  MUX2_X2 U4285 ( .A(n2940), .B(n2939), .S(N10), .Z(n2941) );
  MUX2_X2 U4286 ( .A(\mem[2][26] ), .B(\mem[3][26] ), .S(n3146), .Z(n2942) );
  MUX2_X2 U4287 ( .A(\mem[0][26] ), .B(\mem[1][26] ), .S(n3146), .Z(n2943) );
  MUX2_X2 U4288 ( .A(n2943), .B(n2942), .S(N10), .Z(n2944) );
  MUX2_X2 U4289 ( .A(n2944), .B(n2941), .S(n3182), .Z(n2945) );
  MUX2_X2 U4290 ( .A(n2945), .B(n2938), .S(n3188), .Z(n2946) );
  MUX2_X2 U4291 ( .A(n2946), .B(n2931), .S(N13), .Z(rData[26]) );
  MUX2_X2 U4292 ( .A(\mem[30][27] ), .B(\mem[31][27] ), .S(n3146), .Z(n2947)
         );
  MUX2_X2 U4293 ( .A(\mem[28][27] ), .B(\mem[29][27] ), .S(n3146), .Z(n2948)
         );
  MUX2_X2 U4294 ( .A(n2948), .B(n2947), .S(N10), .Z(n2949) );
  MUX2_X2 U4295 ( .A(\mem[26][27] ), .B(\mem[27][27] ), .S(n3146), .Z(n2950)
         );
  MUX2_X2 U4296 ( .A(\mem[24][27] ), .B(\mem[25][27] ), .S(n3147), .Z(n2951)
         );
  MUX2_X2 U4297 ( .A(n2951), .B(n2950), .S(N10), .Z(n2952) );
  MUX2_X2 U4298 ( .A(n2952), .B(n2949), .S(n3182), .Z(n2953) );
  MUX2_X2 U4299 ( .A(\mem[22][27] ), .B(\mem[23][27] ), .S(n3147), .Z(n2954)
         );
  MUX2_X2 U4300 ( .A(\mem[20][27] ), .B(\mem[21][27] ), .S(n3147), .Z(n2955)
         );
  MUX2_X2 U4301 ( .A(n2955), .B(n2954), .S(N10), .Z(n2956) );
  MUX2_X2 U4302 ( .A(\mem[18][27] ), .B(\mem[19][27] ), .S(n3147), .Z(n2957)
         );
  MUX2_X2 U4303 ( .A(\mem[16][27] ), .B(\mem[17][27] ), .S(n3147), .Z(n2958)
         );
  MUX2_X2 U4304 ( .A(n2958), .B(n2957), .S(N10), .Z(n2959) );
  MUX2_X2 U4305 ( .A(n2959), .B(n2956), .S(n3182), .Z(n2960) );
  MUX2_X2 U4306 ( .A(n2960), .B(n2953), .S(n3189), .Z(n2961) );
  MUX2_X2 U4307 ( .A(\mem[14][27] ), .B(\mem[15][27] ), .S(n3147), .Z(n2962)
         );
  MUX2_X2 U4308 ( .A(\mem[12][27] ), .B(\mem[13][27] ), .S(n3147), .Z(n2963)
         );
  MUX2_X2 U4309 ( .A(n2963), .B(n2962), .S(N10), .Z(n2964) );
  MUX2_X2 U4310 ( .A(\mem[10][27] ), .B(\mem[11][27] ), .S(n3147), .Z(n2965)
         );
  MUX2_X2 U4311 ( .A(\mem[8][27] ), .B(\mem[9][27] ), .S(n3147), .Z(n2966) );
  MUX2_X2 U4312 ( .A(n2966), .B(n2965), .S(N10), .Z(n2967) );
  MUX2_X2 U4313 ( .A(n2967), .B(n2964), .S(n3182), .Z(n2968) );
  MUX2_X2 U4314 ( .A(\mem[6][27] ), .B(\mem[7][27] ), .S(n3147), .Z(n2969) );
  MUX2_X2 U4315 ( .A(\mem[4][27] ), .B(\mem[5][27] ), .S(n3147), .Z(n2970) );
  MUX2_X2 U4316 ( .A(n2970), .B(n2969), .S(N10), .Z(n2971) );
  MUX2_X2 U4317 ( .A(\mem[2][27] ), .B(\mem[3][27] ), .S(n3148), .Z(n2972) );
  MUX2_X2 U4318 ( .A(\mem[0][27] ), .B(\mem[1][27] ), .S(n3148), .Z(n2973) );
  MUX2_X2 U4319 ( .A(n2973), .B(n2972), .S(N10), .Z(n2974) );
  MUX2_X2 U4320 ( .A(n2974), .B(n2971), .S(n3182), .Z(n2975) );
  MUX2_X2 U4321 ( .A(n2975), .B(n2968), .S(n3189), .Z(n2976) );
  MUX2_X2 U4322 ( .A(n2976), .B(n2961), .S(N13), .Z(rData[27]) );
  MUX2_X2 U4323 ( .A(\mem[30][28] ), .B(\mem[31][28] ), .S(n3148), .Z(n2977)
         );
  MUX2_X2 U4324 ( .A(\mem[28][28] ), .B(\mem[29][28] ), .S(n3148), .Z(n2978)
         );
  MUX2_X2 U4325 ( .A(n2978), .B(n2977), .S(N10), .Z(n2979) );
  MUX2_X2 U4326 ( .A(\mem[26][28] ), .B(\mem[27][28] ), .S(n3148), .Z(n2980)
         );
  MUX2_X2 U4327 ( .A(\mem[24][28] ), .B(\mem[25][28] ), .S(n3148), .Z(n2981)
         );
  MUX2_X2 U4328 ( .A(n2981), .B(n2980), .S(N10), .Z(n2982) );
  MUX2_X2 U4329 ( .A(n2982), .B(n2979), .S(n3182), .Z(n2983) );
  MUX2_X2 U4330 ( .A(\mem[22][28] ), .B(\mem[23][28] ), .S(n3148), .Z(n2984)
         );
  MUX2_X2 U4331 ( .A(\mem[20][28] ), .B(\mem[21][28] ), .S(n3148), .Z(n2985)
         );
  MUX2_X2 U4332 ( .A(n2985), .B(n2984), .S(N10), .Z(n2986) );
  MUX2_X2 U4333 ( .A(\mem[18][28] ), .B(\mem[19][28] ), .S(n3148), .Z(n2987)
         );
  MUX2_X2 U4334 ( .A(\mem[16][28] ), .B(\mem[17][28] ), .S(n3148), .Z(n2988)
         );
  MUX2_X2 U4335 ( .A(n2988), .B(n2987), .S(N10), .Z(n2989) );
  MUX2_X2 U4336 ( .A(n2989), .B(n2986), .S(n3182), .Z(n2990) );
  MUX2_X2 U4337 ( .A(n2990), .B(n2983), .S(n3188), .Z(n2991) );
  MUX2_X2 U4338 ( .A(\mem[14][28] ), .B(\mem[15][28] ), .S(n3148), .Z(n2992)
         );
  MUX2_X2 U4339 ( .A(\mem[12][28] ), .B(\mem[13][28] ), .S(n3149), .Z(n2993)
         );
  MUX2_X2 U4340 ( .A(n2993), .B(n2992), .S(N10), .Z(n2994) );
  MUX2_X2 U4341 ( .A(\mem[10][28] ), .B(\mem[11][28] ), .S(n3149), .Z(n2995)
         );
  MUX2_X2 U4342 ( .A(\mem[8][28] ), .B(\mem[9][28] ), .S(n3149), .Z(n2996) );
  MUX2_X2 U4343 ( .A(n2996), .B(n2995), .S(N10), .Z(n2997) );
  MUX2_X2 U4344 ( .A(n2997), .B(n2994), .S(n3182), .Z(n2998) );
  MUX2_X2 U4345 ( .A(\mem[6][28] ), .B(\mem[7][28] ), .S(n3149), .Z(n2999) );
  MUX2_X2 U4346 ( .A(\mem[4][28] ), .B(\mem[5][28] ), .S(n3149), .Z(n3000) );
  MUX2_X2 U4347 ( .A(n3000), .B(n2999), .S(N10), .Z(n3001) );
  MUX2_X2 U4348 ( .A(\mem[2][28] ), .B(\mem[3][28] ), .S(n3149), .Z(n3002) );
  MUX2_X2 U4349 ( .A(\mem[0][28] ), .B(\mem[1][28] ), .S(n3149), .Z(n3003) );
  MUX2_X2 U4350 ( .A(n3003), .B(n3002), .S(N10), .Z(n3004) );
  MUX2_X2 U4351 ( .A(n3004), .B(n3001), .S(n3182), .Z(n3005) );
  MUX2_X2 U4352 ( .A(n3005), .B(n2998), .S(n3188), .Z(n3006) );
  MUX2_X2 U4353 ( .A(n3006), .B(n2991), .S(N13), .Z(rData[28]) );
  MUX2_X2 U4354 ( .A(\mem[30][29] ), .B(\mem[31][29] ), .S(n3149), .Z(n3007)
         );
  MUX2_X2 U4355 ( .A(\mem[28][29] ), .B(\mem[29][29] ), .S(n3149), .Z(n3008)
         );
  MUX2_X2 U4356 ( .A(n3008), .B(n3007), .S(N10), .Z(n3009) );
  MUX2_X2 U4357 ( .A(\mem[26][29] ), .B(\mem[27][29] ), .S(n3149), .Z(n3010)
         );
  MUX2_X2 U4358 ( .A(\mem[24][29] ), .B(\mem[25][29] ), .S(n3149), .Z(n3011)
         );
  MUX2_X2 U4359 ( .A(n3011), .B(n3010), .S(N10), .Z(n3012) );
  MUX2_X2 U4360 ( .A(n3012), .B(n3009), .S(n3182), .Z(n3013) );
  MUX2_X2 U4361 ( .A(\mem[22][29] ), .B(\mem[23][29] ), .S(n3150), .Z(n3014)
         );
  MUX2_X2 U4362 ( .A(\mem[20][29] ), .B(\mem[21][29] ), .S(n3150), .Z(n3015)
         );
  MUX2_X2 U4363 ( .A(n3015), .B(n3014), .S(N10), .Z(n3016) );
  MUX2_X2 U4364 ( .A(\mem[18][29] ), .B(\mem[19][29] ), .S(n3150), .Z(n3017)
         );
  MUX2_X2 U4365 ( .A(\mem[16][29] ), .B(\mem[17][29] ), .S(n3150), .Z(n3018)
         );
  MUX2_X2 U4366 ( .A(n3018), .B(n3017), .S(N10), .Z(n3019) );
  MUX2_X2 U4367 ( .A(n3019), .B(n3016), .S(n3175), .Z(n3020) );
  MUX2_X2 U4368 ( .A(n3020), .B(n3013), .S(n3189), .Z(n3021) );
  MUX2_X2 U4369 ( .A(\mem[14][29] ), .B(\mem[15][29] ), .S(n3150), .Z(n3022)
         );
  MUX2_X2 U4370 ( .A(\mem[12][29] ), .B(\mem[13][29] ), .S(n3150), .Z(n3023)
         );
  MUX2_X2 U4371 ( .A(n3023), .B(n3022), .S(N10), .Z(n3024) );
  MUX2_X2 U4372 ( .A(\mem[10][29] ), .B(\mem[11][29] ), .S(n3150), .Z(n3025)
         );
  MUX2_X2 U4373 ( .A(\mem[8][29] ), .B(\mem[9][29] ), .S(n3150), .Z(n3026) );
  MUX2_X2 U4374 ( .A(n3026), .B(n3025), .S(N10), .Z(n3027) );
  MUX2_X2 U4375 ( .A(n3027), .B(n3024), .S(n3176), .Z(n3028) );
  MUX2_X2 U4376 ( .A(\mem[6][29] ), .B(\mem[7][29] ), .S(n3150), .Z(n3029) );
  MUX2_X2 U4377 ( .A(\mem[4][29] ), .B(\mem[5][29] ), .S(n3150), .Z(n3030) );
  MUX2_X2 U4378 ( .A(n3030), .B(n3029), .S(N10), .Z(n3031) );
  MUX2_X2 U4379 ( .A(\mem[2][29] ), .B(\mem[3][29] ), .S(n3150), .Z(n3032) );
  MUX2_X2 U4380 ( .A(\mem[0][29] ), .B(\mem[1][29] ), .S(n3151), .Z(n3033) );
  MUX2_X2 U4381 ( .A(n3033), .B(n3032), .S(N10), .Z(n3034) );
  MUX2_X2 U4382 ( .A(n3034), .B(n3031), .S(n3176), .Z(n3035) );
  MUX2_X2 U4383 ( .A(n3035), .B(n3028), .S(n3189), .Z(n3036) );
  MUX2_X2 U4384 ( .A(n3036), .B(n3021), .S(N13), .Z(rData[29]) );
  MUX2_X2 U4385 ( .A(\mem[30][30] ), .B(\mem[31][30] ), .S(n3151), .Z(n3037)
         );
  MUX2_X2 U4386 ( .A(\mem[28][30] ), .B(\mem[29][30] ), .S(n3151), .Z(n3038)
         );
  MUX2_X2 U4387 ( .A(n3038), .B(n3037), .S(N10), .Z(n3039) );
  MUX2_X2 U4388 ( .A(\mem[26][30] ), .B(\mem[27][30] ), .S(n3151), .Z(n3040)
         );
  MUX2_X2 U4389 ( .A(\mem[24][30] ), .B(\mem[25][30] ), .S(n3151), .Z(n3041)
         );
  MUX2_X2 U4390 ( .A(n3041), .B(n3040), .S(N10), .Z(n3042) );
  MUX2_X2 U4391 ( .A(n3042), .B(n3039), .S(n3176), .Z(n3043) );
  MUX2_X2 U4392 ( .A(\mem[22][30] ), .B(\mem[23][30] ), .S(n3151), .Z(n3044)
         );
  MUX2_X2 U4393 ( .A(\mem[20][30] ), .B(\mem[21][30] ), .S(n3151), .Z(n3045)
         );
  MUX2_X2 U4394 ( .A(n3045), .B(n3044), .S(N10), .Z(n3046) );
  MUX2_X2 U4395 ( .A(\mem[18][30] ), .B(\mem[19][30] ), .S(n3151), .Z(n3047)
         );
  MUX2_X2 U4396 ( .A(\mem[16][30] ), .B(\mem[17][30] ), .S(n3151), .Z(n3048)
         );
  MUX2_X2 U4397 ( .A(n3048), .B(n3047), .S(N10), .Z(n3049) );
  MUX2_X2 U4398 ( .A(n3049), .B(n3046), .S(n3176), .Z(n3050) );
  MUX2_X2 U4399 ( .A(n3050), .B(n3043), .S(n3188), .Z(n3051) );
  MUX2_X2 U4400 ( .A(\mem[14][30] ), .B(\mem[15][30] ), .S(n3151), .Z(n3052)
         );
  MUX2_X2 U4401 ( .A(\mem[12][30] ), .B(\mem[13][30] ), .S(n3151), .Z(n3053)
         );
  MUX2_X2 U4402 ( .A(n3053), .B(n3052), .S(N10), .Z(n3054) );
  MUX2_X2 U4403 ( .A(\mem[10][30] ), .B(\mem[11][30] ), .S(n3152), .Z(n3055)
         );
  MUX2_X2 U4404 ( .A(\mem[8][30] ), .B(\mem[9][30] ), .S(n3152), .Z(n3056) );
  MUX2_X2 U4405 ( .A(n3056), .B(n3055), .S(N10), .Z(n3057) );
  MUX2_X2 U4406 ( .A(n3057), .B(n3054), .S(n3175), .Z(n3058) );
  MUX2_X2 U4407 ( .A(\mem[6][30] ), .B(\mem[7][30] ), .S(n3152), .Z(n3059) );
  MUX2_X2 U4408 ( .A(\mem[4][30] ), .B(\mem[5][30] ), .S(n3152), .Z(n3060) );
  MUX2_X2 U4409 ( .A(n3060), .B(n3059), .S(N10), .Z(n3061) );
  MUX2_X2 U4410 ( .A(\mem[2][30] ), .B(\mem[3][30] ), .S(n3152), .Z(n3062) );
  MUX2_X2 U4411 ( .A(\mem[0][30] ), .B(\mem[1][30] ), .S(n3152), .Z(n3063) );
  MUX2_X2 U4412 ( .A(n3063), .B(n3062), .S(N10), .Z(n3064) );
  MUX2_X2 U4413 ( .A(n3064), .B(n3061), .S(n3175), .Z(n3065) );
  MUX2_X2 U4414 ( .A(n3065), .B(n3058), .S(n3188), .Z(n3066) );
  MUX2_X2 U4415 ( .A(n3066), .B(n3051), .S(N13), .Z(rData[30]) );
  MUX2_X2 U4416 ( .A(\mem[30][31] ), .B(\mem[31][31] ), .S(n3152), .Z(n3067)
         );
  MUX2_X2 U4417 ( .A(\mem[28][31] ), .B(\mem[29][31] ), .S(n3152), .Z(n3068)
         );
  MUX2_X2 U4418 ( .A(n3068), .B(n3067), .S(N10), .Z(n3069) );
  MUX2_X2 U4419 ( .A(\mem[26][31] ), .B(\mem[27][31] ), .S(n3152), .Z(n3070)
         );
  MUX2_X2 U4420 ( .A(\mem[24][31] ), .B(\mem[25][31] ), .S(n3152), .Z(n3071)
         );
  MUX2_X2 U4421 ( .A(n3071), .B(n3070), .S(N10), .Z(n3072) );
  MUX2_X2 U4422 ( .A(n3072), .B(n3069), .S(n3175), .Z(n3073) );
  MUX2_X2 U4423 ( .A(\mem[22][31] ), .B(\mem[23][31] ), .S(n3152), .Z(n3074)
         );
  MUX2_X2 U4424 ( .A(\mem[20][31] ), .B(\mem[21][31] ), .S(n3153), .Z(n3075)
         );
  MUX2_X2 U4425 ( .A(n3075), .B(n3074), .S(N10), .Z(n3076) );
  MUX2_X2 U4426 ( .A(\mem[18][31] ), .B(\mem[19][31] ), .S(n3153), .Z(n3077)
         );
  MUX2_X2 U4427 ( .A(\mem[16][31] ), .B(\mem[17][31] ), .S(n3153), .Z(n3078)
         );
  MUX2_X2 U4428 ( .A(n3078), .B(n3077), .S(N10), .Z(n3079) );
  MUX2_X2 U4429 ( .A(n3079), .B(n3076), .S(n3175), .Z(n3080) );
  MUX2_X2 U4430 ( .A(n3080), .B(n3073), .S(n3189), .Z(n3081) );
  MUX2_X2 U4431 ( .A(\mem[14][31] ), .B(\mem[15][31] ), .S(n3153), .Z(n3082)
         );
  MUX2_X2 U4432 ( .A(\mem[12][31] ), .B(\mem[13][31] ), .S(n3153), .Z(n3083)
         );
  MUX2_X2 U4433 ( .A(n3083), .B(n3082), .S(N10), .Z(n3084) );
  MUX2_X2 U4434 ( .A(\mem[10][31] ), .B(\mem[11][31] ), .S(n3153), .Z(n3085)
         );
  MUX2_X2 U4435 ( .A(\mem[8][31] ), .B(\mem[9][31] ), .S(n3153), .Z(n3086) );
  MUX2_X2 U4436 ( .A(n3086), .B(n3085), .S(N10), .Z(n3087) );
  MUX2_X2 U4437 ( .A(n3087), .B(n3084), .S(n3176), .Z(n3088) );
  MUX2_X2 U4438 ( .A(\mem[6][31] ), .B(\mem[7][31] ), .S(n3153), .Z(n3089) );
  MUX2_X2 U4439 ( .A(\mem[4][31] ), .B(\mem[5][31] ), .S(n3153), .Z(n3090) );
  MUX2_X2 U4440 ( .A(n3090), .B(n3089), .S(N10), .Z(n3091) );
  MUX2_X2 U4441 ( .A(\mem[2][31] ), .B(\mem[3][31] ), .S(n3153), .Z(n3092) );
  MUX2_X2 U4442 ( .A(\mem[0][31] ), .B(\mem[1][31] ), .S(n3153), .Z(n3093) );
  MUX2_X2 U4443 ( .A(n3093), .B(n3092), .S(N10), .Z(n3094) );
  MUX2_X2 U4444 ( .A(n3094), .B(n3091), .S(n3176), .Z(n3095) );
  MUX2_X2 U4445 ( .A(n3095), .B(n3088), .S(n3189), .Z(n3096) );
  MUX2_X2 U4446 ( .A(n3096), .B(n3081), .S(N13), .Z(rData[31]) );
  INV_X4 U4447 ( .A(rd[4]), .ZN(n4406) );
  INV_X4 U4448 ( .A(rd[3]), .ZN(n4407) );
  INV_X4 U4449 ( .A(rd[2]), .ZN(n4408) );
  INV_X4 U4450 ( .A(rd[0]), .ZN(n4409) );
  INV_X4 U4451 ( .A(regWr), .ZN(n4410) );
endmodule

