
// NOT GATE



module not_gate (a, z);

// Ports

input a;
output z;

// Implementation

assign z = ~a;
endmodule
