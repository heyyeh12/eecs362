
module regfile ( rs1, rs2, rd, rData1, rData2, wData, regWr, clk );
  input [4:0] rs1;
  input [4:0] rs2;
  input [4:0] rd;
  output [31:0] rData1;
  output [31:0] rData2;
  input [31:0] wData;
  input regWr, clk;
  wire   mem_15__31_, mem_15__30_, mem_15__29_, mem_15__28_, mem_15__27_,
         mem_15__26_, mem_15__25_, mem_15__24_, mem_15__23_, mem_15__22_,
         mem_15__21_, mem_15__20_, mem_15__19_, mem_15__18_, mem_15__17_,
         mem_15__16_, mem_15__15_, mem_15__14_, mem_15__13_, mem_15__12_,
         mem_15__11_, mem_15__10_, mem_15__9_, mem_15__8_, mem_15__7_,
         mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_, mem_15__2_,
         mem_15__1_, mem_15__0_, mem_14__31_, mem_14__30_, mem_14__29_,
         mem_14__28_, mem_14__27_, mem_14__26_, mem_14__25_, mem_14__24_,
         mem_14__23_, mem_14__22_, mem_14__21_, mem_14__20_, mem_14__19_,
         mem_14__18_, mem_14__17_, mem_14__16_, mem_14__15_, mem_14__14_,
         mem_14__13_, mem_14__12_, mem_14__11_, mem_14__10_, mem_14__9_,
         mem_14__8_, mem_14__7_, mem_14__6_, mem_14__5_, mem_14__4_,
         mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_, mem_13__31_,
         mem_13__30_, mem_13__29_, mem_13__28_, mem_13__27_, mem_13__26_,
         mem_13__25_, mem_13__24_, mem_13__23_, mem_13__22_, mem_13__21_,
         mem_13__20_, mem_13__19_, mem_13__18_, mem_13__17_, mem_13__16_,
         mem_13__15_, mem_13__14_, mem_13__13_, mem_13__12_, mem_13__11_,
         mem_13__10_, mem_13__9_, mem_13__8_, mem_13__7_, mem_13__6_,
         mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_, mem_13__1_,
         mem_13__0_, mem_12__31_, mem_12__30_, mem_12__29_, mem_12__28_,
         mem_12__27_, mem_12__26_, mem_12__25_, mem_12__24_, mem_12__23_,
         mem_12__22_, mem_12__21_, mem_12__20_, mem_12__19_, mem_12__18_,
         mem_12__17_, mem_12__16_, mem_12__15_, mem_12__14_, mem_12__13_,
         mem_12__12_, mem_12__11_, mem_12__10_, mem_12__9_, mem_12__8_,
         mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_, mem_12__3_,
         mem_12__2_, mem_12__1_, mem_12__0_, mem_11__31_, mem_11__30_,
         mem_11__29_, mem_11__28_, mem_11__27_, mem_11__26_, mem_11__25_,
         mem_11__24_, mem_11__23_, mem_11__22_, mem_11__21_, mem_11__20_,
         mem_11__19_, mem_11__18_, mem_11__17_, mem_11__16_, mem_11__15_,
         mem_11__14_, mem_11__13_, mem_11__12_, mem_11__11_, mem_11__10_,
         mem_11__9_, mem_11__8_, mem_11__7_, mem_11__6_, mem_11__5_,
         mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_, mem_11__0_,
         mem_10__31_, mem_10__30_, mem_10__29_, mem_10__28_, mem_10__27_,
         mem_10__26_, mem_10__25_, mem_10__24_, mem_10__23_, mem_10__22_,
         mem_10__21_, mem_10__20_, mem_10__19_, mem_10__18_, mem_10__17_,
         mem_10__16_, mem_10__15_, mem_10__14_, mem_10__13_, mem_10__12_,
         mem_10__11_, mem_10__10_, mem_10__9_, mem_10__8_, mem_10__7_,
         mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_, mem_10__2_,
         mem_10__1_, mem_10__0_, mem_9__31_, mem_9__30_, mem_9__29_,
         mem_9__28_, mem_9__27_, mem_9__26_, mem_9__25_, mem_9__24_,
         mem_9__23_, mem_9__22_, mem_9__21_, mem_9__20_, mem_9__19_,
         mem_9__18_, mem_9__17_, mem_9__16_, mem_9__15_, mem_9__14_,
         mem_9__13_, mem_9__12_, mem_9__11_, mem_9__10_, mem_9__9_, mem_9__8_,
         mem_9__7_, mem_9__6_, mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_,
         mem_9__1_, mem_9__0_, mem_8__31_, mem_8__30_, mem_8__29_, mem_8__28_,
         mem_8__27_, mem_8__26_, mem_8__25_, mem_8__24_, mem_8__23_,
         mem_8__22_, mem_8__21_, mem_8__20_, mem_8__19_, mem_8__18_,
         mem_8__17_, mem_8__16_, mem_8__15_, mem_8__14_, mem_8__13_,
         mem_8__12_, mem_8__11_, mem_8__10_, mem_8__9_, mem_8__8_, mem_8__7_,
         mem_8__6_, mem_8__5_, mem_8__4_, mem_8__3_, mem_8__2_, mem_8__1_,
         mem_8__0_, mem_7__31_, mem_7__30_, mem_7__29_, mem_7__28_, mem_7__27_,
         mem_7__26_, mem_7__25_, mem_7__24_, mem_7__23_, mem_7__22_,
         mem_7__21_, mem_7__20_, mem_7__19_, mem_7__18_, mem_7__17_,
         mem_7__16_, mem_7__15_, mem_7__14_, mem_7__13_, mem_7__12_,
         mem_7__11_, mem_7__10_, mem_7__9_, mem_7__8_, mem_7__7_, mem_7__6_,
         mem_7__5_, mem_7__4_, mem_7__3_, mem_7__2_, mem_7__1_, mem_7__0_,
         mem_6__31_, mem_6__30_, mem_6__29_, mem_6__28_, mem_6__27_,
         mem_6__26_, mem_6__25_, mem_6__24_, mem_6__23_, mem_6__22_,
         mem_6__21_, mem_6__20_, mem_6__19_, mem_6__18_, mem_6__17_,
         mem_6__16_, mem_6__15_, mem_6__14_, mem_6__13_, mem_6__12_,
         mem_6__11_, mem_6__10_, mem_6__9_, mem_6__8_, mem_6__7_, mem_6__6_,
         mem_6__5_, mem_6__4_, mem_6__3_, mem_6__2_, mem_6__1_, mem_6__0_,
         mem_5__31_, mem_5__30_, mem_5__29_, mem_5__28_, mem_5__27_,
         mem_5__26_, mem_5__25_, mem_5__24_, mem_5__23_, mem_5__22_,
         mem_5__21_, mem_5__20_, mem_5__19_, mem_5__18_, mem_5__17_,
         mem_5__16_, mem_5__15_, mem_5__14_, mem_5__13_, mem_5__12_,
         mem_5__11_, mem_5__10_, mem_5__9_, mem_5__8_, mem_5__7_, mem_5__6_,
         mem_5__5_, mem_5__4_, mem_5__3_, mem_5__2_, mem_5__1_, mem_5__0_,
         mem_4__31_, mem_4__30_, mem_4__29_, mem_4__28_, mem_4__27_,
         mem_4__26_, mem_4__25_, mem_4__24_, mem_4__23_, mem_4__22_,
         mem_4__21_, mem_4__20_, mem_4__19_, mem_4__18_, mem_4__17_,
         mem_4__16_, mem_4__15_, mem_4__14_, mem_4__13_, mem_4__12_,
         mem_4__11_, mem_4__10_, mem_4__9_, mem_4__8_, mem_4__7_, mem_4__6_,
         mem_4__5_, mem_4__4_, mem_4__3_, mem_4__2_, mem_4__1_, mem_4__0_,
         mem_3__31_, mem_3__30_, mem_3__29_, mem_3__28_, mem_3__27_,
         mem_3__26_, mem_3__25_, mem_3__24_, mem_3__23_, mem_3__22_,
         mem_3__21_, mem_3__20_, mem_3__19_, mem_3__18_, mem_3__17_,
         mem_3__16_, mem_3__15_, mem_3__14_, mem_3__13_, mem_3__12_,
         mem_3__11_, mem_3__10_, mem_3__9_, mem_3__8_, mem_3__7_, mem_3__6_,
         mem_3__5_, mem_3__4_, mem_3__3_, mem_3__2_, mem_3__1_, mem_3__0_,
         mem_2__31_, mem_2__30_, mem_2__29_, mem_2__28_, mem_2__27_,
         mem_2__26_, mem_2__25_, mem_2__24_, mem_2__23_, mem_2__22_,
         mem_2__21_, mem_2__20_, mem_2__19_, mem_2__18_, mem_2__17_,
         mem_2__16_, mem_2__15_, mem_2__14_, mem_2__13_, mem_2__12_,
         mem_2__11_, mem_2__10_, mem_2__9_, mem_2__8_, mem_2__7_, mem_2__6_,
         mem_2__5_, mem_2__4_, mem_2__3_, mem_2__2_, mem_2__1_, mem_2__0_,
         mem_1__31_, mem_1__30_, mem_1__29_, mem_1__28_, mem_1__27_,
         mem_1__26_, mem_1__25_, mem_1__24_, mem_1__23_, mem_1__22_,
         mem_1__21_, mem_1__20_, mem_1__19_, mem_1__18_, mem_1__17_,
         mem_1__16_, mem_1__15_, mem_1__14_, mem_1__13_, mem_1__12_,
         mem_1__11_, mem_1__10_, mem_1__9_, mem_1__8_, mem_1__7_, mem_1__6_,
         mem_1__5_, mem_1__4_, mem_1__3_, mem_1__2_, mem_1__1_, mem_1__0_,
         mem_0__31_, mem_0__30_, mem_0__29_, mem_0__28_, mem_0__27_,
         mem_0__26_, mem_0__25_, mem_0__24_, mem_0__23_, mem_0__22_,
         mem_0__21_, mem_0__20_, mem_0__19_, mem_0__18_, mem_0__17_,
         mem_0__16_, mem_0__15_, mem_0__14_, mem_0__13_, mem_0__12_,
         mem_0__11_, mem_0__10_, mem_0__9_, mem_0__8_, mem_0__7_, mem_0__6_,
         mem_0__5_, mem_0__4_, mem_0__3_, mem_0__2_, mem_0__1_, mem_0__0_,
         mem_31__31_, mem_31__30_, mem_31__29_, mem_31__28_, mem_31__27_,
         mem_31__26_, mem_31__25_, mem_31__24_, mem_31__23_, mem_31__22_,
         mem_31__21_, mem_31__20_, mem_31__19_, mem_31__18_, mem_31__17_,
         mem_31__16_, mem_31__15_, mem_31__14_, mem_31__13_, mem_31__12_,
         mem_31__11_, mem_31__10_, mem_31__9_, mem_31__8_, mem_31__7_,
         mem_31__6_, mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_,
         mem_31__1_, mem_31__0_, mem_30__31_, mem_30__30_, mem_30__29_,
         mem_30__28_, mem_30__27_, mem_30__26_, mem_30__25_, mem_30__24_,
         mem_30__23_, mem_30__22_, mem_30__21_, mem_30__20_, mem_30__19_,
         mem_30__18_, mem_30__17_, mem_30__16_, mem_30__15_, mem_30__14_,
         mem_30__13_, mem_30__12_, mem_30__11_, mem_30__10_, mem_30__9_,
         mem_30__8_, mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_,
         mem_30__3_, mem_30__2_, mem_30__1_, mem_30__0_, mem_29__31_,
         mem_29__30_, mem_29__29_, mem_29__28_, mem_29__27_, mem_29__26_,
         mem_29__25_, mem_29__24_, mem_29__23_, mem_29__22_, mem_29__21_,
         mem_29__20_, mem_29__19_, mem_29__18_, mem_29__17_, mem_29__16_,
         mem_29__15_, mem_29__14_, mem_29__13_, mem_29__12_, mem_29__11_,
         mem_29__10_, mem_29__9_, mem_29__8_, mem_29__7_, mem_29__6_,
         mem_29__5_, mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_,
         mem_29__0_, mem_28__31_, mem_28__30_, mem_28__29_, mem_28__28_,
         mem_28__27_, mem_28__26_, mem_28__25_, mem_28__24_, mem_28__23_,
         mem_28__22_, mem_28__21_, mem_28__20_, mem_28__19_, mem_28__18_,
         mem_28__17_, mem_28__16_, mem_28__15_, mem_28__14_, mem_28__13_,
         mem_28__12_, mem_28__11_, mem_28__10_, mem_28__9_, mem_28__8_,
         mem_28__7_, mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_,
         mem_28__2_, mem_28__1_, mem_28__0_, mem_27__31_, mem_27__30_,
         mem_27__29_, mem_27__28_, mem_27__27_, mem_27__26_, mem_27__25_,
         mem_27__24_, mem_27__23_, mem_27__22_, mem_27__21_, mem_27__20_,
         mem_27__19_, mem_27__18_, mem_27__17_, mem_27__16_, mem_27__15_,
         mem_27__14_, mem_27__13_, mem_27__12_, mem_27__11_, mem_27__10_,
         mem_27__9_, mem_27__8_, mem_27__7_, mem_27__6_, mem_27__5_,
         mem_27__4_, mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_,
         mem_26__31_, mem_26__30_, mem_26__29_, mem_26__28_, mem_26__27_,
         mem_26__26_, mem_26__25_, mem_26__24_, mem_26__23_, mem_26__22_,
         mem_26__21_, mem_26__20_, mem_26__19_, mem_26__18_, mem_26__17_,
         mem_26__16_, mem_26__15_, mem_26__14_, mem_26__13_, mem_26__12_,
         mem_26__11_, mem_26__10_, mem_26__9_, mem_26__8_, mem_26__7_,
         mem_26__6_, mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_,
         mem_26__1_, mem_26__0_, mem_25__31_, mem_25__30_, mem_25__29_,
         mem_25__28_, mem_25__27_, mem_25__26_, mem_25__25_, mem_25__24_,
         mem_25__23_, mem_25__22_, mem_25__21_, mem_25__20_, mem_25__19_,
         mem_25__18_, mem_25__17_, mem_25__16_, mem_25__15_, mem_25__14_,
         mem_25__13_, mem_25__12_, mem_25__11_, mem_25__10_, mem_25__9_,
         mem_25__8_, mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_,
         mem_25__3_, mem_25__2_, mem_25__1_, mem_25__0_, mem_24__31_,
         mem_24__30_, mem_24__29_, mem_24__28_, mem_24__27_, mem_24__26_,
         mem_24__25_, mem_24__24_, mem_24__23_, mem_24__22_, mem_24__21_,
         mem_24__20_, mem_24__19_, mem_24__18_, mem_24__17_, mem_24__16_,
         mem_24__15_, mem_24__14_, mem_24__13_, mem_24__12_, mem_24__11_,
         mem_24__10_, mem_24__9_, mem_24__8_, mem_24__7_, mem_24__6_,
         mem_24__5_, mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_,
         mem_24__0_, mem_23__31_, mem_23__30_, mem_23__29_, mem_23__28_,
         mem_23__27_, mem_23__26_, mem_23__25_, mem_23__24_, mem_23__23_,
         mem_23__22_, mem_23__21_, mem_23__20_, mem_23__19_, mem_23__18_,
         mem_23__17_, mem_23__16_, mem_23__15_, mem_23__14_, mem_23__13_,
         mem_23__12_, mem_23__11_, mem_23__10_, mem_23__9_, mem_23__8_,
         mem_23__7_, mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_,
         mem_23__2_, mem_23__1_, mem_23__0_, mem_22__31_, mem_22__30_,
         mem_22__29_, mem_22__28_, mem_22__27_, mem_22__26_, mem_22__25_,
         mem_22__24_, mem_22__23_, mem_22__22_, mem_22__21_, mem_22__20_,
         mem_22__19_, mem_22__18_, mem_22__17_, mem_22__16_, mem_22__15_,
         mem_22__14_, mem_22__13_, mem_22__12_, mem_22__11_, mem_22__10_,
         mem_22__9_, mem_22__8_, mem_22__7_, mem_22__6_, mem_22__5_,
         mem_22__4_, mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_,
         mem_21__31_, mem_21__30_, mem_21__29_, mem_21__28_, mem_21__27_,
         mem_21__26_, mem_21__25_, mem_21__24_, mem_21__23_, mem_21__22_,
         mem_21__21_, mem_21__20_, mem_21__19_, mem_21__18_, mem_21__17_,
         mem_21__16_, mem_21__15_, mem_21__14_, mem_21__13_, mem_21__12_,
         mem_21__11_, mem_21__10_, mem_21__9_, mem_21__8_, mem_21__7_,
         mem_21__6_, mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_,
         mem_21__1_, mem_21__0_, mem_20__31_, mem_20__30_, mem_20__29_,
         mem_20__28_, mem_20__27_, mem_20__26_, mem_20__25_, mem_20__24_,
         mem_20__23_, mem_20__22_, mem_20__21_, mem_20__20_, mem_20__19_,
         mem_20__18_, mem_20__17_, mem_20__16_, mem_20__15_, mem_20__14_,
         mem_20__13_, mem_20__12_, mem_20__11_, mem_20__10_, mem_20__9_,
         mem_20__8_, mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_,
         mem_20__3_, mem_20__2_, mem_20__1_, mem_20__0_, mem_19__31_,
         mem_19__30_, mem_19__29_, mem_19__28_, mem_19__27_, mem_19__26_,
         mem_19__25_, mem_19__24_, mem_19__23_, mem_19__22_, mem_19__21_,
         mem_19__20_, mem_19__19_, mem_19__18_, mem_19__17_, mem_19__16_,
         mem_19__15_, mem_19__14_, mem_19__13_, mem_19__12_, mem_19__11_,
         mem_19__10_, mem_19__9_, mem_19__8_, mem_19__7_, mem_19__6_,
         mem_19__5_, mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_,
         mem_19__0_, mem_18__31_, mem_18__30_, mem_18__29_, mem_18__28_,
         mem_18__27_, mem_18__26_, mem_18__25_, mem_18__24_, mem_18__23_,
         mem_18__22_, mem_18__21_, mem_18__20_, mem_18__19_, mem_18__18_,
         mem_18__17_, mem_18__16_, mem_18__15_, mem_18__14_, mem_18__13_,
         mem_18__12_, mem_18__11_, mem_18__10_, mem_18__9_, mem_18__8_,
         mem_18__7_, mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_,
         mem_18__2_, mem_18__1_, mem_18__0_, mem_17__31_, mem_17__30_,
         mem_17__29_, mem_17__28_, mem_17__27_, mem_17__26_, mem_17__25_,
         mem_17__24_, mem_17__23_, mem_17__22_, mem_17__21_, mem_17__20_,
         mem_17__19_, mem_17__18_, mem_17__17_, mem_17__16_, mem_17__15_,
         mem_17__14_, mem_17__13_, mem_17__12_, mem_17__11_, mem_17__10_,
         mem_17__9_, mem_17__8_, mem_17__7_, mem_17__6_, mem_17__5_,
         mem_17__4_, mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_,
         mem_16__31_, mem_16__30_, mem_16__29_, mem_16__28_, mem_16__27_,
         mem_16__26_, mem_16__25_, mem_16__24_, mem_16__23_, mem_16__22_,
         mem_16__21_, mem_16__20_, mem_16__19_, mem_16__18_, mem_16__17_,
         mem_16__16_, mem_16__15_, mem_16__14_, mem_16__13_, mem_16__12_,
         mem_16__11_, mem_16__10_, mem_16__9_, mem_16__8_, mem_16__7_,
         mem_16__6_, mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_,
         mem_16__1_, mem_16__0_, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N217, N218, N220, N221, N222, N223,
         N224, n6, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29,
         n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57,
         n59, n61, n63, n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2324, n2325, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230;

  DFF_X2 rData1_reg_31_ ( .D(n7195), .CK(n2238), .Q(rData1[31]) );
  DFF_X2 rData1_reg_30_ ( .D(n7196), .CK(n2238), .Q(rData1[30]) );
  DFF_X2 rData1_reg_29_ ( .D(n7197), .CK(n2238), .Q(rData1[29]) );
  DFF_X2 rData1_reg_28_ ( .D(n7198), .CK(n2238), .Q(rData1[28]) );
  DFF_X2 rData1_reg_27_ ( .D(n7199), .CK(n2238), .Q(rData1[27]) );
  DFF_X2 rData1_reg_26_ ( .D(n7200), .CK(n2238), .Q(rData1[26]) );
  DFF_X2 rData1_reg_25_ ( .D(n7201), .CK(n2238), .Q(rData1[25]) );
  DFF_X2 rData1_reg_24_ ( .D(n7202), .CK(n2238), .Q(rData1[24]) );
  DFF_X2 rData1_reg_23_ ( .D(n7203), .CK(n2238), .Q(rData1[23]) );
  DFF_X2 rData1_reg_22_ ( .D(n7204), .CK(n2238), .Q(rData1[22]) );
  DFF_X2 rData1_reg_21_ ( .D(n7205), .CK(n2238), .Q(rData1[21]) );
  DFF_X2 rData1_reg_20_ ( .D(n7206), .CK(n2238), .Q(rData1[20]) );
  DFF_X2 rData1_reg_19_ ( .D(n7207), .CK(n2238), .Q(rData1[19]) );
  DFF_X2 rData1_reg_18_ ( .D(n7208), .CK(n2238), .Q(rData1[18]) );
  DFF_X2 rData1_reg_17_ ( .D(n7209), .CK(n2238), .Q(rData1[17]) );
  DFF_X2 rData1_reg_16_ ( .D(n7210), .CK(n2238), .Q(rData1[16]) );
  DFF_X2 rData1_reg_15_ ( .D(n7211), .CK(n2238), .Q(rData1[15]) );
  DFF_X2 rData1_reg_14_ ( .D(n7212), .CK(n2238), .Q(rData1[14]) );
  DFF_X2 rData1_reg_13_ ( .D(n7213), .CK(n2238), .Q(rData1[13]) );
  DFF_X2 rData1_reg_12_ ( .D(n7214), .CK(n2238), .Q(rData1[12]) );
  DFF_X2 rData1_reg_11_ ( .D(n7215), .CK(n2238), .Q(rData1[11]) );
  DFF_X2 rData1_reg_10_ ( .D(n7216), .CK(n2238), .Q(rData1[10]) );
  DFF_X2 rData1_reg_9_ ( .D(n7217), .CK(n2238), .Q(rData1[9]) );
  DFF_X2 rData1_reg_8_ ( .D(n7218), .CK(n2238), .Q(rData1[8]) );
  DFF_X2 rData1_reg_7_ ( .D(n7219), .CK(n2238), .Q(rData1[7]) );
  DFF_X2 rData1_reg_6_ ( .D(n7220), .CK(n2238), .Q(rData1[6]) );
  DFF_X2 rData1_reg_5_ ( .D(n7221), .CK(n2238), .Q(rData1[5]) );
  DFF_X2 rData1_reg_4_ ( .D(n7222), .CK(n2238), .Q(rData1[4]) );
  DFF_X2 rData1_reg_3_ ( .D(n7223), .CK(n2238), .Q(rData1[3]) );
  DFF_X2 rData1_reg_2_ ( .D(n7224), .CK(n2238), .Q(rData1[2]) );
  DFF_X2 rData1_reg_1_ ( .D(n7225), .CK(n2238), .Q(rData1[1]) );
  DFF_X2 rData1_reg_0_ ( .D(n7226), .CK(n2238), .Q(rData1[0]) );
  DFF_X2 rData2_reg_31_ ( .D(N224), .CK(n2238), .Q(rData2[31]) );
  DFF_X2 rData2_reg_30_ ( .D(N223), .CK(n2238), .Q(rData2[30]) );
  DFF_X2 rData2_reg_29_ ( .D(N222), .CK(n2238), .Q(rData2[29]) );
  DFF_X2 rData2_reg_28_ ( .D(N221), .CK(n2238), .Q(rData2[28]) );
  DFF_X2 rData2_reg_25_ ( .D(N218), .CK(n2238), .Q(rData2[25]) );
  DFF_X2 rData2_reg_22_ ( .D(N215), .CK(n2238), .Q(rData2[22]) );
  DFF_X2 rData2_reg_21_ ( .D(N214), .CK(n2238), .Q(rData2[21]) );
  DFF_X2 rData2_reg_20_ ( .D(N213), .CK(n2238), .Q(rData2[20]) );
  DFF_X2 rData2_reg_19_ ( .D(N212), .CK(n2238), .Q(rData2[19]) );
  DFF_X2 rData2_reg_18_ ( .D(N211), .CK(n2238), .Q(rData2[18]) );
  DFF_X2 rData2_reg_17_ ( .D(N210), .CK(n2238), .Q(rData2[17]) );
  DFF_X2 rData2_reg_16_ ( .D(N209), .CK(n2238), .Q(rData2[16]) );
  DFF_X2 rData2_reg_15_ ( .D(N208), .CK(n2238), .Q(rData2[15]) );
  DFF_X2 rData2_reg_14_ ( .D(N207), .CK(n2238), .Q(rData2[14]) );
  DFF_X2 rData2_reg_13_ ( .D(N206), .CK(n2238), .Q(rData2[13]) );
  DFF_X2 rData2_reg_12_ ( .D(N205), .CK(n2238), .Q(rData2[12]) );
  DFF_X2 rData2_reg_11_ ( .D(N204), .CK(n2238), .Q(rData2[11]) );
  DFF_X2 rData2_reg_10_ ( .D(N203), .CK(n2238), .Q(rData2[10]) );
  DFF_X2 rData2_reg_9_ ( .D(N202), .CK(n2238), .Q(rData2[9]) );
  DFF_X2 rData2_reg_8_ ( .D(N201), .CK(n2238), .Q(rData2[8]) );
  DFF_X2 rData2_reg_7_ ( .D(N200), .CK(n2238), .Q(rData2[7]) );
  DFF_X2 rData2_reg_6_ ( .D(N199), .CK(n2238), .Q(rData2[6]) );
  DFF_X2 rData2_reg_5_ ( .D(N198), .CK(n2238), .Q(rData2[5]) );
  DFF_X2 rData2_reg_4_ ( .D(N197), .CK(n2238), .Q(rData2[4]) );
  DFF_X2 rData2_reg_3_ ( .D(N196), .CK(n2238), .Q(rData2[3]) );
  DFF_X2 rData2_reg_2_ ( .D(N195), .CK(n2238), .Q(rData2[2]) );
  DFF_X2 rData2_reg_1_ ( .D(N194), .CK(n2238), .Q(rData2[1]) );
  DFF_X2 rData2_reg_0_ ( .D(N193), .CK(n2238), .Q(rData2[0]) );
  DFF_X2 mem_reg_31__31_ ( .D(n2173), .CK(clk), .Q(mem_31__31_), .QN(n2746) );
  DFF_X2 mem_reg_31__30_ ( .D(n2172), .CK(clk), .Q(mem_31__30_), .QN(n2744) );
  DFF_X2 mem_reg_31__29_ ( .D(n2171), .CK(clk), .Q(mem_31__29_), .QN(n2742) );
  DFF_X2 mem_reg_31__28_ ( .D(n2170), .CK(clk), .Q(mem_31__28_), .QN(n2634) );
  DFF_X2 mem_reg_31__27_ ( .D(n2169), .CK(clk), .Q(mem_31__27_), .QN(n2658) );
  DFF_X2 mem_reg_31__26_ ( .D(n2168), .CK(clk), .Q(mem_31__26_), .QN(n2630) );
  DFF_X2 mem_reg_31__25_ ( .D(n2167), .CK(clk), .Q(mem_31__25_), .QN(n2636) );
  DFF_X2 mem_reg_31__24_ ( .D(n2166), .CK(clk), .Q(mem_31__24_), .QN(n2660) );
  DFF_X2 mem_reg_31__23_ ( .D(n2165), .CK(clk), .Q(mem_31__23_), .QN(n2652) );
  DFF_X2 mem_reg_31__22_ ( .D(n2164), .CK(clk), .Q(mem_31__22_) );
  DFF_X2 mem_reg_31__21_ ( .D(n2163), .CK(clk), .Q(mem_31__21_) );
  DFF_X2 mem_reg_31__20_ ( .D(n2162), .CK(clk), .Q(mem_31__20_) );
  DFF_X2 mem_reg_31__19_ ( .D(n2161), .CK(clk), .Q(mem_31__19_) );
  DFF_X2 mem_reg_31__18_ ( .D(n2160), .CK(clk), .Q(mem_31__18_) );
  DFF_X2 mem_reg_31__17_ ( .D(n2159), .CK(clk), .Q(mem_31__17_) );
  DFF_X2 mem_reg_31__16_ ( .D(n2158), .CK(clk), .Q(mem_31__16_) );
  DFF_X2 mem_reg_31__15_ ( .D(n2157), .CK(clk), .Q(mem_31__15_) );
  DFF_X2 mem_reg_31__14_ ( .D(n2156), .CK(clk), .Q(mem_31__14_) );
  DFF_X2 mem_reg_31__13_ ( .D(n2155), .CK(clk), .Q(mem_31__13_) );
  DFF_X2 mem_reg_31__12_ ( .D(n2154), .CK(clk), .Q(mem_31__12_) );
  DFF_X2 mem_reg_31__11_ ( .D(n2153), .CK(clk), .Q(mem_31__11_) );
  DFF_X2 mem_reg_31__10_ ( .D(n2152), .CK(clk), .Q(mem_31__10_) );
  DFF_X2 mem_reg_31__9_ ( .D(n2151), .CK(clk), .Q(mem_31__9_) );
  DFF_X2 mem_reg_31__8_ ( .D(n2150), .CK(clk), .Q(mem_31__8_) );
  DFF_X2 mem_reg_31__7_ ( .D(n2149), .CK(clk), .Q(mem_31__7_) );
  DFF_X2 mem_reg_31__6_ ( .D(n2148), .CK(clk), .Q(mem_31__6_) );
  DFF_X2 mem_reg_31__5_ ( .D(n2147), .CK(clk), .Q(mem_31__5_) );
  DFF_X2 mem_reg_31__4_ ( .D(n2146), .CK(clk), .Q(mem_31__4_) );
  DFF_X2 mem_reg_31__3_ ( .D(n2145), .CK(clk), .Q(mem_31__3_) );
  DFF_X2 mem_reg_31__2_ ( .D(n2144), .CK(clk), .Q(mem_31__2_) );
  DFF_X2 mem_reg_31__1_ ( .D(n2143), .CK(clk), .Q(mem_31__1_) );
  DFF_X2 mem_reg_31__0_ ( .D(n2142), .CK(clk), .Q(mem_31__0_) );
  DFF_X2 mem_reg_30__31_ ( .D(n2141), .CK(clk), .Q(mem_30__31_), .QN(n2712) );
  DFF_X2 mem_reg_30__30_ ( .D(n2140), .CK(clk), .Q(mem_30__30_), .QN(n2710) );
  DFF_X2 mem_reg_30__29_ ( .D(n2139), .CK(clk), .Q(mem_30__29_), .QN(n2708) );
  DFF_X2 mem_reg_30__28_ ( .D(n2138), .CK(clk), .Q(mem_30__28_), .QN(n2718) );
  DFF_X2 mem_reg_30__27_ ( .D(n2137), .CK(clk), .Q(mem_30__27_), .QN(n2664) );
  DFF_X2 mem_reg_30__26_ ( .D(n2136), .CK(clk), .Q(mem_30__26_) );
  DFF_X2 mem_reg_30__25_ ( .D(n2135), .CK(clk), .Q(mem_30__25_), .QN(n2720) );
  DFF_X2 mem_reg_30__24_ ( .D(n2134), .CK(clk), .Q(mem_30__24_), .QN(n2666) );
  DFF_X2 mem_reg_30__23_ ( .D(n2133), .CK(clk), .Q(mem_30__23_), .QN(n2730) );
  DFF_X2 mem_reg_30__22_ ( .D(n2132), .CK(clk), .Q(mem_30__22_) );
  DFF_X2 mem_reg_30__21_ ( .D(n2131), .CK(clk), .Q(mem_30__21_) );
  DFF_X2 mem_reg_30__20_ ( .D(n2130), .CK(clk), .Q(mem_30__20_) );
  DFF_X2 mem_reg_30__19_ ( .D(n2129), .CK(clk), .Q(mem_30__19_) );
  DFF_X2 mem_reg_30__18_ ( .D(n2128), .CK(clk), .Q(mem_30__18_) );
  DFF_X2 mem_reg_30__17_ ( .D(n2127), .CK(clk), .Q(mem_30__17_) );
  DFF_X2 mem_reg_30__16_ ( .D(n2126), .CK(clk), .Q(mem_30__16_) );
  DFF_X2 mem_reg_30__15_ ( .D(n2125), .CK(clk), .Q(mem_30__15_) );
  DFF_X2 mem_reg_30__14_ ( .D(n2124), .CK(clk), .Q(mem_30__14_) );
  DFF_X2 mem_reg_30__13_ ( .D(n2123), .CK(clk), .Q(mem_30__13_) );
  DFF_X2 mem_reg_30__12_ ( .D(n2122), .CK(clk), .Q(mem_30__12_) );
  DFF_X2 mem_reg_30__11_ ( .D(n2121), .CK(clk), .Q(mem_30__11_) );
  DFF_X2 mem_reg_30__10_ ( .D(n2120), .CK(clk), .Q(mem_30__10_) );
  DFF_X2 mem_reg_30__9_ ( .D(n2119), .CK(clk), .Q(mem_30__9_) );
  DFF_X2 mem_reg_30__8_ ( .D(n2118), .CK(clk), .Q(mem_30__8_) );
  DFF_X2 mem_reg_30__7_ ( .D(n2117), .CK(clk), .Q(mem_30__7_) );
  DFF_X2 mem_reg_30__6_ ( .D(n2116), .CK(clk), .Q(mem_30__6_) );
  DFF_X2 mem_reg_30__5_ ( .D(n2115), .CK(clk), .Q(mem_30__5_) );
  DFF_X2 mem_reg_30__4_ ( .D(n2114), .CK(clk), .Q(mem_30__4_) );
  DFF_X2 mem_reg_30__3_ ( .D(n2113), .CK(clk), .Q(mem_30__3_) );
  DFF_X2 mem_reg_30__2_ ( .D(n2112), .CK(clk), .Q(mem_30__2_) );
  DFF_X2 mem_reg_30__1_ ( .D(n2111), .CK(clk), .Q(mem_30__1_) );
  DFF_X2 mem_reg_30__0_ ( .D(n2110), .CK(clk), .Q(mem_30__0_) );
  DFF_X2 mem_reg_29__31_ ( .D(n2109), .CK(clk), .Q(mem_29__31_), .QN(n2680) );
  DFF_X2 mem_reg_29__30_ ( .D(n2108), .CK(clk), .Q(mem_29__30_), .QN(n2682) );
  DFF_X2 mem_reg_29__29_ ( .D(n2107), .CK(clk), .Q(mem_29__29_), .QN(n2678) );
  DFF_X2 mem_reg_29__28_ ( .D(n2106), .CK(clk), .Q(mem_29__28_), .QN(n2686) );
  DFF_X2 mem_reg_29__27_ ( .D(n2105), .CK(clk), .Q(mem_29__27_), .QN(n2648) );
  DFF_X2 mem_reg_29__26_ ( .D(n2104), .CK(clk), .Q(mem_29__26_) );
  DFF_X2 mem_reg_29__25_ ( .D(n2103), .CK(clk), .Q(mem_29__25_), .QN(n2688) );
  DFF_X2 mem_reg_29__24_ ( .D(n2102), .CK(clk), .Q(mem_29__24_), .QN(n2650) );
  DFF_X2 mem_reg_29__23_ ( .D(n2101), .CK(clk), .Q(mem_29__23_), .QN(n2714) );
  DFF_X2 mem_reg_29__22_ ( .D(n2100), .CK(clk), .Q(mem_29__22_) );
  DFF_X2 mem_reg_29__21_ ( .D(n2099), .CK(clk), .Q(mem_29__21_) );
  DFF_X2 mem_reg_29__20_ ( .D(n2098), .CK(clk), .Q(mem_29__20_) );
  DFF_X2 mem_reg_29__19_ ( .D(n2097), .CK(clk), .Q(mem_29__19_) );
  DFF_X2 mem_reg_29__18_ ( .D(n2096), .CK(clk), .Q(mem_29__18_) );
  DFF_X2 mem_reg_29__17_ ( .D(n2095), .CK(clk), .Q(mem_29__17_) );
  DFF_X2 mem_reg_29__16_ ( .D(n2094), .CK(clk), .Q(mem_29__16_) );
  DFF_X2 mem_reg_29__15_ ( .D(n2093), .CK(clk), .Q(mem_29__15_) );
  DFF_X2 mem_reg_29__14_ ( .D(n2092), .CK(clk), .Q(mem_29__14_) );
  DFF_X2 mem_reg_29__13_ ( .D(n2091), .CK(clk), .Q(mem_29__13_) );
  DFF_X2 mem_reg_29__12_ ( .D(n2090), .CK(clk), .Q(mem_29__12_) );
  DFF_X2 mem_reg_29__11_ ( .D(n2089), .CK(clk), .Q(mem_29__11_) );
  DFF_X2 mem_reg_29__10_ ( .D(n2088), .CK(clk), .Q(mem_29__10_) );
  DFF_X2 mem_reg_29__9_ ( .D(n2087), .CK(clk), .Q(mem_29__9_) );
  DFF_X2 mem_reg_29__8_ ( .D(n2086), .CK(clk), .Q(mem_29__8_) );
  DFF_X2 mem_reg_29__7_ ( .D(n2085), .CK(clk), .Q(mem_29__7_) );
  DFF_X2 mem_reg_29__6_ ( .D(n2084), .CK(clk), .Q(mem_29__6_) );
  DFF_X2 mem_reg_29__5_ ( .D(n2083), .CK(clk), .Q(mem_29__5_) );
  DFF_X2 mem_reg_29__4_ ( .D(n2082), .CK(clk), .Q(mem_29__4_) );
  DFF_X2 mem_reg_29__3_ ( .D(n2081), .CK(clk), .Q(mem_29__3_) );
  DFF_X2 mem_reg_29__2_ ( .D(n2080), .CK(clk), .Q(mem_29__2_) );
  DFF_X2 mem_reg_29__1_ ( .D(n2079), .CK(clk), .Q(mem_29__1_) );
  DFF_X2 mem_reg_29__0_ ( .D(n2078), .CK(clk), .Q(mem_29__0_) );
  DFF_X2 mem_reg_28__31_ ( .D(n2077), .CK(clk), .Q(mem_28__31_), .QN(n2700) );
  DFF_X2 mem_reg_28__30_ ( .D(n2076), .CK(clk), .Q(mem_28__30_), .QN(n2698) );
  DFF_X2 mem_reg_28__29_ ( .D(n2075), .CK(clk), .Q(mem_28__29_), .QN(n2672) );
  DFF_X2 mem_reg_28__28_ ( .D(n2074), .CK(clk), .Q(mem_28__28_), .QN(n2668) );
  DFF_X2 mem_reg_28__27_ ( .D(n2073), .CK(clk), .Q(mem_28__27_), .QN(n2692) );
  DFF_X2 mem_reg_28__26_ ( .D(n2072), .CK(clk), .Q(mem_28__26_) );
  DFF_X2 mem_reg_28__25_ ( .D(n2071), .CK(clk), .Q(mem_28__25_), .QN(n2670) );
  DFF_X2 mem_reg_28__24_ ( .D(n2070), .CK(clk), .Q(mem_28__24_), .QN(n2694) );
  DFF_X2 mem_reg_28__23_ ( .D(n2069), .CK(clk), .Q(mem_28__23_), .QN(n2696) );
  DFF_X2 mem_reg_28__22_ ( .D(n2068), .CK(clk), .Q(mem_28__22_) );
  DFF_X2 mem_reg_28__21_ ( .D(n2067), .CK(clk), .Q(mem_28__21_) );
  DFF_X2 mem_reg_28__20_ ( .D(n2066), .CK(clk), .Q(mem_28__20_) );
  DFF_X2 mem_reg_28__19_ ( .D(n2065), .CK(clk), .Q(mem_28__19_) );
  DFF_X2 mem_reg_28__18_ ( .D(n2064), .CK(clk), .Q(mem_28__18_) );
  DFF_X2 mem_reg_28__17_ ( .D(n2063), .CK(clk), .Q(mem_28__17_) );
  DFF_X2 mem_reg_28__16_ ( .D(n2062), .CK(clk), .Q(mem_28__16_) );
  DFF_X2 mem_reg_28__15_ ( .D(n2061), .CK(clk), .Q(mem_28__15_) );
  DFF_X2 mem_reg_28__14_ ( .D(n2060), .CK(clk), .Q(mem_28__14_) );
  DFF_X2 mem_reg_28__13_ ( .D(n2059), .CK(clk), .Q(mem_28__13_) );
  DFF_X2 mem_reg_28__12_ ( .D(n2058), .CK(clk), .Q(mem_28__12_) );
  DFF_X2 mem_reg_28__11_ ( .D(n2057), .CK(clk), .Q(mem_28__11_) );
  DFF_X2 mem_reg_28__10_ ( .D(n2056), .CK(clk), .Q(mem_28__10_) );
  DFF_X2 mem_reg_28__9_ ( .D(n2055), .CK(clk), .Q(mem_28__9_) );
  DFF_X2 mem_reg_28__8_ ( .D(n2054), .CK(clk), .Q(mem_28__8_) );
  DFF_X2 mem_reg_28__7_ ( .D(n2053), .CK(clk), .Q(mem_28__7_) );
  DFF_X2 mem_reg_28__6_ ( .D(n2052), .CK(clk), .Q(mem_28__6_) );
  DFF_X2 mem_reg_28__5_ ( .D(n2051), .CK(clk), .Q(mem_28__5_) );
  DFF_X2 mem_reg_28__4_ ( .D(n2050), .CK(clk), .Q(mem_28__4_) );
  DFF_X2 mem_reg_28__3_ ( .D(n2049), .CK(clk), .Q(mem_28__3_) );
  DFF_X2 mem_reg_28__2_ ( .D(n2048), .CK(clk), .Q(mem_28__2_) );
  DFF_X2 mem_reg_28__1_ ( .D(n2047), .CK(clk), .Q(mem_28__1_) );
  DFF_X2 mem_reg_28__0_ ( .D(n2046), .CK(clk), .Q(mem_28__0_) );
  DFF_X2 mem_reg_27__31_ ( .D(n2045), .CK(clk), .Q(mem_27__31_), .QN(n2728) );
  DFF_X2 mem_reg_27__30_ ( .D(n2044), .CK(clk), .Q(mem_27__30_), .QN(n2726) );
  DFF_X2 mem_reg_27__29_ ( .D(n2043), .CK(clk), .Q(mem_27__29_), .QN(n2706) );
  DFF_X2 mem_reg_27__28_ ( .D(n2042), .CK(clk), .Q(mem_27__28_), .QN(n2702) );
  DFF_X2 mem_reg_27__27_ ( .D(n2041), .CK(clk), .Q(mem_27__27_), .QN(n2722) );
  DFF_X2 mem_reg_27__26_ ( .D(n2040), .CK(clk), .Q(mem_27__26_), .QN(n2632) );
  DFF_X2 mem_reg_27__25_ ( .D(n2039), .CK(clk), .Q(mem_27__25_), .QN(n2704) );
  DFF_X2 mem_reg_27__24_ ( .D(n2038), .CK(clk), .Q(mem_27__24_), .QN(n2724) );
  DFF_X2 mem_reg_27__23_ ( .D(n2037), .CK(clk), .Q(mem_27__23_), .QN(n2716) );
  DFF_X2 mem_reg_27__22_ ( .D(n2036), .CK(clk), .Q(mem_27__22_) );
  DFF_X2 mem_reg_27__21_ ( .D(n2035), .CK(clk), .Q(mem_27__21_) );
  DFF_X2 mem_reg_27__20_ ( .D(n2034), .CK(clk), .Q(mem_27__20_) );
  DFF_X2 mem_reg_27__19_ ( .D(n2033), .CK(clk), .Q(mem_27__19_) );
  DFF_X2 mem_reg_27__18_ ( .D(n2032), .CK(clk), .Q(mem_27__18_) );
  DFF_X2 mem_reg_27__17_ ( .D(n2031), .CK(clk), .Q(mem_27__17_) );
  DFF_X2 mem_reg_27__16_ ( .D(n2030), .CK(clk), .Q(mem_27__16_) );
  DFF_X2 mem_reg_27__15_ ( .D(n2029), .CK(clk), .Q(mem_27__15_) );
  DFF_X2 mem_reg_27__14_ ( .D(n2028), .CK(clk), .Q(mem_27__14_) );
  DFF_X2 mem_reg_27__13_ ( .D(n2027), .CK(clk), .Q(mem_27__13_) );
  DFF_X2 mem_reg_27__12_ ( .D(n2026), .CK(clk), .Q(mem_27__12_) );
  DFF_X2 mem_reg_27__11_ ( .D(n2025), .CK(clk), .Q(mem_27__11_) );
  DFF_X2 mem_reg_27__10_ ( .D(n2024), .CK(clk), .Q(mem_27__10_) );
  DFF_X2 mem_reg_27__9_ ( .D(n2023), .CK(clk), .Q(mem_27__9_) );
  DFF_X2 mem_reg_27__8_ ( .D(n2022), .CK(clk), .Q(mem_27__8_) );
  DFF_X2 mem_reg_27__7_ ( .D(n2021), .CK(clk), .Q(mem_27__7_) );
  DFF_X2 mem_reg_27__6_ ( .D(n2020), .CK(clk), .Q(mem_27__6_) );
  DFF_X2 mem_reg_27__5_ ( .D(n2019), .CK(clk), .Q(mem_27__5_) );
  DFF_X2 mem_reg_27__4_ ( .D(n2018), .CK(clk), .Q(mem_27__4_) );
  DFF_X2 mem_reg_27__3_ ( .D(n2017), .CK(clk), .Q(mem_27__3_) );
  DFF_X2 mem_reg_27__2_ ( .D(n2016), .CK(clk), .Q(mem_27__2_) );
  DFF_X2 mem_reg_27__1_ ( .D(n2015), .CK(clk), .Q(mem_27__1_) );
  DFF_X2 mem_reg_27__0_ ( .D(n2014), .CK(clk), .Q(mem_27__0_) );
  DFF_X2 mem_reg_26__31_ ( .D(n2013), .CK(clk), .Q(mem_26__31_), .QN(n2676) );
  DFF_X2 mem_reg_26__30_ ( .D(n2012), .CK(clk), .Q(mem_26__30_), .QN(n2748) );
  DFF_X2 mem_reg_26__29_ ( .D(n2011), .CK(clk), .Q(mem_26__29_), .QN(n2740) );
  DFF_X2 mem_reg_26__28_ ( .D(n2010), .CK(clk), .Q(mem_26__28_), .QN(n2734) );
  DFF_X2 mem_reg_26__27_ ( .D(n2009), .CK(clk), .Q(mem_26__27_), .QN(n2732) );
  DFF_X2 mem_reg_26__26_ ( .D(n2008), .CK(clk), .Q(mem_26__26_), .QN(n2644) );
  DFF_X2 mem_reg_26__25_ ( .D(n2007), .CK(clk), .Q(mem_26__25_), .QN(n2738) );
  DFF_X2 mem_reg_26__24_ ( .D(n2006), .CK(clk), .Q(mem_26__24_), .QN(n2662) );
  DFF_X2 mem_reg_26__23_ ( .D(n2005), .CK(clk), .Q(mem_26__23_), .QN(n2684) );
  DFF_X2 mem_reg_26__22_ ( .D(n2004), .CK(clk), .Q(mem_26__22_) );
  DFF_X2 mem_reg_26__21_ ( .D(n2003), .CK(clk), .Q(mem_26__21_) );
  DFF_X2 mem_reg_26__20_ ( .D(n2002), .CK(clk), .Q(mem_26__20_) );
  DFF_X2 mem_reg_26__19_ ( .D(n2001), .CK(clk), .Q(mem_26__19_) );
  DFF_X2 mem_reg_26__18_ ( .D(n2000), .CK(clk), .Q(mem_26__18_) );
  DFF_X2 mem_reg_26__17_ ( .D(n1999), .CK(clk), .Q(mem_26__17_) );
  DFF_X2 mem_reg_26__16_ ( .D(n1998), .CK(clk), .Q(mem_26__16_) );
  DFF_X2 mem_reg_26__15_ ( .D(n1997), .CK(clk), .Q(mem_26__15_) );
  DFF_X2 mem_reg_26__14_ ( .D(n1996), .CK(clk), .Q(mem_26__14_) );
  DFF_X2 mem_reg_26__13_ ( .D(n1995), .CK(clk), .Q(mem_26__13_) );
  DFF_X2 mem_reg_26__12_ ( .D(n1994), .CK(clk), .Q(mem_26__12_) );
  DFF_X2 mem_reg_26__11_ ( .D(n1993), .CK(clk), .Q(mem_26__11_) );
  DFF_X2 mem_reg_26__10_ ( .D(n1992), .CK(clk), .Q(mem_26__10_) );
  DFF_X2 mem_reg_26__9_ ( .D(n1991), .CK(clk), .Q(mem_26__9_) );
  DFF_X2 mem_reg_26__8_ ( .D(n1990), .CK(clk), .Q(mem_26__8_) );
  DFF_X2 mem_reg_26__7_ ( .D(n1989), .CK(clk), .Q(mem_26__7_) );
  DFF_X2 mem_reg_26__6_ ( .D(n1988), .CK(clk), .Q(mem_26__6_) );
  DFF_X2 mem_reg_26__5_ ( .D(n1987), .CK(clk), .Q(mem_26__5_) );
  DFF_X2 mem_reg_26__4_ ( .D(n1986), .CK(clk), .Q(mem_26__4_) );
  DFF_X2 mem_reg_26__3_ ( .D(n1985), .CK(clk), .Q(mem_26__3_) );
  DFF_X2 mem_reg_26__2_ ( .D(n1984), .CK(clk), .Q(mem_26__2_) );
  DFF_X2 mem_reg_26__1_ ( .D(n1983), .CK(clk), .Q(mem_26__1_) );
  DFF_X2 mem_reg_26__0_ ( .D(n1982), .CK(clk), .Q(mem_26__0_) );
  DFF_X2 mem_reg_25__31_ ( .D(n1981), .CK(clk), .Q(mem_25__31_) );
  DFF_X2 mem_reg_25__30_ ( .D(n1980), .CK(clk), .Q(mem_25__30_) );
  DFF_X2 mem_reg_25__29_ ( .D(n1979), .CK(clk), .Q(mem_25__29_) );
  DFF_X2 mem_reg_25__28_ ( .D(n1978), .CK(clk), .Q(mem_25__28_) );
  DFF_X2 mem_reg_25__27_ ( .D(n1977), .CK(clk), .Q(mem_25__27_) );
  DFF_X2 mem_reg_25__26_ ( .D(n1976), .CK(clk), .Q(mem_25__26_) );
  DFF_X2 mem_reg_25__25_ ( .D(n1975), .CK(clk), .Q(mem_25__25_) );
  DFF_X2 mem_reg_25__24_ ( .D(n1974), .CK(clk), .Q(mem_25__24_) );
  DFF_X2 mem_reg_25__23_ ( .D(n1973), .CK(clk), .Q(mem_25__23_) );
  DFF_X2 mem_reg_25__22_ ( .D(n1972), .CK(clk), .Q(mem_25__22_) );
  DFF_X2 mem_reg_25__21_ ( .D(n1971), .CK(clk), .Q(mem_25__21_) );
  DFF_X2 mem_reg_25__20_ ( .D(n1970), .CK(clk), .Q(mem_25__20_) );
  DFF_X2 mem_reg_25__19_ ( .D(n1969), .CK(clk), .Q(mem_25__19_) );
  DFF_X2 mem_reg_25__18_ ( .D(n1968), .CK(clk), .Q(mem_25__18_) );
  DFF_X2 mem_reg_25__17_ ( .D(n1967), .CK(clk), .Q(mem_25__17_) );
  DFF_X2 mem_reg_25__16_ ( .D(n1966), .CK(clk), .Q(mem_25__16_) );
  DFF_X2 mem_reg_25__15_ ( .D(n1965), .CK(clk), .Q(mem_25__15_) );
  DFF_X2 mem_reg_25__14_ ( .D(n1964), .CK(clk), .Q(mem_25__14_) );
  DFF_X2 mem_reg_25__13_ ( .D(n1963), .CK(clk), .Q(mem_25__13_) );
  DFF_X2 mem_reg_25__12_ ( .D(n1962), .CK(clk), .Q(mem_25__12_) );
  DFF_X2 mem_reg_25__11_ ( .D(n1961), .CK(clk), .Q(mem_25__11_) );
  DFF_X2 mem_reg_25__10_ ( .D(n1960), .CK(clk), .Q(mem_25__10_) );
  DFF_X2 mem_reg_25__9_ ( .D(n1959), .CK(clk), .Q(mem_25__9_) );
  DFF_X2 mem_reg_25__8_ ( .D(n1958), .CK(clk), .Q(mem_25__8_) );
  DFF_X2 mem_reg_25__7_ ( .D(n1957), .CK(clk), .Q(mem_25__7_) );
  DFF_X2 mem_reg_25__6_ ( .D(n1956), .CK(clk), .Q(mem_25__6_) );
  DFF_X2 mem_reg_25__5_ ( .D(n1955), .CK(clk), .Q(mem_25__5_) );
  DFF_X2 mem_reg_25__4_ ( .D(n1954), .CK(clk), .Q(mem_25__4_) );
  DFF_X2 mem_reg_25__3_ ( .D(n1953), .CK(clk), .Q(mem_25__3_) );
  DFF_X2 mem_reg_25__2_ ( .D(n1952), .CK(clk), .Q(mem_25__2_) );
  DFF_X2 mem_reg_25__1_ ( .D(n1951), .CK(clk), .Q(mem_25__1_) );
  DFF_X2 mem_reg_25__0_ ( .D(n1950), .CK(clk), .Q(mem_25__0_) );
  DFF_X2 mem_reg_24__31_ ( .D(n1949), .CK(clk), .Q(mem_24__31_) );
  DFF_X2 mem_reg_24__30_ ( .D(n1948), .CK(clk), .Q(mem_24__30_) );
  DFF_X2 mem_reg_24__29_ ( .D(n1947), .CK(clk), .Q(mem_24__29_) );
  DFF_X2 mem_reg_24__28_ ( .D(n1946), .CK(clk), .Q(mem_24__28_) );
  DFF_X2 mem_reg_24__27_ ( .D(n1945), .CK(clk), .Q(mem_24__27_) );
  DFF_X2 mem_reg_24__26_ ( .D(n1944), .CK(clk), .Q(mem_24__26_) );
  DFF_X2 mem_reg_24__25_ ( .D(n1943), .CK(clk), .Q(mem_24__25_) );
  DFF_X2 mem_reg_24__24_ ( .D(n1942), .CK(clk), .Q(mem_24__24_) );
  DFF_X2 mem_reg_24__23_ ( .D(n1941), .CK(clk), .Q(mem_24__23_) );
  DFF_X2 mem_reg_24__22_ ( .D(n1940), .CK(clk), .Q(mem_24__22_) );
  DFF_X2 mem_reg_24__21_ ( .D(n1939), .CK(clk), .Q(mem_24__21_) );
  DFF_X2 mem_reg_24__20_ ( .D(n1938), .CK(clk), .Q(mem_24__20_) );
  DFF_X2 mem_reg_24__19_ ( .D(n1937), .CK(clk), .Q(mem_24__19_) );
  DFF_X2 mem_reg_24__18_ ( .D(n1936), .CK(clk), .Q(mem_24__18_) );
  DFF_X2 mem_reg_24__17_ ( .D(n1935), .CK(clk), .Q(mem_24__17_) );
  DFF_X2 mem_reg_24__16_ ( .D(n1934), .CK(clk), .Q(mem_24__16_) );
  DFF_X2 mem_reg_24__15_ ( .D(n1933), .CK(clk), .Q(mem_24__15_) );
  DFF_X2 mem_reg_24__14_ ( .D(n1932), .CK(clk), .Q(mem_24__14_) );
  DFF_X2 mem_reg_24__13_ ( .D(n1931), .CK(clk), .Q(mem_24__13_) );
  DFF_X2 mem_reg_24__12_ ( .D(n1930), .CK(clk), .Q(mem_24__12_) );
  DFF_X2 mem_reg_24__11_ ( .D(n1929), .CK(clk), .Q(mem_24__11_) );
  DFF_X2 mem_reg_24__10_ ( .D(n1928), .CK(clk), .Q(mem_24__10_) );
  DFF_X2 mem_reg_24__9_ ( .D(n1927), .CK(clk), .Q(mem_24__9_) );
  DFF_X2 mem_reg_24__8_ ( .D(n1926), .CK(clk), .Q(mem_24__8_) );
  DFF_X2 mem_reg_24__7_ ( .D(n1925), .CK(clk), .Q(mem_24__7_) );
  DFF_X2 mem_reg_24__6_ ( .D(n1924), .CK(clk), .Q(mem_24__6_) );
  DFF_X2 mem_reg_24__5_ ( .D(n1923), .CK(clk), .Q(mem_24__5_) );
  DFF_X2 mem_reg_24__4_ ( .D(n1922), .CK(clk), .Q(mem_24__4_) );
  DFF_X2 mem_reg_24__3_ ( .D(n1921), .CK(clk), .Q(mem_24__3_) );
  DFF_X2 mem_reg_24__2_ ( .D(n1920), .CK(clk), .Q(mem_24__2_) );
  DFF_X2 mem_reg_24__1_ ( .D(n1919), .CK(clk), .Q(mem_24__1_) );
  DFF_X2 mem_reg_24__0_ ( .D(n1918), .CK(clk), .Q(mem_24__0_) );
  DFF_X2 mem_reg_23__31_ ( .D(n1917), .CK(clk), .Q(mem_23__31_) );
  DFF_X2 mem_reg_23__30_ ( .D(n1916), .CK(clk), .Q(mem_23__30_) );
  DFF_X2 mem_reg_23__29_ ( .D(n1915), .CK(clk), .Q(mem_23__29_) );
  DFF_X2 mem_reg_23__28_ ( .D(n1914), .CK(clk), .Q(mem_23__28_) );
  DFF_X2 mem_reg_23__27_ ( .D(n1913), .CK(clk), .Q(mem_23__27_) );
  DFF_X2 mem_reg_23__26_ ( .D(n1912), .CK(clk), .Q(mem_23__26_), .QN(n2638) );
  DFF_X2 mem_reg_23__25_ ( .D(n1911), .CK(clk), .Q(mem_23__25_) );
  DFF_X2 mem_reg_23__24_ ( .D(n1910), .CK(clk), .Q(mem_23__24_) );
  DFF_X2 mem_reg_23__23_ ( .D(n1909), .CK(clk), .Q(mem_23__23_) );
  DFF_X2 mem_reg_23__22_ ( .D(n1908), .CK(clk), .Q(mem_23__22_) );
  DFF_X2 mem_reg_23__21_ ( .D(n1907), .CK(clk), .Q(mem_23__21_) );
  DFF_X2 mem_reg_23__20_ ( .D(n1906), .CK(clk), .Q(mem_23__20_) );
  DFF_X2 mem_reg_23__19_ ( .D(n1905), .CK(clk), .Q(mem_23__19_) );
  DFF_X2 mem_reg_23__18_ ( .D(n1904), .CK(clk), .Q(mem_23__18_) );
  DFF_X2 mem_reg_23__17_ ( .D(n1903), .CK(clk), .Q(mem_23__17_) );
  DFF_X2 mem_reg_23__16_ ( .D(n1902), .CK(clk), .Q(mem_23__16_) );
  DFF_X2 mem_reg_23__15_ ( .D(n1901), .CK(clk), .Q(mem_23__15_) );
  DFF_X2 mem_reg_23__14_ ( .D(n1900), .CK(clk), .Q(mem_23__14_) );
  DFF_X2 mem_reg_23__13_ ( .D(n1899), .CK(clk), .Q(mem_23__13_) );
  DFF_X2 mem_reg_23__12_ ( .D(n1898), .CK(clk), .Q(mem_23__12_) );
  DFF_X2 mem_reg_23__11_ ( .D(n1897), .CK(clk), .Q(mem_23__11_) );
  DFF_X2 mem_reg_23__10_ ( .D(n1896), .CK(clk), .Q(mem_23__10_) );
  DFF_X2 mem_reg_23__9_ ( .D(n1895), .CK(clk), .Q(mem_23__9_) );
  DFF_X2 mem_reg_23__8_ ( .D(n1894), .CK(clk), .Q(mem_23__8_) );
  DFF_X2 mem_reg_23__7_ ( .D(n1893), .CK(clk), .Q(mem_23__7_) );
  DFF_X2 mem_reg_23__6_ ( .D(n1892), .CK(clk), .Q(mem_23__6_) );
  DFF_X2 mem_reg_23__5_ ( .D(n1891), .CK(clk), .Q(mem_23__5_) );
  DFF_X2 mem_reg_23__4_ ( .D(n1890), .CK(clk), .Q(mem_23__4_) );
  DFF_X2 mem_reg_23__3_ ( .D(n1889), .CK(clk), .Q(mem_23__3_) );
  DFF_X2 mem_reg_23__2_ ( .D(n1888), .CK(clk), .Q(mem_23__2_) );
  DFF_X2 mem_reg_23__1_ ( .D(n1887), .CK(clk), .Q(mem_23__1_) );
  DFF_X2 mem_reg_23__0_ ( .D(n1886), .CK(clk), .Q(mem_23__0_) );
  DFF_X2 mem_reg_22__31_ ( .D(n1885), .CK(clk), .Q(mem_22__31_) );
  DFF_X2 mem_reg_22__30_ ( .D(n1884), .CK(clk), .Q(mem_22__30_) );
  DFF_X2 mem_reg_22__29_ ( .D(n1883), .CK(clk), .Q(mem_22__29_) );
  DFF_X2 mem_reg_22__28_ ( .D(n1882), .CK(clk), .Q(mem_22__28_) );
  DFF_X2 mem_reg_22__27_ ( .D(n1881), .CK(clk), .Q(mem_22__27_) );
  DFF_X2 mem_reg_22__26_ ( .D(n1880), .CK(clk), .Q(mem_22__26_), .QN(n2656) );
  DFF_X2 mem_reg_22__25_ ( .D(n1879), .CK(clk), .Q(mem_22__25_) );
  DFF_X2 mem_reg_22__24_ ( .D(n1878), .CK(clk), .Q(mem_22__24_) );
  DFF_X2 mem_reg_22__23_ ( .D(n1877), .CK(clk), .Q(mem_22__23_) );
  DFF_X2 mem_reg_22__22_ ( .D(n1876), .CK(clk), .Q(mem_22__22_) );
  DFF_X2 mem_reg_22__21_ ( .D(n1875), .CK(clk), .Q(mem_22__21_) );
  DFF_X2 mem_reg_22__20_ ( .D(n1874), .CK(clk), .Q(mem_22__20_) );
  DFF_X2 mem_reg_22__19_ ( .D(n1873), .CK(clk), .Q(mem_22__19_) );
  DFF_X2 mem_reg_22__18_ ( .D(n1872), .CK(clk), .Q(mem_22__18_) );
  DFF_X2 mem_reg_22__17_ ( .D(n1871), .CK(clk), .Q(mem_22__17_) );
  DFF_X2 mem_reg_22__16_ ( .D(n1870), .CK(clk), .Q(mem_22__16_) );
  DFF_X2 mem_reg_22__15_ ( .D(n1869), .CK(clk), .Q(mem_22__15_) );
  DFF_X2 mem_reg_22__14_ ( .D(n1868), .CK(clk), .Q(mem_22__14_) );
  DFF_X2 mem_reg_22__13_ ( .D(n1867), .CK(clk), .Q(mem_22__13_) );
  DFF_X2 mem_reg_22__12_ ( .D(n1866), .CK(clk), .Q(mem_22__12_) );
  DFF_X2 mem_reg_22__11_ ( .D(n1865), .CK(clk), .Q(mem_22__11_) );
  DFF_X2 mem_reg_22__10_ ( .D(n1864), .CK(clk), .Q(mem_22__10_) );
  DFF_X2 mem_reg_22__9_ ( .D(n1863), .CK(clk), .Q(mem_22__9_) );
  DFF_X2 mem_reg_22__8_ ( .D(n1862), .CK(clk), .Q(mem_22__8_) );
  DFF_X2 mem_reg_22__7_ ( .D(n1861), .CK(clk), .Q(mem_22__7_) );
  DFF_X2 mem_reg_22__6_ ( .D(n1860), .CK(clk), .Q(mem_22__6_) );
  DFF_X2 mem_reg_22__5_ ( .D(n1859), .CK(clk), .Q(mem_22__5_) );
  DFF_X2 mem_reg_22__4_ ( .D(n1858), .CK(clk), .Q(mem_22__4_) );
  DFF_X2 mem_reg_22__3_ ( .D(n1857), .CK(clk), .Q(mem_22__3_) );
  DFF_X2 mem_reg_22__2_ ( .D(n1856), .CK(clk), .Q(mem_22__2_) );
  DFF_X2 mem_reg_22__1_ ( .D(n1855), .CK(clk), .Q(mem_22__1_) );
  DFF_X2 mem_reg_22__0_ ( .D(n1854), .CK(clk), .Q(mem_22__0_) );
  DFF_X2 mem_reg_21__31_ ( .D(n1853), .CK(clk), .Q(mem_21__31_) );
  DFF_X2 mem_reg_21__30_ ( .D(n1852), .CK(clk), .Q(mem_21__30_) );
  DFF_X2 mem_reg_21__29_ ( .D(n1851), .CK(clk), .Q(mem_21__29_) );
  DFF_X2 mem_reg_21__28_ ( .D(n1850), .CK(clk), .Q(mem_21__28_) );
  DFF_X2 mem_reg_21__27_ ( .D(n1849), .CK(clk), .Q(mem_21__27_) );
  DFF_X2 mem_reg_21__26_ ( .D(n1848), .CK(clk), .Q(mem_21__26_), .QN(n2690) );
  DFF_X2 mem_reg_21__25_ ( .D(n1847), .CK(clk), .Q(mem_21__25_) );
  DFF_X2 mem_reg_21__24_ ( .D(n1846), .CK(clk), .Q(mem_21__24_) );
  DFF_X2 mem_reg_21__23_ ( .D(n1845), .CK(clk), .Q(mem_21__23_) );
  DFF_X2 mem_reg_21__22_ ( .D(n1844), .CK(clk), .Q(mem_21__22_) );
  DFF_X2 mem_reg_21__21_ ( .D(n1843), .CK(clk), .Q(mem_21__21_) );
  DFF_X2 mem_reg_21__20_ ( .D(n1842), .CK(clk), .Q(mem_21__20_) );
  DFF_X2 mem_reg_21__19_ ( .D(n1841), .CK(clk), .Q(mem_21__19_) );
  DFF_X2 mem_reg_21__18_ ( .D(n1840), .CK(clk), .Q(mem_21__18_) );
  DFF_X2 mem_reg_21__17_ ( .D(n1839), .CK(clk), .Q(mem_21__17_) );
  DFF_X2 mem_reg_21__16_ ( .D(n1838), .CK(clk), .Q(mem_21__16_) );
  DFF_X2 mem_reg_21__15_ ( .D(n1837), .CK(clk), .Q(mem_21__15_) );
  DFF_X2 mem_reg_21__14_ ( .D(n1836), .CK(clk), .Q(mem_21__14_) );
  DFF_X2 mem_reg_21__13_ ( .D(n1835), .CK(clk), .Q(mem_21__13_) );
  DFF_X2 mem_reg_21__12_ ( .D(n1834), .CK(clk), .Q(mem_21__12_) );
  DFF_X2 mem_reg_21__11_ ( .D(n1833), .CK(clk), .Q(mem_21__11_) );
  DFF_X2 mem_reg_21__10_ ( .D(n1832), .CK(clk), .Q(mem_21__10_) );
  DFF_X2 mem_reg_21__9_ ( .D(n1831), .CK(clk), .Q(mem_21__9_) );
  DFF_X2 mem_reg_21__8_ ( .D(n1830), .CK(clk), .Q(mem_21__8_) );
  DFF_X2 mem_reg_21__7_ ( .D(n1829), .CK(clk), .Q(mem_21__7_) );
  DFF_X2 mem_reg_21__6_ ( .D(n1828), .CK(clk), .Q(mem_21__6_) );
  DFF_X2 mem_reg_21__5_ ( .D(n1827), .CK(clk), .Q(mem_21__5_) );
  DFF_X2 mem_reg_21__4_ ( .D(n1826), .CK(clk), .Q(mem_21__4_) );
  DFF_X2 mem_reg_21__3_ ( .D(n1825), .CK(clk), .Q(mem_21__3_) );
  DFF_X2 mem_reg_21__2_ ( .D(n1824), .CK(clk), .Q(mem_21__2_) );
  DFF_X2 mem_reg_21__1_ ( .D(n1823), .CK(clk), .Q(mem_21__1_) );
  DFF_X2 mem_reg_21__0_ ( .D(n1822), .CK(clk), .Q(mem_21__0_) );
  DFF_X2 mem_reg_20__31_ ( .D(n1821), .CK(clk), .Q(mem_20__31_) );
  DFF_X2 mem_reg_20__30_ ( .D(n1820), .CK(clk), .Q(mem_20__30_) );
  DFF_X2 mem_reg_20__29_ ( .D(n1819), .CK(clk), .Q(mem_20__29_) );
  DFF_X2 mem_reg_20__28_ ( .D(n1818), .CK(clk), .Q(mem_20__28_) );
  DFF_X2 mem_reg_20__27_ ( .D(n1817), .CK(clk), .Q(mem_20__27_) );
  DFF_X2 mem_reg_20__26_ ( .D(n1816), .CK(clk), .Q(mem_20__26_), .QN(n2674) );
  DFF_X2 mem_reg_20__25_ ( .D(n1815), .CK(clk), .Q(mem_20__25_) );
  DFF_X2 mem_reg_20__24_ ( .D(n1814), .CK(clk), .Q(mem_20__24_) );
  DFF_X2 mem_reg_20__23_ ( .D(n1813), .CK(clk), .Q(mem_20__23_) );
  DFF_X2 mem_reg_20__22_ ( .D(n1812), .CK(clk), .Q(mem_20__22_) );
  DFF_X2 mem_reg_20__21_ ( .D(n1811), .CK(clk), .Q(mem_20__21_) );
  DFF_X2 mem_reg_20__20_ ( .D(n1810), .CK(clk), .Q(mem_20__20_) );
  DFF_X2 mem_reg_20__19_ ( .D(n1809), .CK(clk), .Q(mem_20__19_) );
  DFF_X2 mem_reg_20__18_ ( .D(n1808), .CK(clk), .Q(mem_20__18_) );
  DFF_X2 mem_reg_20__17_ ( .D(n1807), .CK(clk), .Q(mem_20__17_) );
  DFF_X2 mem_reg_20__16_ ( .D(n1806), .CK(clk), .Q(mem_20__16_) );
  DFF_X2 mem_reg_20__15_ ( .D(n1805), .CK(clk), .Q(mem_20__15_) );
  DFF_X2 mem_reg_20__14_ ( .D(n1804), .CK(clk), .Q(mem_20__14_) );
  DFF_X2 mem_reg_20__13_ ( .D(n1803), .CK(clk), .Q(mem_20__13_) );
  DFF_X2 mem_reg_20__12_ ( .D(n1802), .CK(clk), .Q(mem_20__12_) );
  DFF_X2 mem_reg_20__11_ ( .D(n1801), .CK(clk), .Q(mem_20__11_) );
  DFF_X2 mem_reg_20__10_ ( .D(n1800), .CK(clk), .Q(mem_20__10_) );
  DFF_X2 mem_reg_20__9_ ( .D(n1799), .CK(clk), .Q(mem_20__9_) );
  DFF_X2 mem_reg_20__8_ ( .D(n1798), .CK(clk), .Q(mem_20__8_) );
  DFF_X2 mem_reg_20__7_ ( .D(n1797), .CK(clk), .Q(mem_20__7_) );
  DFF_X2 mem_reg_20__6_ ( .D(n1796), .CK(clk), .Q(mem_20__6_) );
  DFF_X2 mem_reg_20__5_ ( .D(n1795), .CK(clk), .Q(mem_20__5_) );
  DFF_X2 mem_reg_20__4_ ( .D(n1794), .CK(clk), .Q(mem_20__4_) );
  DFF_X2 mem_reg_20__3_ ( .D(n1793), .CK(clk), .Q(mem_20__3_) );
  DFF_X2 mem_reg_20__2_ ( .D(n1792), .CK(clk), .Q(mem_20__2_) );
  DFF_X2 mem_reg_20__1_ ( .D(n1791), .CK(clk), .Q(mem_20__1_) );
  DFF_X2 mem_reg_20__0_ ( .D(n1790), .CK(clk), .Q(mem_20__0_) );
  DFF_X2 mem_reg_19__31_ ( .D(n1789), .CK(clk), .Q(mem_19__31_) );
  DFF_X2 mem_reg_19__30_ ( .D(n1788), .CK(clk), .Q(mem_19__30_) );
  DFF_X2 mem_reg_19__29_ ( .D(n1787), .CK(clk), .Q(mem_19__29_) );
  DFF_X2 mem_reg_19__28_ ( .D(n1786), .CK(clk), .Q(mem_19__28_) );
  DFF_X2 mem_reg_19__27_ ( .D(n1785), .CK(clk), .Q(mem_19__27_) );
  DFF_X2 mem_reg_19__26_ ( .D(n1784), .CK(clk), .Q(mem_19__26_), .QN(n2654) );
  DFF_X2 mem_reg_19__25_ ( .D(n1783), .CK(clk), .Q(mem_19__25_) );
  DFF_X2 mem_reg_19__24_ ( .D(n1782), .CK(clk), .Q(mem_19__24_) );
  DFF_X2 mem_reg_19__23_ ( .D(n1781), .CK(clk), .Q(mem_19__23_) );
  DFF_X2 mem_reg_19__22_ ( .D(n1780), .CK(clk), .Q(mem_19__22_) );
  DFF_X2 mem_reg_19__21_ ( .D(n1779), .CK(clk), .Q(mem_19__21_) );
  DFF_X2 mem_reg_19__20_ ( .D(n1778), .CK(clk), .Q(mem_19__20_) );
  DFF_X2 mem_reg_19__19_ ( .D(n1777), .CK(clk), .Q(mem_19__19_) );
  DFF_X2 mem_reg_19__18_ ( .D(n1776), .CK(clk), .Q(mem_19__18_) );
  DFF_X2 mem_reg_19__17_ ( .D(n1775), .CK(clk), .Q(mem_19__17_) );
  DFF_X2 mem_reg_19__16_ ( .D(n1774), .CK(clk), .Q(mem_19__16_) );
  DFF_X2 mem_reg_19__15_ ( .D(n1773), .CK(clk), .Q(mem_19__15_) );
  DFF_X2 mem_reg_19__14_ ( .D(n1772), .CK(clk), .Q(mem_19__14_) );
  DFF_X2 mem_reg_19__13_ ( .D(n1771), .CK(clk), .Q(mem_19__13_) );
  DFF_X2 mem_reg_19__12_ ( .D(n1770), .CK(clk), .Q(mem_19__12_) );
  DFF_X2 mem_reg_19__11_ ( .D(n1769), .CK(clk), .Q(mem_19__11_) );
  DFF_X2 mem_reg_19__10_ ( .D(n1768), .CK(clk), .Q(mem_19__10_) );
  DFF_X2 mem_reg_19__9_ ( .D(n1767), .CK(clk), .Q(mem_19__9_) );
  DFF_X2 mem_reg_19__8_ ( .D(n1766), .CK(clk), .Q(mem_19__8_) );
  DFF_X2 mem_reg_19__7_ ( .D(n1765), .CK(clk), .Q(mem_19__7_) );
  DFF_X2 mem_reg_19__6_ ( .D(n1764), .CK(clk), .Q(mem_19__6_) );
  DFF_X2 mem_reg_19__5_ ( .D(n1763), .CK(clk), .Q(mem_19__5_) );
  DFF_X2 mem_reg_19__4_ ( .D(n1762), .CK(clk), .Q(mem_19__4_) );
  DFF_X2 mem_reg_19__3_ ( .D(n1761), .CK(clk), .Q(mem_19__3_) );
  DFF_X2 mem_reg_19__2_ ( .D(n1760), .CK(clk), .Q(mem_19__2_) );
  DFF_X2 mem_reg_19__1_ ( .D(n1759), .CK(clk), .Q(mem_19__1_) );
  DFF_X2 mem_reg_19__0_ ( .D(n1758), .CK(clk), .Q(mem_19__0_) );
  DFF_X2 mem_reg_18__31_ ( .D(n1757), .CK(clk), .Q(mem_18__31_) );
  DFF_X2 mem_reg_18__30_ ( .D(n1756), .CK(clk), .Q(mem_18__30_) );
  DFF_X2 mem_reg_18__29_ ( .D(n1755), .CK(clk), .Q(mem_18__29_), .QN(n2640) );
  DFF_X2 mem_reg_18__28_ ( .D(n1754), .CK(clk), .Q(mem_18__28_), .QN(n2642) );
  DFF_X2 mem_reg_18__27_ ( .D(n1753), .CK(clk), .Q(mem_18__27_) );
  DFF_X2 mem_reg_18__26_ ( .D(n1752), .CK(clk), .Q(mem_18__26_), .QN(n2736) );
  DFF_X2 mem_reg_18__25_ ( .D(n1751), .CK(clk), .Q(mem_18__25_), .QN(n2646) );
  DFF_X2 mem_reg_18__24_ ( .D(n1750), .CK(clk), .Q(mem_18__24_) );
  DFF_X2 mem_reg_18__23_ ( .D(n1749), .CK(clk), .Q(mem_18__23_) );
  DFF_X2 mem_reg_18__22_ ( .D(n1748), .CK(clk), .Q(mem_18__22_) );
  DFF_X2 mem_reg_18__21_ ( .D(n1747), .CK(clk), .Q(mem_18__21_) );
  DFF_X2 mem_reg_18__20_ ( .D(n1746), .CK(clk), .Q(mem_18__20_) );
  DFF_X2 mem_reg_18__19_ ( .D(n1745), .CK(clk), .Q(mem_18__19_) );
  DFF_X2 mem_reg_18__18_ ( .D(n1744), .CK(clk), .Q(mem_18__18_) );
  DFF_X2 mem_reg_18__17_ ( .D(n1743), .CK(clk), .Q(mem_18__17_) );
  DFF_X2 mem_reg_18__16_ ( .D(n1742), .CK(clk), .Q(mem_18__16_) );
  DFF_X2 mem_reg_18__15_ ( .D(n1741), .CK(clk), .Q(mem_18__15_) );
  DFF_X2 mem_reg_18__14_ ( .D(n1740), .CK(clk), .Q(mem_18__14_) );
  DFF_X2 mem_reg_18__13_ ( .D(n1739), .CK(clk), .Q(mem_18__13_) );
  DFF_X2 mem_reg_18__12_ ( .D(n1738), .CK(clk), .Q(mem_18__12_) );
  DFF_X2 mem_reg_18__11_ ( .D(n1737), .CK(clk), .Q(mem_18__11_) );
  DFF_X2 mem_reg_18__10_ ( .D(n1736), .CK(clk), .Q(mem_18__10_) );
  DFF_X2 mem_reg_18__9_ ( .D(n1735), .CK(clk), .Q(mem_18__9_) );
  DFF_X2 mem_reg_18__8_ ( .D(n1734), .CK(clk), .Q(mem_18__8_) );
  DFF_X2 mem_reg_18__7_ ( .D(n1733), .CK(clk), .Q(mem_18__7_) );
  DFF_X2 mem_reg_18__6_ ( .D(n1732), .CK(clk), .Q(mem_18__6_) );
  DFF_X2 mem_reg_18__5_ ( .D(n1731), .CK(clk), .Q(mem_18__5_) );
  DFF_X2 mem_reg_18__4_ ( .D(n1730), .CK(clk), .Q(mem_18__4_) );
  DFF_X2 mem_reg_18__3_ ( .D(n1729), .CK(clk), .Q(mem_18__3_) );
  DFF_X2 mem_reg_18__2_ ( .D(n1728), .CK(clk), .Q(mem_18__2_) );
  DFF_X2 mem_reg_18__1_ ( .D(n1727), .CK(clk), .Q(mem_18__1_) );
  DFF_X2 mem_reg_18__0_ ( .D(n1726), .CK(clk), .Q(mem_18__0_) );
  DFF_X2 mem_reg_17__31_ ( .D(n1725), .CK(clk), .Q(mem_17__31_) );
  DFF_X2 mem_reg_17__30_ ( .D(n1724), .CK(clk), .Q(mem_17__30_) );
  DFF_X2 mem_reg_17__29_ ( .D(n1723), .CK(clk), .Q(mem_17__29_) );
  DFF_X2 mem_reg_17__28_ ( .D(n1722), .CK(clk), .Q(mem_17__28_) );
  DFF_X2 mem_reg_17__27_ ( .D(n1721), .CK(clk), .Q(mem_17__27_) );
  DFF_X2 mem_reg_17__26_ ( .D(n1720), .CK(clk), .Q(mem_17__26_) );
  DFF_X2 mem_reg_17__25_ ( .D(n1719), .CK(clk), .Q(mem_17__25_) );
  DFF_X2 mem_reg_17__24_ ( .D(n1718), .CK(clk), .Q(mem_17__24_) );
  DFF_X2 mem_reg_17__23_ ( .D(n1717), .CK(clk), .Q(mem_17__23_) );
  DFF_X2 mem_reg_17__22_ ( .D(n1716), .CK(clk), .Q(mem_17__22_) );
  DFF_X2 mem_reg_17__21_ ( .D(n1715), .CK(clk), .Q(mem_17__21_) );
  DFF_X2 mem_reg_17__20_ ( .D(n1714), .CK(clk), .Q(mem_17__20_) );
  DFF_X2 mem_reg_17__19_ ( .D(n1713), .CK(clk), .Q(mem_17__19_) );
  DFF_X2 mem_reg_17__18_ ( .D(n1712), .CK(clk), .Q(mem_17__18_) );
  DFF_X2 mem_reg_17__17_ ( .D(n1711), .CK(clk), .Q(mem_17__17_) );
  DFF_X2 mem_reg_17__16_ ( .D(n1710), .CK(clk), .Q(mem_17__16_) );
  DFF_X2 mem_reg_17__15_ ( .D(n1709), .CK(clk), .Q(mem_17__15_) );
  DFF_X2 mem_reg_17__14_ ( .D(n1708), .CK(clk), .Q(mem_17__14_) );
  DFF_X2 mem_reg_17__13_ ( .D(n1707), .CK(clk), .Q(mem_17__13_) );
  DFF_X2 mem_reg_17__12_ ( .D(n1706), .CK(clk), .Q(mem_17__12_) );
  DFF_X2 mem_reg_17__11_ ( .D(n1705), .CK(clk), .Q(mem_17__11_) );
  DFF_X2 mem_reg_17__10_ ( .D(n1704), .CK(clk), .Q(mem_17__10_) );
  DFF_X2 mem_reg_17__9_ ( .D(n1703), .CK(clk), .Q(mem_17__9_) );
  DFF_X2 mem_reg_17__8_ ( .D(n1702), .CK(clk), .Q(mem_17__8_) );
  DFF_X2 mem_reg_17__7_ ( .D(n1701), .CK(clk), .Q(mem_17__7_) );
  DFF_X2 mem_reg_17__6_ ( .D(n1700), .CK(clk), .Q(mem_17__6_) );
  DFF_X2 mem_reg_17__5_ ( .D(n1699), .CK(clk), .Q(mem_17__5_) );
  DFF_X2 mem_reg_17__4_ ( .D(n1698), .CK(clk), .Q(mem_17__4_) );
  DFF_X2 mem_reg_17__3_ ( .D(n1697), .CK(clk), .Q(mem_17__3_) );
  DFF_X2 mem_reg_17__2_ ( .D(n1696), .CK(clk), .Q(mem_17__2_) );
  DFF_X2 mem_reg_17__1_ ( .D(n1695), .CK(clk), .Q(mem_17__1_) );
  DFF_X2 mem_reg_17__0_ ( .D(n1694), .CK(clk), .Q(mem_17__0_) );
  DFF_X2 mem_reg_16__31_ ( .D(n1693), .CK(clk), .Q(mem_16__31_) );
  DFF_X2 mem_reg_16__30_ ( .D(n1692), .CK(clk), .Q(mem_16__30_) );
  DFF_X2 mem_reg_16__29_ ( .D(n1691), .CK(clk), .Q(mem_16__29_) );
  DFF_X2 mem_reg_16__28_ ( .D(n1690), .CK(clk), .Q(mem_16__28_) );
  DFF_X2 mem_reg_16__27_ ( .D(n1689), .CK(clk), .Q(mem_16__27_) );
  DFF_X2 mem_reg_16__26_ ( .D(n1688), .CK(clk), .Q(mem_16__26_) );
  DFF_X2 mem_reg_16__25_ ( .D(n1687), .CK(clk), .Q(mem_16__25_) );
  DFF_X2 mem_reg_16__24_ ( .D(n1686), .CK(clk), .Q(mem_16__24_) );
  DFF_X2 mem_reg_16__23_ ( .D(n1685), .CK(clk), .Q(mem_16__23_) );
  DFF_X2 mem_reg_16__22_ ( .D(n1684), .CK(clk), .Q(mem_16__22_) );
  DFF_X2 mem_reg_16__21_ ( .D(n1683), .CK(clk), .Q(mem_16__21_) );
  DFF_X2 mem_reg_16__20_ ( .D(n1682), .CK(clk), .Q(mem_16__20_) );
  DFF_X2 mem_reg_16__19_ ( .D(n1681), .CK(clk), .Q(mem_16__19_) );
  DFF_X2 mem_reg_16__18_ ( .D(n1680), .CK(clk), .Q(mem_16__18_) );
  DFF_X2 mem_reg_16__17_ ( .D(n1679), .CK(clk), .Q(mem_16__17_) );
  DFF_X2 mem_reg_16__16_ ( .D(n1678), .CK(clk), .Q(mem_16__16_) );
  DFF_X2 mem_reg_16__15_ ( .D(n1677), .CK(clk), .Q(mem_16__15_) );
  DFF_X2 mem_reg_16__14_ ( .D(n1676), .CK(clk), .Q(mem_16__14_) );
  DFF_X2 mem_reg_16__13_ ( .D(n1675), .CK(clk), .Q(mem_16__13_) );
  DFF_X2 mem_reg_16__12_ ( .D(n1674), .CK(clk), .Q(mem_16__12_) );
  DFF_X2 mem_reg_16__11_ ( .D(n1673), .CK(clk), .Q(mem_16__11_) );
  DFF_X2 mem_reg_16__10_ ( .D(n1672), .CK(clk), .Q(mem_16__10_) );
  DFF_X2 mem_reg_16__9_ ( .D(n1671), .CK(clk), .Q(mem_16__9_) );
  DFF_X2 mem_reg_16__8_ ( .D(n1670), .CK(clk), .Q(mem_16__8_) );
  DFF_X2 mem_reg_16__7_ ( .D(n1669), .CK(clk), .Q(mem_16__7_) );
  DFF_X2 mem_reg_16__6_ ( .D(n1668), .CK(clk), .Q(mem_16__6_) );
  DFF_X2 mem_reg_16__5_ ( .D(n1667), .CK(clk), .Q(mem_16__5_) );
  DFF_X2 mem_reg_16__4_ ( .D(n1666), .CK(clk), .Q(mem_16__4_) );
  DFF_X2 mem_reg_16__3_ ( .D(n1665), .CK(clk), .Q(mem_16__3_) );
  DFF_X2 mem_reg_16__2_ ( .D(n1664), .CK(clk), .Q(mem_16__2_) );
  DFF_X2 mem_reg_16__1_ ( .D(n1663), .CK(clk), .Q(mem_16__1_) );
  DFF_X2 mem_reg_16__0_ ( .D(n1662), .CK(clk), .Q(mem_16__0_) );
  DFF_X2 mem_reg_15__31_ ( .D(n1661), .CK(clk), .Q(mem_15__31_) );
  DFF_X2 mem_reg_15__30_ ( .D(n1660), .CK(clk), .Q(mem_15__30_) );
  DFF_X2 mem_reg_15__29_ ( .D(n1659), .CK(clk), .Q(mem_15__29_) );
  DFF_X2 mem_reg_15__28_ ( .D(n1658), .CK(clk), .Q(mem_15__28_), .QN(n2324) );
  DFF_X2 mem_reg_15__27_ ( .D(n1657), .CK(clk), .Q(mem_15__27_) );
  DFF_X2 mem_reg_15__26_ ( .D(n1656), .CK(clk), .Q(mem_15__26_) );
  DFF_X2 mem_reg_15__25_ ( .D(n1655), .CK(clk), .Q(mem_15__25_) );
  DFF_X2 mem_reg_15__24_ ( .D(n1654), .CK(clk), .Q(mem_15__24_) );
  DFF_X2 mem_reg_15__23_ ( .D(n1653), .CK(clk), .Q(mem_15__23_) );
  DFF_X2 mem_reg_15__22_ ( .D(n1652), .CK(clk), .Q(mem_15__22_) );
  DFF_X2 mem_reg_15__21_ ( .D(n1651), .CK(clk), .Q(mem_15__21_) );
  DFF_X2 mem_reg_15__20_ ( .D(n1650), .CK(clk), .Q(mem_15__20_) );
  DFF_X2 mem_reg_15__19_ ( .D(n1649), .CK(clk), .Q(mem_15__19_) );
  DFF_X2 mem_reg_15__18_ ( .D(n1648), .CK(clk), .Q(mem_15__18_) );
  DFF_X2 mem_reg_15__17_ ( .D(n1647), .CK(clk), .Q(mem_15__17_) );
  DFF_X2 mem_reg_15__16_ ( .D(n1646), .CK(clk), .Q(mem_15__16_) );
  DFF_X2 mem_reg_15__15_ ( .D(n1645), .CK(clk), .Q(mem_15__15_) );
  DFF_X2 mem_reg_15__14_ ( .D(n1644), .CK(clk), .Q(mem_15__14_) );
  DFF_X2 mem_reg_15__13_ ( .D(n1643), .CK(clk), .Q(mem_15__13_) );
  DFF_X2 mem_reg_15__12_ ( .D(n1642), .CK(clk), .Q(mem_15__12_) );
  DFF_X2 mem_reg_15__11_ ( .D(n1641), .CK(clk), .Q(mem_15__11_) );
  DFF_X2 mem_reg_15__10_ ( .D(n1640), .CK(clk), .Q(mem_15__10_) );
  DFF_X2 mem_reg_15__9_ ( .D(n1639), .CK(clk), .Q(mem_15__9_) );
  DFF_X2 mem_reg_15__8_ ( .D(n1638), .CK(clk), .Q(mem_15__8_) );
  DFF_X2 mem_reg_15__7_ ( .D(n1637), .CK(clk), .Q(mem_15__7_) );
  DFF_X2 mem_reg_15__6_ ( .D(n1636), .CK(clk), .Q(mem_15__6_) );
  DFF_X2 mem_reg_15__5_ ( .D(n1635), .CK(clk), .Q(mem_15__5_) );
  DFF_X2 mem_reg_15__4_ ( .D(n1634), .CK(clk), .Q(mem_15__4_) );
  DFF_X2 mem_reg_15__3_ ( .D(n1633), .CK(clk), .Q(mem_15__3_) );
  DFF_X2 mem_reg_15__2_ ( .D(n1632), .CK(clk), .Q(mem_15__2_) );
  DFF_X2 mem_reg_15__1_ ( .D(n1631), .CK(clk), .Q(mem_15__1_) );
  DFF_X2 mem_reg_15__0_ ( .D(n1630), .CK(clk), .Q(mem_15__0_) );
  DFF_X2 mem_reg_14__31_ ( .D(n1629), .CK(clk), .Q(mem_14__31_) );
  DFF_X2 mem_reg_14__30_ ( .D(n1628), .CK(clk), .Q(mem_14__30_) );
  DFF_X2 mem_reg_14__29_ ( .D(n1627), .CK(clk), .Q(mem_14__29_) );
  DFF_X2 mem_reg_14__28_ ( .D(n1626), .CK(clk), .Q(mem_14__28_) );
  DFF_X2 mem_reg_14__27_ ( .D(n1625), .CK(clk), .Q(mem_14__27_) );
  DFF_X2 mem_reg_14__26_ ( .D(n1624), .CK(clk), .Q(mem_14__26_) );
  DFF_X2 mem_reg_14__25_ ( .D(n1623), .CK(clk), .Q(mem_14__25_) );
  DFF_X2 mem_reg_14__24_ ( .D(n1622), .CK(clk), .Q(mem_14__24_) );
  DFF_X2 mem_reg_14__23_ ( .D(n1621), .CK(clk), .Q(mem_14__23_) );
  DFF_X2 mem_reg_14__22_ ( .D(n1620), .CK(clk), .Q(mem_14__22_) );
  DFF_X2 mem_reg_14__21_ ( .D(n1619), .CK(clk), .Q(mem_14__21_) );
  DFF_X2 mem_reg_14__20_ ( .D(n1618), .CK(clk), .Q(mem_14__20_) );
  DFF_X2 mem_reg_14__19_ ( .D(n1617), .CK(clk), .Q(mem_14__19_) );
  DFF_X2 mem_reg_14__18_ ( .D(n1616), .CK(clk), .Q(mem_14__18_) );
  DFF_X2 mem_reg_14__17_ ( .D(n1615), .CK(clk), .Q(mem_14__17_) );
  DFF_X2 mem_reg_14__16_ ( .D(n1614), .CK(clk), .Q(mem_14__16_) );
  DFF_X2 mem_reg_14__15_ ( .D(n1613), .CK(clk), .Q(mem_14__15_) );
  DFF_X2 mem_reg_14__14_ ( .D(n1612), .CK(clk), .Q(mem_14__14_) );
  DFF_X2 mem_reg_14__13_ ( .D(n1611), .CK(clk), .Q(mem_14__13_) );
  DFF_X2 mem_reg_14__12_ ( .D(n1610), .CK(clk), .Q(mem_14__12_) );
  DFF_X2 mem_reg_14__11_ ( .D(n1609), .CK(clk), .Q(mem_14__11_) );
  DFF_X2 mem_reg_14__10_ ( .D(n1608), .CK(clk), .Q(mem_14__10_) );
  DFF_X2 mem_reg_14__9_ ( .D(n1607), .CK(clk), .Q(mem_14__9_) );
  DFF_X2 mem_reg_14__8_ ( .D(n1606), .CK(clk), .Q(mem_14__8_) );
  DFF_X2 mem_reg_14__7_ ( .D(n1605), .CK(clk), .Q(mem_14__7_) );
  DFF_X2 mem_reg_14__6_ ( .D(n1604), .CK(clk), .Q(mem_14__6_) );
  DFF_X2 mem_reg_14__5_ ( .D(n1603), .CK(clk), .Q(mem_14__5_) );
  DFF_X2 mem_reg_14__4_ ( .D(n1602), .CK(clk), .Q(mem_14__4_) );
  DFF_X2 mem_reg_14__3_ ( .D(n1601), .CK(clk), .Q(mem_14__3_) );
  DFF_X2 mem_reg_14__2_ ( .D(n1600), .CK(clk), .Q(mem_14__2_) );
  DFF_X2 mem_reg_14__1_ ( .D(n1599), .CK(clk), .Q(mem_14__1_) );
  DFF_X2 mem_reg_14__0_ ( .D(n1598), .CK(clk), .Q(mem_14__0_) );
  DFF_X2 mem_reg_13__31_ ( .D(n1597), .CK(clk), .Q(mem_13__31_) );
  DFF_X2 mem_reg_13__30_ ( .D(n1596), .CK(clk), .Q(mem_13__30_) );
  DFF_X2 mem_reg_13__29_ ( .D(n1595), .CK(clk), .Q(mem_13__29_) );
  DFF_X2 mem_reg_13__28_ ( .D(n1594), .CK(clk), .Q(mem_13__28_) );
  DFF_X2 mem_reg_13__27_ ( .D(n1593), .CK(clk), .Q(mem_13__27_) );
  DFF_X2 mem_reg_13__26_ ( .D(n1592), .CK(clk), .Q(mem_13__26_) );
  DFF_X2 mem_reg_13__25_ ( .D(n1591), .CK(clk), .Q(mem_13__25_) );
  DFF_X2 mem_reg_13__24_ ( .D(n1590), .CK(clk), .Q(mem_13__24_) );
  DFF_X2 mem_reg_13__23_ ( .D(n1589), .CK(clk), .Q(mem_13__23_) );
  DFF_X2 mem_reg_13__22_ ( .D(n1588), .CK(clk), .Q(mem_13__22_) );
  DFF_X2 mem_reg_13__21_ ( .D(n1587), .CK(clk), .Q(mem_13__21_) );
  DFF_X2 mem_reg_13__20_ ( .D(n1586), .CK(clk), .Q(mem_13__20_) );
  DFF_X2 mem_reg_13__19_ ( .D(n1585), .CK(clk), .Q(mem_13__19_) );
  DFF_X2 mem_reg_13__18_ ( .D(n1584), .CK(clk), .Q(mem_13__18_) );
  DFF_X2 mem_reg_13__17_ ( .D(n1583), .CK(clk), .Q(mem_13__17_) );
  DFF_X2 mem_reg_13__16_ ( .D(n1582), .CK(clk), .Q(mem_13__16_) );
  DFF_X2 mem_reg_13__15_ ( .D(n1581), .CK(clk), .Q(mem_13__15_) );
  DFF_X2 mem_reg_13__14_ ( .D(n1580), .CK(clk), .Q(mem_13__14_) );
  DFF_X2 mem_reg_13__13_ ( .D(n1579), .CK(clk), .Q(mem_13__13_) );
  DFF_X2 mem_reg_13__12_ ( .D(n1578), .CK(clk), .Q(mem_13__12_) );
  DFF_X2 mem_reg_13__11_ ( .D(n1577), .CK(clk), .Q(mem_13__11_) );
  DFF_X2 mem_reg_13__10_ ( .D(n1576), .CK(clk), .Q(mem_13__10_) );
  DFF_X2 mem_reg_13__9_ ( .D(n1575), .CK(clk), .Q(mem_13__9_) );
  DFF_X2 mem_reg_13__8_ ( .D(n1574), .CK(clk), .Q(mem_13__8_) );
  DFF_X2 mem_reg_13__7_ ( .D(n1573), .CK(clk), .Q(mem_13__7_) );
  DFF_X2 mem_reg_13__6_ ( .D(n1572), .CK(clk), .Q(mem_13__6_) );
  DFF_X2 mem_reg_13__5_ ( .D(n1571), .CK(clk), .Q(mem_13__5_) );
  DFF_X2 mem_reg_13__4_ ( .D(n1570), .CK(clk), .Q(mem_13__4_) );
  DFF_X2 mem_reg_13__3_ ( .D(n1569), .CK(clk), .Q(mem_13__3_) );
  DFF_X2 mem_reg_13__2_ ( .D(n1568), .CK(clk), .Q(mem_13__2_) );
  DFF_X2 mem_reg_13__1_ ( .D(n1567), .CK(clk), .Q(mem_13__1_) );
  DFF_X2 mem_reg_13__0_ ( .D(n1566), .CK(clk), .Q(mem_13__0_) );
  DFF_X2 mem_reg_12__31_ ( .D(n1565), .CK(clk), .Q(mem_12__31_) );
  DFF_X2 mem_reg_12__30_ ( .D(n1564), .CK(clk), .Q(mem_12__30_) );
  DFF_X2 mem_reg_12__29_ ( .D(n1563), .CK(clk), .Q(mem_12__29_) );
  DFF_X2 mem_reg_12__28_ ( .D(n1562), .CK(clk), .Q(mem_12__28_) );
  DFF_X2 mem_reg_12__27_ ( .D(n1561), .CK(clk), .Q(mem_12__27_) );
  DFF_X2 mem_reg_12__26_ ( .D(n1560), .CK(clk), .Q(mem_12__26_) );
  DFF_X2 mem_reg_12__25_ ( .D(n1559), .CK(clk), .Q(mem_12__25_) );
  DFF_X2 mem_reg_12__24_ ( .D(n1558), .CK(clk), .Q(mem_12__24_) );
  DFF_X2 mem_reg_12__23_ ( .D(n1557), .CK(clk), .Q(mem_12__23_) );
  DFF_X2 mem_reg_12__22_ ( .D(n1556), .CK(clk), .Q(mem_12__22_) );
  DFF_X2 mem_reg_12__21_ ( .D(n1555), .CK(clk), .Q(mem_12__21_) );
  DFF_X2 mem_reg_12__20_ ( .D(n1554), .CK(clk), .Q(mem_12__20_) );
  DFF_X2 mem_reg_12__19_ ( .D(n1553), .CK(clk), .Q(mem_12__19_) );
  DFF_X2 mem_reg_12__18_ ( .D(n1552), .CK(clk), .Q(mem_12__18_) );
  DFF_X2 mem_reg_12__17_ ( .D(n1551), .CK(clk), .Q(mem_12__17_) );
  DFF_X2 mem_reg_12__16_ ( .D(n1550), .CK(clk), .Q(mem_12__16_) );
  DFF_X2 mem_reg_12__15_ ( .D(n1549), .CK(clk), .Q(mem_12__15_) );
  DFF_X2 mem_reg_12__14_ ( .D(n1548), .CK(clk), .Q(mem_12__14_) );
  DFF_X2 mem_reg_12__13_ ( .D(n1547), .CK(clk), .Q(mem_12__13_) );
  DFF_X2 mem_reg_12__12_ ( .D(n1546), .CK(clk), .Q(mem_12__12_) );
  DFF_X2 mem_reg_12__11_ ( .D(n1545), .CK(clk), .Q(mem_12__11_) );
  DFF_X2 mem_reg_12__10_ ( .D(n1544), .CK(clk), .Q(mem_12__10_) );
  DFF_X2 mem_reg_12__9_ ( .D(n1543), .CK(clk), .Q(mem_12__9_) );
  DFF_X2 mem_reg_12__8_ ( .D(n1542), .CK(clk), .Q(mem_12__8_) );
  DFF_X2 mem_reg_12__7_ ( .D(n1541), .CK(clk), .Q(mem_12__7_) );
  DFF_X2 mem_reg_12__6_ ( .D(n1540), .CK(clk), .Q(mem_12__6_) );
  DFF_X2 mem_reg_12__5_ ( .D(n1539), .CK(clk), .Q(mem_12__5_) );
  DFF_X2 mem_reg_12__4_ ( .D(n1538), .CK(clk), .Q(mem_12__4_) );
  DFF_X2 mem_reg_12__3_ ( .D(n1537), .CK(clk), .Q(mem_12__3_) );
  DFF_X2 mem_reg_12__2_ ( .D(n1536), .CK(clk), .Q(mem_12__2_) );
  DFF_X2 mem_reg_12__1_ ( .D(n1535), .CK(clk), .Q(mem_12__1_) );
  DFF_X2 mem_reg_12__0_ ( .D(n1534), .CK(clk), .Q(mem_12__0_) );
  DFF_X2 mem_reg_11__31_ ( .D(n1533), .CK(clk), .Q(mem_11__31_) );
  DFF_X2 mem_reg_11__30_ ( .D(n1532), .CK(clk), .Q(mem_11__30_) );
  DFF_X2 mem_reg_11__29_ ( .D(n1531), .CK(clk), .Q(mem_11__29_) );
  DFF_X2 mem_reg_11__28_ ( .D(n1530), .CK(clk), .Q(mem_11__28_) );
  DFF_X2 mem_reg_11__27_ ( .D(n1529), .CK(clk), .Q(mem_11__27_) );
  DFF_X2 mem_reg_11__26_ ( .D(n1528), .CK(clk), .Q(mem_11__26_) );
  DFF_X2 mem_reg_11__25_ ( .D(n1527), .CK(clk), .Q(mem_11__25_) );
  DFF_X2 mem_reg_11__24_ ( .D(n1526), .CK(clk), .Q(mem_11__24_) );
  DFF_X2 mem_reg_11__23_ ( .D(n1525), .CK(clk), .Q(mem_11__23_) );
  DFF_X2 mem_reg_11__22_ ( .D(n1524), .CK(clk), .Q(mem_11__22_) );
  DFF_X2 mem_reg_11__21_ ( .D(n1523), .CK(clk), .Q(mem_11__21_) );
  DFF_X2 mem_reg_11__20_ ( .D(n1522), .CK(clk), .Q(mem_11__20_) );
  DFF_X2 mem_reg_11__19_ ( .D(n1521), .CK(clk), .Q(mem_11__19_) );
  DFF_X2 mem_reg_11__18_ ( .D(n1520), .CK(clk), .Q(mem_11__18_) );
  DFF_X2 mem_reg_11__17_ ( .D(n1519), .CK(clk), .Q(mem_11__17_) );
  DFF_X2 mem_reg_11__16_ ( .D(n1518), .CK(clk), .Q(mem_11__16_) );
  DFF_X2 mem_reg_11__15_ ( .D(n1517), .CK(clk), .Q(mem_11__15_) );
  DFF_X2 mem_reg_11__14_ ( .D(n1516), .CK(clk), .Q(mem_11__14_) );
  DFF_X2 mem_reg_11__13_ ( .D(n1515), .CK(clk), .Q(mem_11__13_) );
  DFF_X2 mem_reg_11__12_ ( .D(n1514), .CK(clk), .Q(mem_11__12_) );
  DFF_X2 mem_reg_11__11_ ( .D(n1513), .CK(clk), .Q(mem_11__11_) );
  DFF_X2 mem_reg_11__10_ ( .D(n1512), .CK(clk), .Q(mem_11__10_) );
  DFF_X2 mem_reg_11__9_ ( .D(n1511), .CK(clk), .Q(mem_11__9_) );
  DFF_X2 mem_reg_11__8_ ( .D(n1510), .CK(clk), .Q(mem_11__8_) );
  DFF_X2 mem_reg_11__7_ ( .D(n1509), .CK(clk), .Q(mem_11__7_) );
  DFF_X2 mem_reg_11__6_ ( .D(n1508), .CK(clk), .Q(mem_11__6_) );
  DFF_X2 mem_reg_11__5_ ( .D(n1507), .CK(clk), .Q(mem_11__5_) );
  DFF_X2 mem_reg_11__4_ ( .D(n1506), .CK(clk), .Q(mem_11__4_) );
  DFF_X2 mem_reg_11__3_ ( .D(n1505), .CK(clk), .Q(mem_11__3_) );
  DFF_X2 mem_reg_11__2_ ( .D(n1504), .CK(clk), .Q(mem_11__2_) );
  DFF_X2 mem_reg_11__1_ ( .D(n1503), .CK(clk), .Q(mem_11__1_) );
  DFF_X2 mem_reg_11__0_ ( .D(n1502), .CK(clk), .Q(mem_11__0_) );
  DFF_X2 mem_reg_10__31_ ( .D(n1501), .CK(clk), .Q(mem_10__31_) );
  DFF_X2 mem_reg_10__30_ ( .D(n1500), .CK(clk), .Q(mem_10__30_) );
  DFF_X2 mem_reg_10__29_ ( .D(n1499), .CK(clk), .Q(mem_10__29_) );
  DFF_X2 mem_reg_10__28_ ( .D(n1498), .CK(clk), .Q(mem_10__28_) );
  DFF_X2 mem_reg_10__27_ ( .D(n1497), .CK(clk), .Q(mem_10__27_) );
  DFF_X2 mem_reg_10__26_ ( .D(n1496), .CK(clk), .Q(mem_10__26_) );
  DFF_X2 mem_reg_10__25_ ( .D(n1495), .CK(clk), .Q(mem_10__25_) );
  DFF_X2 mem_reg_10__24_ ( .D(n1494), .CK(clk), .Q(mem_10__24_) );
  DFF_X2 mem_reg_10__23_ ( .D(n1493), .CK(clk), .Q(mem_10__23_) );
  DFF_X2 mem_reg_10__22_ ( .D(n1492), .CK(clk), .Q(mem_10__22_) );
  DFF_X2 mem_reg_10__21_ ( .D(n1491), .CK(clk), .Q(mem_10__21_) );
  DFF_X2 mem_reg_10__20_ ( .D(n1490), .CK(clk), .Q(mem_10__20_) );
  DFF_X2 mem_reg_10__19_ ( .D(n1489), .CK(clk), .Q(mem_10__19_) );
  DFF_X2 mem_reg_10__18_ ( .D(n1488), .CK(clk), .Q(mem_10__18_) );
  DFF_X2 mem_reg_10__17_ ( .D(n1487), .CK(clk), .Q(mem_10__17_) );
  DFF_X2 mem_reg_10__16_ ( .D(n1486), .CK(clk), .Q(mem_10__16_) );
  DFF_X2 mem_reg_10__15_ ( .D(n1485), .CK(clk), .Q(mem_10__15_) );
  DFF_X2 mem_reg_10__14_ ( .D(n1484), .CK(clk), .Q(mem_10__14_) );
  DFF_X2 mem_reg_10__13_ ( .D(n1483), .CK(clk), .Q(mem_10__13_) );
  DFF_X2 mem_reg_10__12_ ( .D(n1482), .CK(clk), .Q(mem_10__12_) );
  DFF_X2 mem_reg_10__11_ ( .D(n1481), .CK(clk), .Q(mem_10__11_) );
  DFF_X2 mem_reg_10__10_ ( .D(n1480), .CK(clk), .Q(mem_10__10_) );
  DFF_X2 mem_reg_10__9_ ( .D(n1479), .CK(clk), .Q(mem_10__9_) );
  DFF_X2 mem_reg_10__8_ ( .D(n1478), .CK(clk), .Q(mem_10__8_) );
  DFF_X2 mem_reg_10__7_ ( .D(n1477), .CK(clk), .Q(mem_10__7_) );
  DFF_X2 mem_reg_10__6_ ( .D(n1476), .CK(clk), .Q(mem_10__6_) );
  DFF_X2 mem_reg_10__5_ ( .D(n1475), .CK(clk), .Q(mem_10__5_) );
  DFF_X2 mem_reg_10__4_ ( .D(n1474), .CK(clk), .Q(mem_10__4_) );
  DFF_X2 mem_reg_10__3_ ( .D(n1473), .CK(clk), .Q(mem_10__3_) );
  DFF_X2 mem_reg_10__2_ ( .D(n1472), .CK(clk), .Q(mem_10__2_) );
  DFF_X2 mem_reg_10__1_ ( .D(n1471), .CK(clk), .Q(mem_10__1_) );
  DFF_X2 mem_reg_10__0_ ( .D(n1470), .CK(clk), .Q(mem_10__0_) );
  DFF_X2 mem_reg_9__31_ ( .D(n1469), .CK(clk), .Q(mem_9__31_) );
  DFF_X2 mem_reg_9__30_ ( .D(n1468), .CK(clk), .Q(mem_9__30_) );
  DFF_X2 mem_reg_9__29_ ( .D(n1467), .CK(clk), .Q(mem_9__29_) );
  DFF_X2 mem_reg_9__28_ ( .D(n1466), .CK(clk), .Q(mem_9__28_) );
  DFF_X2 mem_reg_9__27_ ( .D(n1465), .CK(clk), .Q(mem_9__27_) );
  DFF_X2 mem_reg_9__26_ ( .D(n1464), .CK(clk), .Q(mem_9__26_) );
  DFF_X2 mem_reg_9__25_ ( .D(n1463), .CK(clk), .Q(mem_9__25_) );
  DFF_X2 mem_reg_9__24_ ( .D(n1462), .CK(clk), .Q(mem_9__24_) );
  DFF_X2 mem_reg_9__23_ ( .D(n1461), .CK(clk), .Q(mem_9__23_) );
  DFF_X2 mem_reg_9__22_ ( .D(n1460), .CK(clk), .Q(mem_9__22_) );
  DFF_X2 mem_reg_9__21_ ( .D(n1459), .CK(clk), .Q(mem_9__21_) );
  DFF_X2 mem_reg_9__20_ ( .D(n1458), .CK(clk), .Q(mem_9__20_) );
  DFF_X2 mem_reg_9__19_ ( .D(n1457), .CK(clk), .Q(mem_9__19_) );
  DFF_X2 mem_reg_9__18_ ( .D(n1456), .CK(clk), .Q(mem_9__18_) );
  DFF_X2 mem_reg_9__17_ ( .D(n1455), .CK(clk), .Q(mem_9__17_) );
  DFF_X2 mem_reg_9__16_ ( .D(n1454), .CK(clk), .Q(mem_9__16_) );
  DFF_X2 mem_reg_9__15_ ( .D(n1453), .CK(clk), .Q(mem_9__15_) );
  DFF_X2 mem_reg_9__14_ ( .D(n1452), .CK(clk), .Q(mem_9__14_) );
  DFF_X2 mem_reg_9__13_ ( .D(n1451), .CK(clk), .Q(mem_9__13_) );
  DFF_X2 mem_reg_9__12_ ( .D(n1450), .CK(clk), .Q(mem_9__12_) );
  DFF_X2 mem_reg_9__11_ ( .D(n1449), .CK(clk), .Q(mem_9__11_) );
  DFF_X2 mem_reg_9__10_ ( .D(n1448), .CK(clk), .Q(mem_9__10_) );
  DFF_X2 mem_reg_9__9_ ( .D(n1447), .CK(clk), .Q(mem_9__9_) );
  DFF_X2 mem_reg_9__8_ ( .D(n1446), .CK(clk), .Q(mem_9__8_) );
  DFF_X2 mem_reg_9__7_ ( .D(n1445), .CK(clk), .Q(mem_9__7_) );
  DFF_X2 mem_reg_9__6_ ( .D(n1444), .CK(clk), .Q(mem_9__6_) );
  DFF_X2 mem_reg_9__5_ ( .D(n1443), .CK(clk), .Q(mem_9__5_) );
  DFF_X2 mem_reg_9__4_ ( .D(n1442), .CK(clk), .Q(mem_9__4_) );
  DFF_X2 mem_reg_9__3_ ( .D(n1441), .CK(clk), .Q(mem_9__3_) );
  DFF_X2 mem_reg_9__2_ ( .D(n1440), .CK(clk), .Q(mem_9__2_) );
  DFF_X2 mem_reg_9__1_ ( .D(n1439), .CK(clk), .Q(mem_9__1_) );
  DFF_X2 mem_reg_9__0_ ( .D(n1438), .CK(clk), .Q(mem_9__0_) );
  DFF_X2 mem_reg_8__31_ ( .D(n1437), .CK(clk), .Q(mem_8__31_) );
  DFF_X2 mem_reg_8__30_ ( .D(n1436), .CK(clk), .Q(mem_8__30_) );
  DFF_X2 mem_reg_8__29_ ( .D(n1435), .CK(clk), .Q(mem_8__29_) );
  DFF_X2 mem_reg_8__28_ ( .D(n1434), .CK(clk), .Q(mem_8__28_) );
  DFF_X2 mem_reg_8__27_ ( .D(n1433), .CK(clk), .Q(mem_8__27_) );
  DFF_X2 mem_reg_8__26_ ( .D(n1432), .CK(clk), .Q(mem_8__26_) );
  DFF_X2 mem_reg_8__25_ ( .D(n1431), .CK(clk), .Q(mem_8__25_) );
  DFF_X2 mem_reg_8__24_ ( .D(n1430), .CK(clk), .Q(mem_8__24_) );
  DFF_X2 mem_reg_8__23_ ( .D(n1429), .CK(clk), .Q(mem_8__23_) );
  DFF_X2 mem_reg_8__22_ ( .D(n1428), .CK(clk), .Q(mem_8__22_) );
  DFF_X2 mem_reg_8__21_ ( .D(n1427), .CK(clk), .Q(mem_8__21_) );
  DFF_X2 mem_reg_8__20_ ( .D(n1426), .CK(clk), .Q(mem_8__20_) );
  DFF_X2 mem_reg_8__19_ ( .D(n1425), .CK(clk), .Q(mem_8__19_) );
  DFF_X2 mem_reg_8__18_ ( .D(n1424), .CK(clk), .Q(mem_8__18_) );
  DFF_X2 mem_reg_8__17_ ( .D(n1423), .CK(clk), .Q(mem_8__17_) );
  DFF_X2 mem_reg_8__16_ ( .D(n1422), .CK(clk), .Q(mem_8__16_) );
  DFF_X2 mem_reg_8__15_ ( .D(n1421), .CK(clk), .Q(mem_8__15_) );
  DFF_X2 mem_reg_8__14_ ( .D(n1420), .CK(clk), .Q(mem_8__14_) );
  DFF_X2 mem_reg_8__13_ ( .D(n1419), .CK(clk), .Q(mem_8__13_) );
  DFF_X2 mem_reg_8__12_ ( .D(n1418), .CK(clk), .Q(mem_8__12_) );
  DFF_X2 mem_reg_8__11_ ( .D(n1417), .CK(clk), .Q(mem_8__11_) );
  DFF_X2 mem_reg_8__10_ ( .D(n1416), .CK(clk), .Q(mem_8__10_) );
  DFF_X2 mem_reg_8__9_ ( .D(n1415), .CK(clk), .Q(mem_8__9_) );
  DFF_X2 mem_reg_8__8_ ( .D(n1414), .CK(clk), .Q(mem_8__8_) );
  DFF_X2 mem_reg_8__7_ ( .D(n1413), .CK(clk), .Q(mem_8__7_) );
  DFF_X2 mem_reg_8__6_ ( .D(n1412), .CK(clk), .Q(mem_8__6_) );
  DFF_X2 mem_reg_8__5_ ( .D(n1411), .CK(clk), .Q(mem_8__5_) );
  DFF_X2 mem_reg_8__4_ ( .D(n1410), .CK(clk), .Q(mem_8__4_) );
  DFF_X2 mem_reg_8__3_ ( .D(n1409), .CK(clk), .Q(mem_8__3_) );
  DFF_X2 mem_reg_8__2_ ( .D(n1408), .CK(clk), .Q(mem_8__2_) );
  DFF_X2 mem_reg_8__1_ ( .D(n1407), .CK(clk), .Q(mem_8__1_) );
  DFF_X2 mem_reg_8__0_ ( .D(n1406), .CK(clk), .Q(mem_8__0_) );
  DFF_X2 mem_reg_7__31_ ( .D(n1405), .CK(clk), .Q(mem_7__31_) );
  DFF_X2 mem_reg_7__30_ ( .D(n1404), .CK(clk), .Q(mem_7__30_) );
  DFF_X2 mem_reg_7__29_ ( .D(n1403), .CK(clk), .Q(mem_7__29_) );
  DFF_X2 mem_reg_7__28_ ( .D(n1402), .CK(clk), .Q(mem_7__28_) );
  DFF_X2 mem_reg_7__27_ ( .D(n1401), .CK(clk), .Q(mem_7__27_) );
  DFF_X2 mem_reg_7__26_ ( .D(n1400), .CK(clk), .Q(mem_7__26_) );
  DFF_X2 mem_reg_7__25_ ( .D(n1399), .CK(clk), .Q(mem_7__25_) );
  DFF_X2 mem_reg_7__24_ ( .D(n1398), .CK(clk), .Q(mem_7__24_) );
  DFF_X2 mem_reg_7__23_ ( .D(n1397), .CK(clk), .Q(mem_7__23_) );
  DFF_X2 mem_reg_7__22_ ( .D(n1396), .CK(clk), .Q(mem_7__22_) );
  DFF_X2 mem_reg_7__21_ ( .D(n1395), .CK(clk), .Q(mem_7__21_) );
  DFF_X2 mem_reg_7__20_ ( .D(n1394), .CK(clk), .Q(mem_7__20_) );
  DFF_X2 mem_reg_7__19_ ( .D(n1393), .CK(clk), .Q(mem_7__19_) );
  DFF_X2 mem_reg_7__18_ ( .D(n1392), .CK(clk), .Q(mem_7__18_) );
  DFF_X2 mem_reg_7__17_ ( .D(n1391), .CK(clk), .Q(mem_7__17_) );
  DFF_X2 mem_reg_7__16_ ( .D(n1390), .CK(clk), .Q(mem_7__16_) );
  DFF_X2 mem_reg_7__15_ ( .D(n1389), .CK(clk), .Q(mem_7__15_) );
  DFF_X2 mem_reg_7__14_ ( .D(n1388), .CK(clk), .Q(mem_7__14_) );
  DFF_X2 mem_reg_7__13_ ( .D(n1387), .CK(clk), .Q(mem_7__13_) );
  DFF_X2 mem_reg_7__12_ ( .D(n1386), .CK(clk), .Q(mem_7__12_) );
  DFF_X2 mem_reg_7__11_ ( .D(n1385), .CK(clk), .Q(mem_7__11_) );
  DFF_X2 mem_reg_7__10_ ( .D(n1384), .CK(clk), .Q(mem_7__10_) );
  DFF_X2 mem_reg_7__9_ ( .D(n1383), .CK(clk), .Q(mem_7__9_) );
  DFF_X2 mem_reg_7__8_ ( .D(n1382), .CK(clk), .Q(mem_7__8_) );
  DFF_X2 mem_reg_7__7_ ( .D(n1381), .CK(clk), .Q(mem_7__7_) );
  DFF_X2 mem_reg_7__6_ ( .D(n1380), .CK(clk), .Q(mem_7__6_) );
  DFF_X2 mem_reg_7__5_ ( .D(n1379), .CK(clk), .Q(mem_7__5_) );
  DFF_X2 mem_reg_7__4_ ( .D(n1378), .CK(clk), .Q(mem_7__4_) );
  DFF_X2 mem_reg_7__3_ ( .D(n1377), .CK(clk), .Q(mem_7__3_) );
  DFF_X2 mem_reg_7__2_ ( .D(n1376), .CK(clk), .Q(mem_7__2_) );
  DFF_X2 mem_reg_7__1_ ( .D(n1375), .CK(clk), .Q(mem_7__1_) );
  DFF_X2 mem_reg_7__0_ ( .D(n1374), .CK(clk), .Q(mem_7__0_) );
  DFF_X2 mem_reg_6__31_ ( .D(n1373), .CK(clk), .Q(mem_6__31_) );
  DFF_X2 mem_reg_6__30_ ( .D(n1372), .CK(clk), .Q(mem_6__30_) );
  DFF_X2 mem_reg_6__29_ ( .D(n1371), .CK(clk), .Q(mem_6__29_) );
  DFF_X2 mem_reg_6__28_ ( .D(n1370), .CK(clk), .Q(mem_6__28_) );
  DFF_X2 mem_reg_6__27_ ( .D(n1369), .CK(clk), .Q(mem_6__27_) );
  DFF_X2 mem_reg_6__26_ ( .D(n1368), .CK(clk), .Q(mem_6__26_) );
  DFF_X2 mem_reg_6__25_ ( .D(n1367), .CK(clk), .Q(mem_6__25_) );
  DFF_X2 mem_reg_6__24_ ( .D(n1366), .CK(clk), .Q(mem_6__24_) );
  DFF_X2 mem_reg_6__23_ ( .D(n1365), .CK(clk), .Q(mem_6__23_) );
  DFF_X2 mem_reg_6__22_ ( .D(n1364), .CK(clk), .Q(mem_6__22_) );
  DFF_X2 mem_reg_6__21_ ( .D(n1363), .CK(clk), .Q(mem_6__21_) );
  DFF_X2 mem_reg_6__20_ ( .D(n1362), .CK(clk), .Q(mem_6__20_) );
  DFF_X2 mem_reg_6__19_ ( .D(n1361), .CK(clk), .Q(mem_6__19_) );
  DFF_X2 mem_reg_6__18_ ( .D(n1360), .CK(clk), .Q(mem_6__18_) );
  DFF_X2 mem_reg_6__17_ ( .D(n1359), .CK(clk), .Q(mem_6__17_) );
  DFF_X2 mem_reg_6__16_ ( .D(n1358), .CK(clk), .Q(mem_6__16_) );
  DFF_X2 mem_reg_6__15_ ( .D(n1357), .CK(clk), .Q(mem_6__15_) );
  DFF_X2 mem_reg_6__14_ ( .D(n1356), .CK(clk), .Q(mem_6__14_) );
  DFF_X2 mem_reg_6__13_ ( .D(n1355), .CK(clk), .Q(mem_6__13_) );
  DFF_X2 mem_reg_6__12_ ( .D(n1354), .CK(clk), .Q(mem_6__12_) );
  DFF_X2 mem_reg_6__11_ ( .D(n1353), .CK(clk), .Q(mem_6__11_) );
  DFF_X2 mem_reg_6__10_ ( .D(n1352), .CK(clk), .Q(mem_6__10_) );
  DFF_X2 mem_reg_6__9_ ( .D(n1351), .CK(clk), .Q(mem_6__9_) );
  DFF_X2 mem_reg_6__8_ ( .D(n1350), .CK(clk), .Q(mem_6__8_) );
  DFF_X2 mem_reg_6__7_ ( .D(n1349), .CK(clk), .Q(mem_6__7_) );
  DFF_X2 mem_reg_6__6_ ( .D(n1348), .CK(clk), .Q(mem_6__6_) );
  DFF_X2 mem_reg_6__5_ ( .D(n1347), .CK(clk), .Q(mem_6__5_) );
  DFF_X2 mem_reg_6__4_ ( .D(n1346), .CK(clk), .Q(mem_6__4_) );
  DFF_X2 mem_reg_6__3_ ( .D(n1345), .CK(clk), .Q(mem_6__3_) );
  DFF_X2 mem_reg_6__2_ ( .D(n1344), .CK(clk), .Q(mem_6__2_) );
  DFF_X2 mem_reg_6__1_ ( .D(n1343), .CK(clk), .Q(mem_6__1_) );
  DFF_X2 mem_reg_6__0_ ( .D(n1342), .CK(clk), .Q(mem_6__0_) );
  DFF_X2 mem_reg_5__31_ ( .D(n1341), .CK(clk), .Q(mem_5__31_) );
  DFF_X2 mem_reg_5__30_ ( .D(n1340), .CK(clk), .Q(mem_5__30_) );
  DFF_X2 mem_reg_5__29_ ( .D(n1339), .CK(clk), .Q(mem_5__29_) );
  DFF_X2 mem_reg_5__28_ ( .D(n1338), .CK(clk), .Q(mem_5__28_) );
  DFF_X2 mem_reg_5__27_ ( .D(n1337), .CK(clk), .Q(mem_5__27_) );
  DFF_X2 mem_reg_5__26_ ( .D(n1336), .CK(clk), .Q(mem_5__26_) );
  DFF_X2 mem_reg_5__25_ ( .D(n1335), .CK(clk), .Q(mem_5__25_) );
  DFF_X2 mem_reg_5__24_ ( .D(n1334), .CK(clk), .Q(mem_5__24_) );
  DFF_X2 mem_reg_5__23_ ( .D(n1333), .CK(clk), .Q(mem_5__23_) );
  DFF_X2 mem_reg_5__22_ ( .D(n1332), .CK(clk), .Q(mem_5__22_) );
  DFF_X2 mem_reg_5__21_ ( .D(n1331), .CK(clk), .Q(mem_5__21_) );
  DFF_X2 mem_reg_5__20_ ( .D(n1330), .CK(clk), .Q(mem_5__20_) );
  DFF_X2 mem_reg_5__19_ ( .D(n1329), .CK(clk), .Q(mem_5__19_) );
  DFF_X2 mem_reg_5__18_ ( .D(n1328), .CK(clk), .Q(mem_5__18_) );
  DFF_X2 mem_reg_5__17_ ( .D(n1327), .CK(clk), .Q(mem_5__17_) );
  DFF_X2 mem_reg_5__16_ ( .D(n1326), .CK(clk), .Q(mem_5__16_) );
  DFF_X2 mem_reg_5__15_ ( .D(n1325), .CK(clk), .Q(mem_5__15_) );
  DFF_X2 mem_reg_5__14_ ( .D(n1324), .CK(clk), .Q(mem_5__14_) );
  DFF_X2 mem_reg_5__13_ ( .D(n1323), .CK(clk), .Q(mem_5__13_) );
  DFF_X2 mem_reg_5__12_ ( .D(n1322), .CK(clk), .Q(mem_5__12_) );
  DFF_X2 mem_reg_5__11_ ( .D(n1321), .CK(clk), .Q(mem_5__11_) );
  DFF_X2 mem_reg_5__10_ ( .D(n1320), .CK(clk), .Q(mem_5__10_) );
  DFF_X2 mem_reg_5__9_ ( .D(n1319), .CK(clk), .Q(mem_5__9_) );
  DFF_X2 mem_reg_5__8_ ( .D(n1318), .CK(clk), .Q(mem_5__8_) );
  DFF_X2 mem_reg_5__7_ ( .D(n1317), .CK(clk), .Q(mem_5__7_) );
  DFF_X2 mem_reg_5__6_ ( .D(n1316), .CK(clk), .Q(mem_5__6_) );
  DFF_X2 mem_reg_5__5_ ( .D(n1315), .CK(clk), .Q(mem_5__5_) );
  DFF_X2 mem_reg_5__4_ ( .D(n1314), .CK(clk), .Q(mem_5__4_) );
  DFF_X2 mem_reg_5__3_ ( .D(n1313), .CK(clk), .Q(mem_5__3_) );
  DFF_X2 mem_reg_5__2_ ( .D(n1312), .CK(clk), .Q(mem_5__2_) );
  DFF_X2 mem_reg_5__1_ ( .D(n1311), .CK(clk), .Q(mem_5__1_) );
  DFF_X2 mem_reg_5__0_ ( .D(n1310), .CK(clk), .Q(mem_5__0_) );
  DFF_X2 mem_reg_4__31_ ( .D(n1309), .CK(clk), .Q(mem_4__31_) );
  DFF_X2 mem_reg_4__30_ ( .D(n1308), .CK(clk), .Q(mem_4__30_) );
  DFF_X2 mem_reg_4__29_ ( .D(n1307), .CK(clk), .Q(mem_4__29_) );
  DFF_X2 mem_reg_4__28_ ( .D(n1306), .CK(clk), .Q(mem_4__28_) );
  DFF_X2 mem_reg_4__27_ ( .D(n1305), .CK(clk), .Q(mem_4__27_) );
  DFF_X2 mem_reg_4__26_ ( .D(n1304), .CK(clk), .Q(mem_4__26_) );
  DFF_X2 mem_reg_4__25_ ( .D(n1303), .CK(clk), .Q(mem_4__25_) );
  DFF_X2 mem_reg_4__24_ ( .D(n1302), .CK(clk), .Q(mem_4__24_) );
  DFF_X2 mem_reg_4__23_ ( .D(n1301), .CK(clk), .Q(mem_4__23_) );
  DFF_X2 mem_reg_4__22_ ( .D(n1300), .CK(clk), .Q(mem_4__22_) );
  DFF_X2 mem_reg_4__21_ ( .D(n1299), .CK(clk), .Q(mem_4__21_) );
  DFF_X2 mem_reg_4__20_ ( .D(n1298), .CK(clk), .Q(mem_4__20_) );
  DFF_X2 mem_reg_4__19_ ( .D(n1297), .CK(clk), .Q(mem_4__19_) );
  DFF_X2 mem_reg_4__18_ ( .D(n1296), .CK(clk), .Q(mem_4__18_) );
  DFF_X2 mem_reg_4__17_ ( .D(n1295), .CK(clk), .Q(mem_4__17_) );
  DFF_X2 mem_reg_4__16_ ( .D(n1294), .CK(clk), .Q(mem_4__16_) );
  DFF_X2 mem_reg_4__15_ ( .D(n1293), .CK(clk), .Q(mem_4__15_) );
  DFF_X2 mem_reg_4__14_ ( .D(n1292), .CK(clk), .Q(mem_4__14_) );
  DFF_X2 mem_reg_4__13_ ( .D(n1291), .CK(clk), .Q(mem_4__13_) );
  DFF_X2 mem_reg_4__12_ ( .D(n1290), .CK(clk), .Q(mem_4__12_) );
  DFF_X2 mem_reg_4__11_ ( .D(n1289), .CK(clk), .Q(mem_4__11_) );
  DFF_X2 mem_reg_4__10_ ( .D(n1288), .CK(clk), .Q(mem_4__10_) );
  DFF_X2 mem_reg_4__9_ ( .D(n1287), .CK(clk), .Q(mem_4__9_) );
  DFF_X2 mem_reg_4__8_ ( .D(n1286), .CK(clk), .Q(mem_4__8_) );
  DFF_X2 mem_reg_4__7_ ( .D(n1285), .CK(clk), .Q(mem_4__7_) );
  DFF_X2 mem_reg_4__6_ ( .D(n1284), .CK(clk), .Q(mem_4__6_) );
  DFF_X2 mem_reg_4__5_ ( .D(n1283), .CK(clk), .Q(mem_4__5_) );
  DFF_X2 mem_reg_4__4_ ( .D(n1282), .CK(clk), .Q(mem_4__4_) );
  DFF_X2 mem_reg_4__3_ ( .D(n1281), .CK(clk), .Q(mem_4__3_) );
  DFF_X2 mem_reg_4__2_ ( .D(n1280), .CK(clk), .Q(mem_4__2_) );
  DFF_X2 mem_reg_4__1_ ( .D(n1279), .CK(clk), .Q(mem_4__1_) );
  DFF_X2 mem_reg_4__0_ ( .D(n1278), .CK(clk), .Q(mem_4__0_) );
  DFF_X2 mem_reg_3__31_ ( .D(n1277), .CK(clk), .Q(mem_3__31_) );
  DFF_X2 mem_reg_3__30_ ( .D(n1276), .CK(clk), .Q(mem_3__30_) );
  DFF_X2 mem_reg_3__29_ ( .D(n1275), .CK(clk), .Q(mem_3__29_) );
  DFF_X2 mem_reg_3__28_ ( .D(n1274), .CK(clk), .Q(mem_3__28_) );
  DFF_X2 mem_reg_3__27_ ( .D(n1273), .CK(clk), .Q(mem_3__27_) );
  DFF_X2 mem_reg_3__26_ ( .D(n1272), .CK(clk), .Q(mem_3__26_) );
  DFF_X2 mem_reg_3__25_ ( .D(n1271), .CK(clk), .Q(mem_3__25_) );
  DFF_X2 mem_reg_3__24_ ( .D(n1270), .CK(clk), .Q(mem_3__24_) );
  DFF_X2 mem_reg_3__23_ ( .D(n1269), .CK(clk), .Q(mem_3__23_) );
  DFF_X2 mem_reg_3__22_ ( .D(n1268), .CK(clk), .Q(mem_3__22_) );
  DFF_X2 mem_reg_3__21_ ( .D(n1267), .CK(clk), .Q(mem_3__21_) );
  DFF_X2 mem_reg_3__20_ ( .D(n1266), .CK(clk), .Q(mem_3__20_) );
  DFF_X2 mem_reg_3__19_ ( .D(n1265), .CK(clk), .Q(mem_3__19_) );
  DFF_X2 mem_reg_3__18_ ( .D(n1264), .CK(clk), .Q(mem_3__18_) );
  DFF_X2 mem_reg_3__17_ ( .D(n1263), .CK(clk), .Q(mem_3__17_) );
  DFF_X2 mem_reg_3__16_ ( .D(n1262), .CK(clk), .Q(mem_3__16_) );
  DFF_X2 mem_reg_3__15_ ( .D(n1261), .CK(clk), .Q(mem_3__15_) );
  DFF_X2 mem_reg_3__14_ ( .D(n1260), .CK(clk), .Q(mem_3__14_) );
  DFF_X2 mem_reg_3__13_ ( .D(n1259), .CK(clk), .Q(mem_3__13_) );
  DFF_X2 mem_reg_3__12_ ( .D(n1258), .CK(clk), .Q(mem_3__12_) );
  DFF_X2 mem_reg_3__11_ ( .D(n1257), .CK(clk), .Q(mem_3__11_) );
  DFF_X2 mem_reg_3__10_ ( .D(n1256), .CK(clk), .Q(mem_3__10_) );
  DFF_X2 mem_reg_3__9_ ( .D(n1255), .CK(clk), .Q(mem_3__9_) );
  DFF_X2 mem_reg_3__8_ ( .D(n1254), .CK(clk), .Q(mem_3__8_) );
  DFF_X2 mem_reg_3__7_ ( .D(n1253), .CK(clk), .Q(mem_3__7_) );
  DFF_X2 mem_reg_3__6_ ( .D(n1252), .CK(clk), .Q(mem_3__6_) );
  DFF_X2 mem_reg_3__5_ ( .D(n1251), .CK(clk), .Q(mem_3__5_) );
  DFF_X2 mem_reg_3__4_ ( .D(n1250), .CK(clk), .Q(mem_3__4_) );
  DFF_X2 mem_reg_3__3_ ( .D(n1249), .CK(clk), .Q(mem_3__3_) );
  DFF_X2 mem_reg_3__2_ ( .D(n1248), .CK(clk), .Q(mem_3__2_) );
  DFF_X2 mem_reg_3__1_ ( .D(n1247), .CK(clk), .Q(mem_3__1_) );
  DFF_X2 mem_reg_3__0_ ( .D(n1246), .CK(clk), .Q(mem_3__0_) );
  DFF_X2 mem_reg_2__31_ ( .D(n1245), .CK(clk), .Q(mem_2__31_) );
  DFF_X2 mem_reg_2__30_ ( .D(n1244), .CK(clk), .Q(mem_2__30_) );
  DFF_X2 mem_reg_2__29_ ( .D(n1243), .CK(clk), .Q(mem_2__29_) );
  DFF_X2 mem_reg_2__28_ ( .D(n1242), .CK(clk), .Q(mem_2__28_) );
  DFF_X2 mem_reg_2__27_ ( .D(n1241), .CK(clk), .Q(mem_2__27_) );
  DFF_X2 mem_reg_2__26_ ( .D(n1240), .CK(clk), .Q(mem_2__26_) );
  DFF_X2 mem_reg_2__25_ ( .D(n1239), .CK(clk), .Q(mem_2__25_) );
  DFF_X2 mem_reg_2__24_ ( .D(n1238), .CK(clk), .Q(mem_2__24_) );
  DFF_X2 mem_reg_2__23_ ( .D(n1237), .CK(clk), .Q(mem_2__23_) );
  DFF_X2 mem_reg_2__22_ ( .D(n1236), .CK(clk), .Q(mem_2__22_) );
  DFF_X2 mem_reg_2__21_ ( .D(n1235), .CK(clk), .Q(mem_2__21_) );
  DFF_X2 mem_reg_2__20_ ( .D(n1234), .CK(clk), .Q(mem_2__20_) );
  DFF_X2 mem_reg_2__19_ ( .D(n1233), .CK(clk), .Q(mem_2__19_) );
  DFF_X2 mem_reg_2__18_ ( .D(n1232), .CK(clk), .Q(mem_2__18_) );
  DFF_X2 mem_reg_2__17_ ( .D(n1231), .CK(clk), .Q(mem_2__17_) );
  DFF_X2 mem_reg_2__16_ ( .D(n1230), .CK(clk), .Q(mem_2__16_) );
  DFF_X2 mem_reg_2__15_ ( .D(n1229), .CK(clk), .Q(mem_2__15_) );
  DFF_X2 mem_reg_2__14_ ( .D(n1228), .CK(clk), .Q(mem_2__14_) );
  DFF_X2 mem_reg_2__13_ ( .D(n1227), .CK(clk), .Q(mem_2__13_) );
  DFF_X2 mem_reg_2__12_ ( .D(n1226), .CK(clk), .Q(mem_2__12_) );
  DFF_X2 mem_reg_2__11_ ( .D(n1225), .CK(clk), .Q(mem_2__11_) );
  DFF_X2 mem_reg_2__10_ ( .D(n1224), .CK(clk), .Q(mem_2__10_) );
  DFF_X2 mem_reg_2__9_ ( .D(n1223), .CK(clk), .Q(mem_2__9_) );
  DFF_X2 mem_reg_2__8_ ( .D(n1222), .CK(clk), .Q(mem_2__8_) );
  DFF_X2 mem_reg_2__7_ ( .D(n1221), .CK(clk), .Q(mem_2__7_) );
  DFF_X2 mem_reg_2__6_ ( .D(n1220), .CK(clk), .Q(mem_2__6_) );
  DFF_X2 mem_reg_2__5_ ( .D(n1219), .CK(clk), .Q(mem_2__5_) );
  DFF_X2 mem_reg_2__4_ ( .D(n1218), .CK(clk), .Q(mem_2__4_) );
  DFF_X2 mem_reg_2__3_ ( .D(n1217), .CK(clk), .Q(mem_2__3_) );
  DFF_X2 mem_reg_2__2_ ( .D(n1216), .CK(clk), .Q(mem_2__2_) );
  DFF_X2 mem_reg_2__1_ ( .D(n1215), .CK(clk), .Q(mem_2__1_) );
  DFF_X2 mem_reg_2__0_ ( .D(n1214), .CK(clk), .Q(mem_2__0_) );
  DFF_X2 mem_reg_1__31_ ( .D(n1213), .CK(clk), .Q(mem_1__31_) );
  DFF_X2 mem_reg_1__30_ ( .D(n1212), .CK(clk), .Q(mem_1__30_) );
  DFF_X2 mem_reg_1__29_ ( .D(n1211), .CK(clk), .Q(mem_1__29_) );
  DFF_X2 mem_reg_1__28_ ( .D(n1210), .CK(clk), .Q(mem_1__28_) );
  DFF_X2 mem_reg_1__27_ ( .D(n1209), .CK(clk), .Q(mem_1__27_) );
  DFF_X2 mem_reg_1__26_ ( .D(n1208), .CK(clk), .Q(mem_1__26_) );
  DFF_X2 mem_reg_1__25_ ( .D(n1207), .CK(clk), .Q(mem_1__25_) );
  DFF_X2 mem_reg_1__24_ ( .D(n1206), .CK(clk), .Q(mem_1__24_) );
  DFF_X2 mem_reg_1__23_ ( .D(n1205), .CK(clk), .Q(mem_1__23_) );
  DFF_X2 mem_reg_1__22_ ( .D(n1204), .CK(clk), .Q(mem_1__22_) );
  DFF_X2 mem_reg_1__21_ ( .D(n1203), .CK(clk), .Q(mem_1__21_) );
  DFF_X2 mem_reg_1__20_ ( .D(n1202), .CK(clk), .Q(mem_1__20_) );
  DFF_X2 mem_reg_1__19_ ( .D(n1201), .CK(clk), .Q(mem_1__19_) );
  DFF_X2 mem_reg_1__18_ ( .D(n1200), .CK(clk), .Q(mem_1__18_) );
  DFF_X2 mem_reg_1__17_ ( .D(n1199), .CK(clk), .Q(mem_1__17_) );
  DFF_X2 mem_reg_1__16_ ( .D(n1198), .CK(clk), .Q(mem_1__16_) );
  DFF_X2 mem_reg_1__15_ ( .D(n1197), .CK(clk), .Q(mem_1__15_) );
  DFF_X2 mem_reg_1__14_ ( .D(n1196), .CK(clk), .Q(mem_1__14_) );
  DFF_X2 mem_reg_1__13_ ( .D(n1195), .CK(clk), .Q(mem_1__13_) );
  DFF_X2 mem_reg_1__12_ ( .D(n1194), .CK(clk), .Q(mem_1__12_) );
  DFF_X2 mem_reg_1__11_ ( .D(n1193), .CK(clk), .Q(mem_1__11_) );
  DFF_X2 mem_reg_1__10_ ( .D(n1192), .CK(clk), .Q(mem_1__10_) );
  DFF_X2 mem_reg_1__9_ ( .D(n1191), .CK(clk), .Q(mem_1__9_) );
  DFF_X2 mem_reg_1__8_ ( .D(n1190), .CK(clk), .Q(mem_1__8_) );
  DFF_X2 mem_reg_1__7_ ( .D(n1189), .CK(clk), .Q(mem_1__7_) );
  DFF_X2 mem_reg_1__6_ ( .D(n1188), .CK(clk), .Q(mem_1__6_) );
  DFF_X2 mem_reg_1__5_ ( .D(n1187), .CK(clk), .Q(mem_1__5_) );
  DFF_X2 mem_reg_1__4_ ( .D(n1186), .CK(clk), .Q(mem_1__4_) );
  DFF_X2 mem_reg_1__3_ ( .D(n1185), .CK(clk), .Q(mem_1__3_) );
  DFF_X2 mem_reg_1__2_ ( .D(n1184), .CK(clk), .Q(mem_1__2_) );
  DFF_X2 mem_reg_1__1_ ( .D(n1183), .CK(clk), .Q(mem_1__1_) );
  DFF_X2 mem_reg_1__0_ ( .D(n1182), .CK(clk), .Q(mem_1__0_) );
  DFF_X2 mem_reg_0__31_ ( .D(n1181), .CK(clk), .Q(mem_0__31_) );
  DFF_X2 mem_reg_0__30_ ( .D(n1180), .CK(clk), .Q(mem_0__30_) );
  DFF_X2 mem_reg_0__29_ ( .D(n1179), .CK(clk), .Q(mem_0__29_) );
  DFF_X2 mem_reg_0__28_ ( .D(n1178), .CK(clk), .Q(mem_0__28_) );
  DFF_X2 mem_reg_0__27_ ( .D(n1177), .CK(clk), .Q(mem_0__27_) );
  DFF_X2 mem_reg_0__26_ ( .D(n1176), .CK(clk), .Q(mem_0__26_) );
  DFF_X2 mem_reg_0__25_ ( .D(n1175), .CK(clk), .Q(mem_0__25_) );
  DFF_X2 mem_reg_0__24_ ( .D(n1174), .CK(clk), .Q(mem_0__24_) );
  DFF_X2 mem_reg_0__23_ ( .D(n1173), .CK(clk), .Q(mem_0__23_) );
  DFF_X2 mem_reg_0__22_ ( .D(n1172), .CK(clk), .Q(mem_0__22_) );
  DFF_X2 mem_reg_0__21_ ( .D(n1171), .CK(clk), .Q(mem_0__21_) );
  DFF_X2 mem_reg_0__20_ ( .D(n1170), .CK(clk), .Q(mem_0__20_) );
  DFF_X2 mem_reg_0__19_ ( .D(n1169), .CK(clk), .Q(mem_0__19_) );
  DFF_X2 mem_reg_0__18_ ( .D(n1168), .CK(clk), .Q(mem_0__18_) );
  DFF_X2 mem_reg_0__17_ ( .D(n1167), .CK(clk), .Q(mem_0__17_) );
  DFF_X2 mem_reg_0__16_ ( .D(n1166), .CK(clk), .Q(mem_0__16_) );
  DFF_X2 mem_reg_0__15_ ( .D(n1165), .CK(clk), .Q(mem_0__15_) );
  DFF_X2 mem_reg_0__14_ ( .D(n1164), .CK(clk), .Q(mem_0__14_) );
  DFF_X2 mem_reg_0__13_ ( .D(n1163), .CK(clk), .Q(mem_0__13_) );
  DFF_X2 mem_reg_0__12_ ( .D(n1162), .CK(clk), .Q(mem_0__12_) );
  DFF_X2 mem_reg_0__11_ ( .D(n1161), .CK(clk), .Q(mem_0__11_) );
  DFF_X2 mem_reg_0__10_ ( .D(n1160), .CK(clk), .Q(mem_0__10_) );
  DFF_X2 mem_reg_0__9_ ( .D(n1159), .CK(clk), .Q(mem_0__9_) );
  DFF_X2 mem_reg_0__8_ ( .D(n1158), .CK(clk), .Q(mem_0__8_) );
  DFF_X2 mem_reg_0__7_ ( .D(n1157), .CK(clk), .Q(mem_0__7_) );
  DFF_X2 mem_reg_0__6_ ( .D(n1156), .CK(clk), .Q(mem_0__6_) );
  DFF_X2 mem_reg_0__5_ ( .D(n1155), .CK(clk), .Q(mem_0__5_) );
  DFF_X2 mem_reg_0__4_ ( .D(n1154), .CK(clk), .Q(mem_0__4_) );
  DFF_X2 mem_reg_0__3_ ( .D(n1153), .CK(clk), .Q(mem_0__3_) );
  DFF_X2 mem_reg_0__2_ ( .D(n1152), .CK(clk), .Q(mem_0__2_) );
  DFF_X2 mem_reg_0__1_ ( .D(n1151), .CK(clk), .Q(mem_0__1_) );
  DFF_X2 mem_reg_0__0_ ( .D(n1150), .CK(clk), .Q(mem_0__0_) );
  INV_X4 U3 ( .A(clk), .ZN(n2238) );
  NAND2_X2 U7 ( .A1(mem_9__9_), .A2(n3058), .ZN(n7) );
  NAND2_X2 U9 ( .A1(mem_9__8_), .A2(n3057), .ZN(n9) );
  NAND2_X2 U11 ( .A1(mem_9__7_), .A2(n3057), .ZN(n11) );
  NAND2_X2 U13 ( .A1(mem_9__6_), .A2(n3057), .ZN(n13) );
  NAND2_X2 U15 ( .A1(mem_9__5_), .A2(n3058), .ZN(n15) );
  NAND2_X2 U17 ( .A1(mem_9__4_), .A2(n3057), .ZN(n17) );
  NAND2_X2 U19 ( .A1(mem_9__3_), .A2(n3056), .ZN(n19) );
  NAND2_X2 U21 ( .A1(mem_9__31_), .A2(n3056), .ZN(n21) );
  NAND2_X2 U23 ( .A1(mem_9__30_), .A2(n3058), .ZN(n23) );
  NAND2_X2 U25 ( .A1(mem_9__2_), .A2(n3058), .ZN(n25) );
  NAND2_X2 U27 ( .A1(mem_9__29_), .A2(n3058), .ZN(n27) );
  NAND2_X2 U29 ( .A1(mem_9__28_), .A2(n3056), .ZN(n29) );
  NAND2_X2 U31 ( .A1(mem_9__27_), .A2(n3058), .ZN(n31) );
  NAND2_X2 U33 ( .A1(mem_9__26_), .A2(n3056), .ZN(n33) );
  NAND2_X2 U35 ( .A1(mem_9__25_), .A2(n3058), .ZN(n35) );
  NAND2_X2 U37 ( .A1(mem_9__24_), .A2(n3056), .ZN(n37) );
  NAND2_X2 U39 ( .A1(mem_9__23_), .A2(n3058), .ZN(n39) );
  NAND2_X2 U41 ( .A1(mem_9__22_), .A2(n3057), .ZN(n41) );
  NAND2_X2 U43 ( .A1(mem_9__21_), .A2(n6), .ZN(n43) );
  NAND2_X2 U45 ( .A1(mem_9__20_), .A2(n6), .ZN(n45) );
  NAND2_X2 U47 ( .A1(mem_9__1_), .A2(n6), .ZN(n47) );
  NAND2_X2 U49 ( .A1(mem_9__19_), .A2(n6), .ZN(n49) );
  NAND2_X2 U51 ( .A1(mem_9__18_), .A2(n6), .ZN(n51) );
  NAND2_X2 U53 ( .A1(mem_9__17_), .A2(n6), .ZN(n53) );
  NAND2_X2 U55 ( .A1(mem_9__16_), .A2(n3058), .ZN(n55) );
  NAND2_X2 U57 ( .A1(mem_9__15_), .A2(n3058), .ZN(n57) );
  NAND2_X2 U59 ( .A1(mem_9__14_), .A2(n6), .ZN(n59) );
  NAND2_X2 U61 ( .A1(mem_9__13_), .A2(n3058), .ZN(n61) );
  NAND2_X2 U63 ( .A1(mem_9__12_), .A2(n3058), .ZN(n63) );
  NAND2_X2 U65 ( .A1(mem_9__11_), .A2(n6), .ZN(n65) );
  NAND2_X2 U67 ( .A1(mem_9__10_), .A2(n3058), .ZN(n67) );
  NAND2_X2 U69 ( .A1(mem_9__0_), .A2(n6), .ZN(n69) );
  NAND2_X2 U70 ( .A1(n70), .A2(n71), .ZN(n6) );
  NAND2_X2 U72 ( .A1(mem_8__9_), .A2(n3054), .ZN(n73) );
  NAND2_X2 U74 ( .A1(mem_8__8_), .A2(n3053), .ZN(n74) );
  NAND2_X2 U76 ( .A1(mem_8__7_), .A2(n3053), .ZN(n75) );
  NAND2_X2 U78 ( .A1(mem_8__6_), .A2(n3053), .ZN(n76) );
  NAND2_X2 U80 ( .A1(mem_8__5_), .A2(n3054), .ZN(n77) );
  NAND2_X2 U82 ( .A1(mem_8__4_), .A2(n3052), .ZN(n78) );
  NAND2_X2 U84 ( .A1(mem_8__3_), .A2(n3053), .ZN(n79) );
  NAND2_X2 U86 ( .A1(mem_8__31_), .A2(n3052), .ZN(n80) );
  NAND2_X2 U88 ( .A1(mem_8__30_), .A2(n3054), .ZN(n81) );
  NAND2_X2 U90 ( .A1(mem_8__2_), .A2(n72), .ZN(n82) );
  NAND2_X2 U92 ( .A1(mem_8__29_), .A2(n3054), .ZN(n83) );
  NAND2_X2 U94 ( .A1(mem_8__28_), .A2(n3054), .ZN(n84) );
  NAND2_X2 U96 ( .A1(mem_8__27_), .A2(n3052), .ZN(n85) );
  NAND2_X2 U98 ( .A1(mem_8__26_), .A2(n3054), .ZN(n86) );
  NAND2_X2 U100 ( .A1(mem_8__25_), .A2(n3052), .ZN(n87) );
  NAND2_X2 U102 ( .A1(mem_8__24_), .A2(n3054), .ZN(n88) );
  NAND2_X2 U104 ( .A1(mem_8__23_), .A2(n3052), .ZN(n89) );
  NAND2_X2 U106 ( .A1(mem_8__22_), .A2(n3054), .ZN(n90) );
  NAND2_X2 U108 ( .A1(mem_8__21_), .A2(n72), .ZN(n91) );
  NAND2_X2 U110 ( .A1(mem_8__20_), .A2(n72), .ZN(n92) );
  NAND2_X2 U112 ( .A1(mem_8__1_), .A2(n3053), .ZN(n93) );
  NAND2_X2 U114 ( .A1(mem_8__19_), .A2(n72), .ZN(n94) );
  NAND2_X2 U116 ( .A1(mem_8__18_), .A2(n72), .ZN(n95) );
  NAND2_X2 U118 ( .A1(mem_8__17_), .A2(n72), .ZN(n96) );
  NAND2_X2 U120 ( .A1(mem_8__16_), .A2(n3054), .ZN(n97) );
  NAND2_X2 U122 ( .A1(mem_8__15_), .A2(n3054), .ZN(n98) );
  NAND2_X2 U124 ( .A1(mem_8__14_), .A2(n72), .ZN(n99) );
  NAND2_X2 U126 ( .A1(mem_8__13_), .A2(n3054), .ZN(n100) );
  NAND2_X2 U128 ( .A1(mem_8__12_), .A2(n3054), .ZN(n101) );
  NAND2_X2 U130 ( .A1(mem_8__11_), .A2(n72), .ZN(n102) );
  NAND2_X2 U132 ( .A1(mem_8__10_), .A2(n3054), .ZN(n103) );
  NAND2_X2 U134 ( .A1(mem_8__0_), .A2(n72), .ZN(n104) );
  NAND2_X2 U135 ( .A1(n105), .A2(n71), .ZN(n72) );
  NAND2_X2 U137 ( .A1(mem_7__9_), .A2(n3050), .ZN(n107) );
  NAND2_X2 U139 ( .A1(mem_7__8_), .A2(n3049), .ZN(n108) );
  NAND2_X2 U141 ( .A1(mem_7__7_), .A2(n3049), .ZN(n109) );
  NAND2_X2 U143 ( .A1(mem_7__6_), .A2(n3049), .ZN(n110) );
  NAND2_X2 U145 ( .A1(mem_7__5_), .A2(n3048), .ZN(n111) );
  NAND2_X2 U147 ( .A1(mem_7__4_), .A2(n3049), .ZN(n112) );
  NAND2_X2 U149 ( .A1(mem_7__3_), .A2(n3048), .ZN(n113) );
  NAND2_X2 U151 ( .A1(mem_7__31_), .A2(n3048), .ZN(n114) );
  NAND2_X2 U153 ( .A1(mem_7__30_), .A2(n3050), .ZN(n115) );
  NAND2_X2 U155 ( .A1(mem_7__2_), .A2(n3050), .ZN(n116) );
  NAND2_X2 U157 ( .A1(mem_7__29_), .A2(n3050), .ZN(n117) );
  NAND2_X2 U159 ( .A1(mem_7__28_), .A2(n3050), .ZN(n118) );
  NAND2_X2 U161 ( .A1(mem_7__27_), .A2(n3050), .ZN(n119) );
  NAND2_X2 U163 ( .A1(mem_7__26_), .A2(n3050), .ZN(n120) );
  NAND2_X2 U165 ( .A1(mem_7__25_), .A2(n3050), .ZN(n121) );
  NAND2_X2 U167 ( .A1(mem_7__24_), .A2(n3050), .ZN(n122) );
  NAND2_X2 U169 ( .A1(mem_7__23_), .A2(n3050), .ZN(n123) );
  NAND2_X2 U171 ( .A1(mem_7__22_), .A2(n3050), .ZN(n124) );
  NAND2_X2 U173 ( .A1(mem_7__21_), .A2(n3050), .ZN(n125) );
  NAND2_X2 U175 ( .A1(mem_7__20_), .A2(n3050), .ZN(n126) );
  NAND2_X2 U177 ( .A1(mem_7__1_), .A2(n3050), .ZN(n127) );
  NAND2_X2 U179 ( .A1(mem_7__19_), .A2(n3050), .ZN(n128) );
  NAND2_X2 U181 ( .A1(mem_7__18_), .A2(n3050), .ZN(n129) );
  NAND2_X2 U183 ( .A1(mem_7__17_), .A2(n3050), .ZN(n130) );
  NAND2_X2 U185 ( .A1(mem_7__16_), .A2(n3050), .ZN(n131) );
  NAND2_X2 U187 ( .A1(mem_7__15_), .A2(n3050), .ZN(n132) );
  NAND2_X2 U189 ( .A1(mem_7__14_), .A2(n3050), .ZN(n133) );
  NAND2_X2 U191 ( .A1(mem_7__13_), .A2(n3050), .ZN(n134) );
  NAND2_X2 U193 ( .A1(mem_7__12_), .A2(n3050), .ZN(n135) );
  NAND2_X2 U195 ( .A1(mem_7__11_), .A2(n3050), .ZN(n136) );
  NAND2_X2 U197 ( .A1(mem_7__10_), .A2(n3050), .ZN(n137) );
  NAND2_X2 U199 ( .A1(mem_7__0_), .A2(n3050), .ZN(n138) );
  NAND2_X2 U202 ( .A1(mem_6__9_), .A2(n3047), .ZN(n142) );
  NAND2_X2 U204 ( .A1(mem_6__8_), .A2(n3046), .ZN(n143) );
  NAND2_X2 U206 ( .A1(mem_6__7_), .A2(n3046), .ZN(n144) );
  NAND2_X2 U208 ( .A1(mem_6__6_), .A2(n3045), .ZN(n145) );
  NAND2_X2 U210 ( .A1(mem_6__5_), .A2(n3046), .ZN(n146) );
  NAND2_X2 U212 ( .A1(mem_6__4_), .A2(n3045), .ZN(n147) );
  NAND2_X2 U214 ( .A1(mem_6__3_), .A2(n3046), .ZN(n148) );
  NAND2_X2 U216 ( .A1(mem_6__31_), .A2(n3045), .ZN(n149) );
  NAND2_X2 U218 ( .A1(mem_6__30_), .A2(n3047), .ZN(n150) );
  NAND2_X2 U220 ( .A1(mem_6__2_), .A2(n3047), .ZN(n151) );
  NAND2_X2 U222 ( .A1(mem_6__29_), .A2(n3047), .ZN(n152) );
  NAND2_X2 U224 ( .A1(mem_6__28_), .A2(n3047), .ZN(n153) );
  NAND2_X2 U226 ( .A1(mem_6__27_), .A2(n3047), .ZN(n154) );
  NAND2_X2 U228 ( .A1(mem_6__26_), .A2(n3047), .ZN(n155) );
  NAND2_X2 U230 ( .A1(mem_6__25_), .A2(n3047), .ZN(n156) );
  NAND2_X2 U232 ( .A1(mem_6__24_), .A2(n3047), .ZN(n157) );
  NAND2_X2 U234 ( .A1(mem_6__23_), .A2(n3047), .ZN(n158) );
  NAND2_X2 U236 ( .A1(mem_6__22_), .A2(n3047), .ZN(n159) );
  NAND2_X2 U238 ( .A1(mem_6__21_), .A2(n3047), .ZN(n160) );
  NAND2_X2 U240 ( .A1(mem_6__20_), .A2(n3047), .ZN(n161) );
  NAND2_X2 U242 ( .A1(mem_6__1_), .A2(n3047), .ZN(n162) );
  NAND2_X2 U244 ( .A1(mem_6__19_), .A2(n3047), .ZN(n163) );
  NAND2_X2 U246 ( .A1(mem_6__18_), .A2(n3047), .ZN(n164) );
  NAND2_X2 U248 ( .A1(mem_6__17_), .A2(n3047), .ZN(n165) );
  NAND2_X2 U250 ( .A1(mem_6__16_), .A2(n3047), .ZN(n166) );
  NAND2_X2 U252 ( .A1(mem_6__15_), .A2(n3047), .ZN(n167) );
  NAND2_X2 U254 ( .A1(mem_6__14_), .A2(n3047), .ZN(n168) );
  NAND2_X2 U256 ( .A1(mem_6__13_), .A2(n3047), .ZN(n169) );
  NAND2_X2 U258 ( .A1(mem_6__12_), .A2(n3047), .ZN(n170) );
  NAND2_X2 U260 ( .A1(mem_6__11_), .A2(n3047), .ZN(n171) );
  NAND2_X2 U262 ( .A1(mem_6__10_), .A2(n3047), .ZN(n172) );
  NAND2_X2 U264 ( .A1(mem_6__0_), .A2(n3047), .ZN(n173) );
  NAND2_X2 U267 ( .A1(mem_5__9_), .A2(n3044), .ZN(n176) );
  NAND2_X2 U269 ( .A1(mem_5__8_), .A2(n3043), .ZN(n177) );
  NAND2_X2 U271 ( .A1(mem_5__7_), .A2(n3043), .ZN(n178) );
  NAND2_X2 U273 ( .A1(mem_5__6_), .A2(n3043), .ZN(n179) );
  NAND2_X2 U275 ( .A1(mem_5__5_), .A2(n3042), .ZN(n180) );
  NAND2_X2 U277 ( .A1(mem_5__4_), .A2(n3043), .ZN(n181) );
  NAND2_X2 U279 ( .A1(mem_5__3_), .A2(n3042), .ZN(n182) );
  NAND2_X2 U281 ( .A1(mem_5__31_), .A2(n3042), .ZN(n183) );
  NAND2_X2 U283 ( .A1(mem_5__30_), .A2(n3044), .ZN(n184) );
  NAND2_X2 U285 ( .A1(mem_5__2_), .A2(n3044), .ZN(n185) );
  NAND2_X2 U287 ( .A1(mem_5__29_), .A2(n3044), .ZN(n186) );
  NAND2_X2 U289 ( .A1(mem_5__28_), .A2(n3044), .ZN(n187) );
  NAND2_X2 U291 ( .A1(mem_5__27_), .A2(n3044), .ZN(n188) );
  NAND2_X2 U293 ( .A1(mem_5__26_), .A2(n3044), .ZN(n189) );
  NAND2_X2 U295 ( .A1(mem_5__25_), .A2(n3044), .ZN(n190) );
  NAND2_X2 U297 ( .A1(mem_5__24_), .A2(n3044), .ZN(n191) );
  NAND2_X2 U299 ( .A1(mem_5__23_), .A2(n3044), .ZN(n192) );
  NAND2_X2 U301 ( .A1(mem_5__22_), .A2(n3044), .ZN(n193) );
  NAND2_X2 U303 ( .A1(mem_5__21_), .A2(n3044), .ZN(n194) );
  NAND2_X2 U305 ( .A1(mem_5__20_), .A2(n3044), .ZN(n195) );
  NAND2_X2 U307 ( .A1(mem_5__1_), .A2(n3044), .ZN(n196) );
  NAND2_X2 U309 ( .A1(mem_5__19_), .A2(n3044), .ZN(n197) );
  NAND2_X2 U311 ( .A1(mem_5__18_), .A2(n3044), .ZN(n198) );
  NAND2_X2 U313 ( .A1(mem_5__17_), .A2(n3044), .ZN(n199) );
  NAND2_X2 U315 ( .A1(mem_5__16_), .A2(n3044), .ZN(n200) );
  NAND2_X2 U317 ( .A1(mem_5__15_), .A2(n3044), .ZN(n201) );
  NAND2_X2 U319 ( .A1(mem_5__14_), .A2(n3044), .ZN(n202) );
  NAND2_X2 U321 ( .A1(mem_5__13_), .A2(n3044), .ZN(n203) );
  NAND2_X2 U323 ( .A1(mem_5__12_), .A2(n3044), .ZN(n204) );
  NAND2_X2 U325 ( .A1(mem_5__11_), .A2(n3044), .ZN(n205) );
  NAND2_X2 U327 ( .A1(mem_5__10_), .A2(n3044), .ZN(n206) );
  NAND2_X2 U329 ( .A1(mem_5__0_), .A2(n3044), .ZN(n207) );
  NAND2_X2 U332 ( .A1(mem_4__9_), .A2(n3041), .ZN(n209) );
  NAND2_X2 U334 ( .A1(mem_4__8_), .A2(n3040), .ZN(n210) );
  NAND2_X2 U336 ( .A1(mem_4__7_), .A2(n3040), .ZN(n211) );
  NAND2_X2 U338 ( .A1(mem_4__6_), .A2(n3039), .ZN(n212) );
  NAND2_X2 U340 ( .A1(mem_4__5_), .A2(n3040), .ZN(n213) );
  NAND2_X2 U342 ( .A1(mem_4__4_), .A2(n3039), .ZN(n214) );
  NAND2_X2 U344 ( .A1(mem_4__3_), .A2(n3040), .ZN(n215) );
  NAND2_X2 U346 ( .A1(mem_4__31_), .A2(n3039), .ZN(n216) );
  NAND2_X2 U348 ( .A1(mem_4__30_), .A2(n3041), .ZN(n217) );
  NAND2_X2 U350 ( .A1(mem_4__2_), .A2(n3041), .ZN(n218) );
  NAND2_X2 U352 ( .A1(mem_4__29_), .A2(n3041), .ZN(n219) );
  NAND2_X2 U354 ( .A1(mem_4__28_), .A2(n3041), .ZN(n220) );
  NAND2_X2 U356 ( .A1(mem_4__27_), .A2(n3041), .ZN(n221) );
  NAND2_X2 U358 ( .A1(mem_4__26_), .A2(n3041), .ZN(n222) );
  NAND2_X2 U360 ( .A1(mem_4__25_), .A2(n3041), .ZN(n223) );
  NAND2_X2 U362 ( .A1(mem_4__24_), .A2(n3041), .ZN(n224) );
  NAND2_X2 U364 ( .A1(mem_4__23_), .A2(n3041), .ZN(n225) );
  NAND2_X2 U366 ( .A1(mem_4__22_), .A2(n3041), .ZN(n226) );
  NAND2_X2 U368 ( .A1(mem_4__21_), .A2(n3041), .ZN(n227) );
  NAND2_X2 U370 ( .A1(mem_4__20_), .A2(n3041), .ZN(n228) );
  NAND2_X2 U372 ( .A1(mem_4__1_), .A2(n3041), .ZN(n229) );
  NAND2_X2 U374 ( .A1(mem_4__19_), .A2(n3041), .ZN(n230) );
  NAND2_X2 U376 ( .A1(mem_4__18_), .A2(n3041), .ZN(n231) );
  NAND2_X2 U378 ( .A1(mem_4__17_), .A2(n3041), .ZN(n232) );
  NAND2_X2 U380 ( .A1(mem_4__16_), .A2(n3041), .ZN(n233) );
  NAND2_X2 U382 ( .A1(mem_4__15_), .A2(n3041), .ZN(n234) );
  NAND2_X2 U384 ( .A1(mem_4__14_), .A2(n3041), .ZN(n235) );
  NAND2_X2 U386 ( .A1(mem_4__13_), .A2(n3041), .ZN(n236) );
  NAND2_X2 U388 ( .A1(mem_4__12_), .A2(n3041), .ZN(n237) );
  NAND2_X2 U390 ( .A1(mem_4__11_), .A2(n3041), .ZN(n238) );
  NAND2_X2 U392 ( .A1(mem_4__10_), .A2(n3041), .ZN(n239) );
  NAND2_X2 U394 ( .A1(mem_4__0_), .A2(n3041), .ZN(n240) );
  AND2_X2 U396 ( .A1(n241), .A2(n242), .ZN(n140) );
  NAND2_X2 U398 ( .A1(mem_3__9_), .A2(n3038), .ZN(n244) );
  NAND2_X2 U400 ( .A1(mem_3__8_), .A2(n3037), .ZN(n245) );
  NAND2_X2 U402 ( .A1(mem_3__7_), .A2(n3037), .ZN(n246) );
  NAND2_X2 U404 ( .A1(mem_3__6_), .A2(n3037), .ZN(n247) );
  NAND2_X2 U406 ( .A1(mem_3__5_), .A2(n3036), .ZN(n248) );
  NAND2_X2 U408 ( .A1(mem_3__4_), .A2(n3037), .ZN(n249) );
  NAND2_X2 U410 ( .A1(mem_3__3_), .A2(n3036), .ZN(n250) );
  NAND2_X2 U412 ( .A1(mem_3__31_), .A2(n3036), .ZN(n251) );
  NAND2_X2 U414 ( .A1(mem_3__30_), .A2(n3038), .ZN(n252) );
  NAND2_X2 U416 ( .A1(mem_3__2_), .A2(n3038), .ZN(n253) );
  NAND2_X2 U418 ( .A1(mem_3__29_), .A2(n3038), .ZN(n254) );
  NAND2_X2 U420 ( .A1(mem_3__28_), .A2(n3038), .ZN(n255) );
  NAND2_X2 U422 ( .A1(mem_3__27_), .A2(n3038), .ZN(n256) );
  NAND2_X2 U424 ( .A1(mem_3__26_), .A2(n3038), .ZN(n257) );
  NAND2_X2 U426 ( .A1(mem_3__25_), .A2(n3038), .ZN(n258) );
  NAND2_X2 U428 ( .A1(mem_3__24_), .A2(n3038), .ZN(n259) );
  NAND2_X2 U430 ( .A1(mem_3__23_), .A2(n3038), .ZN(n260) );
  NAND2_X2 U432 ( .A1(mem_3__22_), .A2(n3038), .ZN(n261) );
  NAND2_X2 U434 ( .A1(mem_3__21_), .A2(n3038), .ZN(n262) );
  NAND2_X2 U436 ( .A1(mem_3__20_), .A2(n3038), .ZN(n263) );
  NAND2_X2 U438 ( .A1(mem_3__1_), .A2(n3038), .ZN(n264) );
  NAND2_X2 U440 ( .A1(mem_3__19_), .A2(n3038), .ZN(n265) );
  NAND2_X2 U442 ( .A1(mem_3__18_), .A2(n3038), .ZN(n266) );
  NAND2_X2 U444 ( .A1(mem_3__17_), .A2(n3038), .ZN(n267) );
  NAND2_X2 U446 ( .A1(mem_3__16_), .A2(n3038), .ZN(n268) );
  NAND2_X2 U448 ( .A1(mem_3__15_), .A2(n3038), .ZN(n269) );
  NAND2_X2 U450 ( .A1(mem_3__14_), .A2(n3038), .ZN(n270) );
  NAND2_X2 U452 ( .A1(mem_3__13_), .A2(n3038), .ZN(n271) );
  NAND2_X2 U454 ( .A1(mem_3__12_), .A2(n3038), .ZN(n272) );
  NAND2_X2 U456 ( .A1(mem_3__11_), .A2(n3038), .ZN(n273) );
  NAND2_X2 U458 ( .A1(mem_3__10_), .A2(n3038), .ZN(n274) );
  NAND2_X2 U460 ( .A1(mem_3__0_), .A2(n3038), .ZN(n275) );
  NAND2_X2 U463 ( .A1(mem_31__9_), .A2(n3035), .ZN(n278) );
  NAND2_X2 U465 ( .A1(mem_31__8_), .A2(n3034), .ZN(n279) );
  NAND2_X2 U467 ( .A1(mem_31__7_), .A2(n3033), .ZN(n280) );
  NAND2_X2 U469 ( .A1(mem_31__6_), .A2(n3034), .ZN(n281) );
  NAND2_X2 U471 ( .A1(mem_31__5_), .A2(n3033), .ZN(n282) );
  NAND2_X2 U473 ( .A1(mem_31__4_), .A2(n3034), .ZN(n283) );
  NAND2_X2 U475 ( .A1(mem_31__3_), .A2(n3033), .ZN(n284) );
  NAND2_X2 U477 ( .A1(mem_31__31_), .A2(n3035), .ZN(n285) );
  NAND2_X2 U479 ( .A1(mem_31__30_), .A2(n3033), .ZN(n286) );
  NAND2_X2 U481 ( .A1(mem_31__2_), .A2(n3034), .ZN(n287) );
  NAND2_X2 U483 ( .A1(mem_31__29_), .A2(n277), .ZN(n288) );
  NAND2_X2 U497 ( .A1(mem_31__22_), .A2(n277), .ZN(n295) );
  NAND2_X2 U499 ( .A1(mem_31__21_), .A2(n277), .ZN(n296) );
  NAND2_X2 U501 ( .A1(mem_31__20_), .A2(n277), .ZN(n297) );
  NAND2_X2 U503 ( .A1(mem_31__1_), .A2(n277), .ZN(n298) );
  NAND2_X2 U505 ( .A1(mem_31__19_), .A2(n277), .ZN(n299) );
  NAND2_X2 U507 ( .A1(mem_31__18_), .A2(n277), .ZN(n300) );
  NAND2_X2 U509 ( .A1(mem_31__17_), .A2(n277), .ZN(n301) );
  NAND2_X2 U511 ( .A1(mem_31__16_), .A2(n3035), .ZN(n302) );
  NAND2_X2 U513 ( .A1(mem_31__15_), .A2(n3035), .ZN(n303) );
  NAND2_X2 U515 ( .A1(mem_31__14_), .A2(n277), .ZN(n304) );
  NAND2_X2 U517 ( .A1(mem_31__13_), .A2(n3035), .ZN(n305) );
  NAND2_X2 U519 ( .A1(mem_31__12_), .A2(n3035), .ZN(n306) );
  NAND2_X2 U521 ( .A1(mem_31__11_), .A2(n277), .ZN(n307) );
  NAND2_X2 U523 ( .A1(mem_31__10_), .A2(n3035), .ZN(n308) );
  NAND2_X2 U525 ( .A1(mem_31__0_), .A2(n277), .ZN(n309) );
  NAND2_X2 U526 ( .A1(n310), .A2(n139), .ZN(n277) );
  NAND2_X2 U528 ( .A1(mem_30__9_), .A2(n3031), .ZN(n312) );
  NAND2_X2 U530 ( .A1(mem_30__8_), .A2(n3030), .ZN(n313) );
  NAND2_X2 U532 ( .A1(mem_30__7_), .A2(n3029), .ZN(n314) );
  NAND2_X2 U534 ( .A1(mem_30__6_), .A2(n3030), .ZN(n315) );
  NAND2_X2 U536 ( .A1(mem_30__5_), .A2(n3029), .ZN(n316) );
  NAND2_X2 U538 ( .A1(mem_30__4_), .A2(n3030), .ZN(n317) );
  NAND2_X2 U540 ( .A1(mem_30__3_), .A2(n3029), .ZN(n318) );
  NAND2_X2 U542 ( .A1(mem_30__31_), .A2(n3031), .ZN(n319) );
  NAND2_X2 U544 ( .A1(mem_30__30_), .A2(n3031), .ZN(n320) );
  NAND2_X2 U546 ( .A1(mem_30__2_), .A2(n3031), .ZN(n321) );
  NAND2_X2 U548 ( .A1(mem_30__29_), .A2(n3031), .ZN(n322) );
  NAND2_X2 U550 ( .A1(mem_30__28_), .A2(n3031), .ZN(n323) );
  NAND2_X2 U552 ( .A1(mem_30__27_), .A2(n3029), .ZN(n324) );
  NAND2_X2 U556 ( .A1(mem_30__25_), .A2(n3030), .ZN(n326) );
  NAND2_X2 U558 ( .A1(mem_30__24_), .A2(n311), .ZN(n327) );
  NAND2_X2 U560 ( .A1(mem_30__23_), .A2(n311), .ZN(n328) );
  NAND2_X2 U562 ( .A1(mem_30__22_), .A2(n311), .ZN(n329) );
  NAND2_X2 U564 ( .A1(mem_30__21_), .A2(n311), .ZN(n330) );
  NAND2_X2 U566 ( .A1(mem_30__20_), .A2(n311), .ZN(n331) );
  NAND2_X2 U568 ( .A1(mem_30__1_), .A2(n311), .ZN(n332) );
  NAND2_X2 U570 ( .A1(mem_30__19_), .A2(n311), .ZN(n333) );
  NAND2_X2 U572 ( .A1(mem_30__18_), .A2(n311), .ZN(n334) );
  NAND2_X2 U574 ( .A1(mem_30__17_), .A2(n311), .ZN(n335) );
  NAND2_X2 U576 ( .A1(mem_30__16_), .A2(n3031), .ZN(n336) );
  NAND2_X2 U578 ( .A1(mem_30__15_), .A2(n3031), .ZN(n337) );
  NAND2_X2 U580 ( .A1(mem_30__14_), .A2(n311), .ZN(n338) );
  NAND2_X2 U582 ( .A1(mem_30__13_), .A2(n3031), .ZN(n339) );
  NAND2_X2 U584 ( .A1(mem_30__12_), .A2(n3031), .ZN(n340) );
  NAND2_X2 U586 ( .A1(mem_30__11_), .A2(n311), .ZN(n341) );
  NAND2_X2 U588 ( .A1(mem_30__10_), .A2(n3031), .ZN(n342) );
  NAND2_X2 U590 ( .A1(mem_30__0_), .A2(n311), .ZN(n343) );
  NAND2_X2 U591 ( .A1(n310), .A2(n174), .ZN(n311) );
  NAND2_X2 U593 ( .A1(mem_2__9_), .A2(n3027), .ZN(n345) );
  NAND2_X2 U595 ( .A1(mem_2__8_), .A2(n3026), .ZN(n346) );
  NAND2_X2 U597 ( .A1(mem_2__7_), .A2(n3026), .ZN(n347) );
  NAND2_X2 U599 ( .A1(mem_2__6_), .A2(n3025), .ZN(n348) );
  NAND2_X2 U601 ( .A1(mem_2__5_), .A2(n3026), .ZN(n349) );
  NAND2_X2 U603 ( .A1(mem_2__4_), .A2(n3025), .ZN(n350) );
  NAND2_X2 U605 ( .A1(mem_2__3_), .A2(n3026), .ZN(n351) );
  NAND2_X2 U607 ( .A1(mem_2__31_), .A2(n3025), .ZN(n352) );
  NAND2_X2 U609 ( .A1(mem_2__30_), .A2(n3027), .ZN(n353) );
  NAND2_X2 U611 ( .A1(mem_2__2_), .A2(n3027), .ZN(n354) );
  NAND2_X2 U613 ( .A1(mem_2__29_), .A2(n3027), .ZN(n355) );
  NAND2_X2 U615 ( .A1(mem_2__28_), .A2(n3027), .ZN(n356) );
  NAND2_X2 U617 ( .A1(mem_2__27_), .A2(n3027), .ZN(n357) );
  NAND2_X2 U619 ( .A1(mem_2__26_), .A2(n3027), .ZN(n358) );
  NAND2_X2 U621 ( .A1(mem_2__25_), .A2(n3027), .ZN(n359) );
  NAND2_X2 U623 ( .A1(mem_2__24_), .A2(n3027), .ZN(n360) );
  NAND2_X2 U625 ( .A1(mem_2__23_), .A2(n3027), .ZN(n361) );
  NAND2_X2 U627 ( .A1(mem_2__22_), .A2(n3027), .ZN(n362) );
  NAND2_X2 U629 ( .A1(mem_2__21_), .A2(n3027), .ZN(n363) );
  NAND2_X2 U631 ( .A1(mem_2__20_), .A2(n3027), .ZN(n364) );
  NAND2_X2 U633 ( .A1(mem_2__1_), .A2(n3027), .ZN(n365) );
  NAND2_X2 U635 ( .A1(mem_2__19_), .A2(n3027), .ZN(n366) );
  NAND2_X2 U637 ( .A1(mem_2__18_), .A2(n3027), .ZN(n367) );
  NAND2_X2 U639 ( .A1(mem_2__17_), .A2(n3027), .ZN(n368) );
  NAND2_X2 U641 ( .A1(mem_2__16_), .A2(n3027), .ZN(n369) );
  NAND2_X2 U643 ( .A1(mem_2__15_), .A2(n3027), .ZN(n370) );
  NAND2_X2 U645 ( .A1(mem_2__14_), .A2(n3027), .ZN(n371) );
  NAND2_X2 U647 ( .A1(mem_2__13_), .A2(n3027), .ZN(n372) );
  NAND2_X2 U649 ( .A1(mem_2__12_), .A2(n3027), .ZN(n373) );
  NAND2_X2 U651 ( .A1(mem_2__11_), .A2(n3027), .ZN(n374) );
  NAND2_X2 U653 ( .A1(mem_2__10_), .A2(n3027), .ZN(n375) );
  NAND2_X2 U655 ( .A1(mem_2__0_), .A2(n3027), .ZN(n376) );
  NAND2_X2 U658 ( .A1(mem_29__9_), .A2(n3023), .ZN(n378) );
  NAND2_X2 U660 ( .A1(mem_29__8_), .A2(n3021), .ZN(n379) );
  NAND2_X2 U662 ( .A1(mem_29__7_), .A2(n3022), .ZN(n380) );
  NAND2_X2 U664 ( .A1(mem_29__6_), .A2(n3021), .ZN(n381) );
  NAND2_X2 U666 ( .A1(mem_29__5_), .A2(n3022), .ZN(n382) );
  NAND2_X2 U668 ( .A1(mem_29__4_), .A2(n3021), .ZN(n383) );
  NAND2_X2 U670 ( .A1(mem_29__3_), .A2(n3022), .ZN(n384) );
  NAND2_X2 U672 ( .A1(mem_29__31_), .A2(n3023), .ZN(n385) );
  NAND2_X2 U674 ( .A1(mem_29__30_), .A2(n3023), .ZN(n386) );
  NAND2_X2 U676 ( .A1(mem_29__2_), .A2(n3023), .ZN(n387) );
  NAND2_X2 U678 ( .A1(mem_29__29_), .A2(n3023), .ZN(n388) );
  NAND2_X2 U680 ( .A1(mem_29__28_), .A2(n3022), .ZN(n389) );
  NAND2_X2 U682 ( .A1(mem_29__27_), .A2(n3021), .ZN(n390) );
  NAND2_X2 U684 ( .A1(mem_29__26_), .A2(n3023), .ZN(n391) );
  NAND2_X2 U686 ( .A1(mem_29__25_), .A2(n377), .ZN(n392) );
  NAND2_X2 U688 ( .A1(mem_29__24_), .A2(n377), .ZN(n393) );
  NAND2_X2 U690 ( .A1(mem_29__23_), .A2(n377), .ZN(n394) );
  NAND2_X2 U692 ( .A1(mem_29__22_), .A2(n377), .ZN(n395) );
  NAND2_X2 U694 ( .A1(mem_29__21_), .A2(n377), .ZN(n396) );
  NAND2_X2 U696 ( .A1(mem_29__20_), .A2(n377), .ZN(n397) );
  NAND2_X2 U698 ( .A1(mem_29__1_), .A2(n377), .ZN(n398) );
  NAND2_X2 U700 ( .A1(mem_29__19_), .A2(n377), .ZN(n399) );
  NAND2_X2 U702 ( .A1(mem_29__18_), .A2(n377), .ZN(n400) );
  NAND2_X2 U704 ( .A1(mem_29__17_), .A2(n377), .ZN(n401) );
  NAND2_X2 U706 ( .A1(mem_29__16_), .A2(n3023), .ZN(n402) );
  NAND2_X2 U708 ( .A1(mem_29__15_), .A2(n3023), .ZN(n403) );
  NAND2_X2 U710 ( .A1(mem_29__14_), .A2(n377), .ZN(n404) );
  NAND2_X2 U712 ( .A1(mem_29__13_), .A2(n3023), .ZN(n405) );
  NAND2_X2 U714 ( .A1(mem_29__12_), .A2(n3023), .ZN(n406) );
  NAND2_X2 U716 ( .A1(mem_29__11_), .A2(n377), .ZN(n407) );
  NAND2_X2 U718 ( .A1(mem_29__10_), .A2(n3023), .ZN(n408) );
  NAND2_X2 U720 ( .A1(mem_29__0_), .A2(n377), .ZN(n409) );
  NAND2_X2 U721 ( .A1(n310), .A2(n70), .ZN(n377) );
  NAND2_X2 U723 ( .A1(mem_28__9_), .A2(n3020), .ZN(n411) );
  NAND2_X2 U725 ( .A1(mem_28__8_), .A2(n3019), .ZN(n412) );
  NAND2_X2 U727 ( .A1(mem_28__7_), .A2(n3018), .ZN(n413) );
  NAND2_X2 U729 ( .A1(mem_28__6_), .A2(n3019), .ZN(n414) );
  NAND2_X2 U731 ( .A1(mem_28__5_), .A2(n3018), .ZN(n415) );
  NAND2_X2 U733 ( .A1(mem_28__4_), .A2(n3019), .ZN(n416) );
  NAND2_X2 U735 ( .A1(mem_28__3_), .A2(n3018), .ZN(n417) );
  NAND2_X2 U737 ( .A1(mem_28__31_), .A2(n3020), .ZN(n418) );
  NAND2_X2 U739 ( .A1(mem_28__30_), .A2(n3020), .ZN(n419) );
  NAND2_X2 U741 ( .A1(mem_28__2_), .A2(n3020), .ZN(n420) );
  NAND2_X2 U743 ( .A1(mem_28__29_), .A2(n3020), .ZN(n421) );
  NAND2_X2 U745 ( .A1(mem_28__28_), .A2(n3020), .ZN(n422) );
  NAND2_X2 U747 ( .A1(mem_28__27_), .A2(n3018), .ZN(n423) );
  NAND2_X2 U751 ( .A1(mem_28__25_), .A2(n3019), .ZN(n425) );
  NAND2_X2 U753 ( .A1(mem_28__24_), .A2(n410), .ZN(n426) );
  NAND2_X2 U755 ( .A1(mem_28__23_), .A2(n410), .ZN(n427) );
  NAND2_X2 U757 ( .A1(mem_28__22_), .A2(n410), .ZN(n428) );
  NAND2_X2 U759 ( .A1(mem_28__21_), .A2(n410), .ZN(n429) );
  NAND2_X2 U761 ( .A1(mem_28__20_), .A2(n410), .ZN(n430) );
  NAND2_X2 U763 ( .A1(mem_28__1_), .A2(n410), .ZN(n431) );
  NAND2_X2 U765 ( .A1(mem_28__19_), .A2(n410), .ZN(n432) );
  NAND2_X2 U767 ( .A1(mem_28__18_), .A2(n410), .ZN(n433) );
  NAND2_X2 U769 ( .A1(mem_28__17_), .A2(n410), .ZN(n434) );
  NAND2_X2 U771 ( .A1(mem_28__16_), .A2(n3020), .ZN(n435) );
  NAND2_X2 U773 ( .A1(mem_28__15_), .A2(n3020), .ZN(n436) );
  NAND2_X2 U775 ( .A1(mem_28__14_), .A2(n410), .ZN(n437) );
  NAND2_X2 U777 ( .A1(mem_28__13_), .A2(n3020), .ZN(n438) );
  NAND2_X2 U779 ( .A1(mem_28__12_), .A2(n3020), .ZN(n439) );
  NAND2_X2 U781 ( .A1(mem_28__11_), .A2(n410), .ZN(n440) );
  NAND2_X2 U783 ( .A1(mem_28__10_), .A2(n3020), .ZN(n441) );
  NAND2_X2 U785 ( .A1(mem_28__0_), .A2(n410), .ZN(n442) );
  NAND2_X2 U786 ( .A1(n310), .A2(n105), .ZN(n410) );
  AND2_X2 U787 ( .A1(n443), .A2(n444), .ZN(n310) );
  NAND2_X2 U789 ( .A1(mem_27__9_), .A2(n3015), .ZN(n446) );
  NAND2_X2 U791 ( .A1(mem_27__8_), .A2(n3014), .ZN(n447) );
  NAND2_X2 U793 ( .A1(mem_27__7_), .A2(n3015), .ZN(n448) );
  NAND2_X2 U795 ( .A1(mem_27__6_), .A2(n3014), .ZN(n449) );
  NAND2_X2 U797 ( .A1(mem_27__5_), .A2(n3015), .ZN(n450) );
  NAND2_X2 U799 ( .A1(mem_27__4_), .A2(n3014), .ZN(n451) );
  NAND2_X2 U801 ( .A1(mem_27__3_), .A2(n3015), .ZN(n452) );
  NAND2_X2 U803 ( .A1(mem_27__31_), .A2(n3016), .ZN(n453) );
  NAND2_X2 U805 ( .A1(mem_27__30_), .A2(n3016), .ZN(n454) );
  NAND2_X2 U807 ( .A1(mem_27__2_), .A2(n3016), .ZN(n455) );
  NAND2_X2 U809 ( .A1(mem_27__29_), .A2(n3016), .ZN(n456) );
  NAND2_X2 U811 ( .A1(mem_27__28_), .A2(n3016), .ZN(n457) );
  NAND2_X2 U813 ( .A1(mem_27__27_), .A2(n3016), .ZN(n458) );
  NAND2_X2 U815 ( .A1(mem_27__26_), .A2(n3016), .ZN(n459) );
  NAND2_X2 U817 ( .A1(mem_27__25_), .A2(n3016), .ZN(n460) );
  NAND2_X2 U819 ( .A1(mem_27__24_), .A2(n3016), .ZN(n461) );
  NAND2_X2 U821 ( .A1(mem_27__23_), .A2(n3016), .ZN(n462) );
  NAND2_X2 U823 ( .A1(mem_27__22_), .A2(n3016), .ZN(n463) );
  NAND2_X2 U825 ( .A1(mem_27__21_), .A2(n3016), .ZN(n464) );
  NAND2_X2 U827 ( .A1(mem_27__20_), .A2(n3016), .ZN(n465) );
  NAND2_X2 U829 ( .A1(mem_27__1_), .A2(n3016), .ZN(n466) );
  NAND2_X2 U831 ( .A1(mem_27__19_), .A2(n3016), .ZN(n467) );
  NAND2_X2 U833 ( .A1(mem_27__18_), .A2(n3016), .ZN(n468) );
  NAND2_X2 U835 ( .A1(mem_27__17_), .A2(n3016), .ZN(n469) );
  NAND2_X2 U837 ( .A1(mem_27__16_), .A2(n3016), .ZN(n470) );
  NAND2_X2 U839 ( .A1(mem_27__15_), .A2(n3016), .ZN(n471) );
  NAND2_X2 U841 ( .A1(mem_27__14_), .A2(n3016), .ZN(n472) );
  NAND2_X2 U843 ( .A1(mem_27__13_), .A2(n3016), .ZN(n473) );
  NAND2_X2 U845 ( .A1(mem_27__12_), .A2(n3016), .ZN(n474) );
  NAND2_X2 U847 ( .A1(mem_27__11_), .A2(n3016), .ZN(n475) );
  NAND2_X2 U849 ( .A1(mem_27__10_), .A2(n3016), .ZN(n476) );
  NAND2_X2 U851 ( .A1(mem_27__0_), .A2(n3016), .ZN(n477) );
  NAND2_X2 U852 ( .A1(n478), .A2(n139), .ZN(n445) );
  NAND2_X2 U854 ( .A1(mem_26__9_), .A2(n3012), .ZN(n480) );
  NAND2_X2 U856 ( .A1(mem_26__8_), .A2(n3011), .ZN(n481) );
  NAND2_X2 U858 ( .A1(mem_26__7_), .A2(n3010), .ZN(n482) );
  NAND2_X2 U860 ( .A1(mem_26__6_), .A2(n3011), .ZN(n483) );
  NAND2_X2 U862 ( .A1(mem_26__5_), .A2(n3010), .ZN(n484) );
  NAND2_X2 U864 ( .A1(mem_26__4_), .A2(n3011), .ZN(n485) );
  NAND2_X2 U866 ( .A1(mem_26__3_), .A2(n3010), .ZN(n486) );
  NAND2_X2 U870 ( .A1(mem_26__30_), .A2(n3011), .ZN(n488) );
  NAND2_X2 U872 ( .A1(mem_26__2_), .A2(n3012), .ZN(n489) );
  NAND2_X2 U874 ( .A1(mem_26__29_), .A2(n479), .ZN(n490) );
  NAND2_X2 U876 ( .A1(mem_26__28_), .A2(n479), .ZN(n491) );
  NAND2_X2 U878 ( .A1(mem_26__27_), .A2(n479), .ZN(n492) );
  NAND2_X2 U880 ( .A1(mem_26__26_), .A2(n479), .ZN(n493) );
  NAND2_X2 U882 ( .A1(mem_26__25_), .A2(n479), .ZN(n494) );
  NAND2_X2 U888 ( .A1(mem_26__22_), .A2(n479), .ZN(n497) );
  NAND2_X2 U890 ( .A1(mem_26__21_), .A2(n479), .ZN(n498) );
  NAND2_X2 U892 ( .A1(mem_26__20_), .A2(n479), .ZN(n499) );
  NAND2_X2 U894 ( .A1(mem_26__1_), .A2(n479), .ZN(n500) );
  NAND2_X2 U896 ( .A1(mem_26__19_), .A2(n479), .ZN(n501) );
  NAND2_X2 U898 ( .A1(mem_26__18_), .A2(n479), .ZN(n502) );
  NAND2_X2 U900 ( .A1(mem_26__17_), .A2(n479), .ZN(n503) );
  NAND2_X2 U902 ( .A1(mem_26__16_), .A2(n3012), .ZN(n504) );
  NAND2_X2 U904 ( .A1(mem_26__15_), .A2(n3012), .ZN(n505) );
  NAND2_X2 U906 ( .A1(mem_26__14_), .A2(n479), .ZN(n506) );
  NAND2_X2 U908 ( .A1(mem_26__13_), .A2(n3012), .ZN(n507) );
  NAND2_X2 U910 ( .A1(mem_26__12_), .A2(n3012), .ZN(n508) );
  NAND2_X2 U912 ( .A1(mem_26__11_), .A2(n479), .ZN(n509) );
  NAND2_X2 U914 ( .A1(mem_26__10_), .A2(n3012), .ZN(n510) );
  NAND2_X2 U916 ( .A1(mem_26__0_), .A2(n479), .ZN(n511) );
  NAND2_X2 U917 ( .A1(n478), .A2(n174), .ZN(n479) );
  NAND2_X2 U919 ( .A1(mem_25__9_), .A2(n3007), .ZN(n513) );
  NAND2_X2 U921 ( .A1(mem_25__8_), .A2(n3006), .ZN(n514) );
  NAND2_X2 U923 ( .A1(mem_25__7_), .A2(n3006), .ZN(n515) );
  NAND2_X2 U925 ( .A1(mem_25__6_), .A2(n3006), .ZN(n516) );
  NAND2_X2 U927 ( .A1(mem_25__5_), .A2(n3007), .ZN(n517) );
  NAND2_X2 U929 ( .A1(mem_25__4_), .A2(n3006), .ZN(n518) );
  NAND2_X2 U931 ( .A1(mem_25__3_), .A2(n3005), .ZN(n519) );
  NAND2_X2 U933 ( .A1(mem_25__31_), .A2(n3005), .ZN(n520) );
  NAND2_X2 U935 ( .A1(mem_25__30_), .A2(n3007), .ZN(n521) );
  NAND2_X2 U937 ( .A1(mem_25__2_), .A2(n3007), .ZN(n522) );
  NAND2_X2 U939 ( .A1(mem_25__29_), .A2(n3005), .ZN(n523) );
  NAND2_X2 U941 ( .A1(mem_25__28_), .A2(n3007), .ZN(n524) );
  NAND2_X2 U943 ( .A1(mem_25__27_), .A2(n3005), .ZN(n525) );
  NAND2_X2 U945 ( .A1(mem_25__26_), .A2(n3007), .ZN(n526) );
  NAND2_X2 U947 ( .A1(mem_25__25_), .A2(n3005), .ZN(n527) );
  NAND2_X2 U949 ( .A1(mem_25__24_), .A2(n3006), .ZN(n528) );
  NAND2_X2 U951 ( .A1(mem_25__23_), .A2(n3007), .ZN(n529) );
  NAND2_X2 U953 ( .A1(mem_25__22_), .A2(n512), .ZN(n530) );
  NAND2_X2 U955 ( .A1(mem_25__21_), .A2(n512), .ZN(n531) );
  NAND2_X2 U957 ( .A1(mem_25__20_), .A2(n512), .ZN(n532) );
  NAND2_X2 U959 ( .A1(mem_25__1_), .A2(n512), .ZN(n533) );
  NAND2_X2 U961 ( .A1(mem_25__19_), .A2(n512), .ZN(n534) );
  NAND2_X2 U963 ( .A1(mem_25__18_), .A2(n512), .ZN(n535) );
  NAND2_X2 U965 ( .A1(mem_25__17_), .A2(n512), .ZN(n536) );
  NAND2_X2 U967 ( .A1(mem_25__16_), .A2(n3007), .ZN(n537) );
  NAND2_X2 U969 ( .A1(mem_25__15_), .A2(n3007), .ZN(n538) );
  NAND2_X2 U971 ( .A1(mem_25__14_), .A2(n512), .ZN(n539) );
  NAND2_X2 U973 ( .A1(mem_25__13_), .A2(n3007), .ZN(n540) );
  NAND2_X2 U975 ( .A1(mem_25__12_), .A2(n3007), .ZN(n541) );
  NAND2_X2 U977 ( .A1(mem_25__11_), .A2(n512), .ZN(n542) );
  NAND2_X2 U979 ( .A1(mem_25__10_), .A2(n3007), .ZN(n543) );
  NAND2_X2 U981 ( .A1(mem_25__0_), .A2(n512), .ZN(n544) );
  NAND2_X2 U982 ( .A1(n478), .A2(n70), .ZN(n512) );
  NAND2_X2 U984 ( .A1(mem_24__9_), .A2(n3003), .ZN(n546) );
  NAND2_X2 U986 ( .A1(mem_24__8_), .A2(n3002), .ZN(n547) );
  NAND2_X2 U988 ( .A1(mem_24__7_), .A2(n3002), .ZN(n548) );
  NAND2_X2 U990 ( .A1(mem_24__6_), .A2(n3002), .ZN(n549) );
  NAND2_X2 U992 ( .A1(mem_24__5_), .A2(n3003), .ZN(n550) );
  NAND2_X2 U994 ( .A1(mem_24__4_), .A2(n3001), .ZN(n551) );
  NAND2_X2 U996 ( .A1(mem_24__3_), .A2(n3002), .ZN(n552) );
  NAND2_X2 U998 ( .A1(mem_24__31_), .A2(n3001), .ZN(n553) );
  NAND2_X2 U1000 ( .A1(mem_24__30_), .A2(n3003), .ZN(n554) );
  NAND2_X2 U1002 ( .A1(mem_24__2_), .A2(n3003), .ZN(n555) );
  NAND2_X2 U1004 ( .A1(mem_24__29_), .A2(n3001), .ZN(n556) );
  NAND2_X2 U1006 ( .A1(mem_24__28_), .A2(n3003), .ZN(n557) );
  NAND2_X2 U1008 ( .A1(mem_24__27_), .A2(n3001), .ZN(n558) );
  NAND2_X2 U1010 ( .A1(mem_24__26_), .A2(n3003), .ZN(n559) );
  NAND2_X2 U1012 ( .A1(mem_24__25_), .A2(n3001), .ZN(n560) );
  NAND2_X2 U1014 ( .A1(mem_24__24_), .A2(n3002), .ZN(n561) );
  NAND2_X2 U1016 ( .A1(mem_24__23_), .A2(n3003), .ZN(n562) );
  NAND2_X2 U1018 ( .A1(mem_24__22_), .A2(n545), .ZN(n563) );
  NAND2_X2 U1020 ( .A1(mem_24__21_), .A2(n545), .ZN(n564) );
  NAND2_X2 U1022 ( .A1(mem_24__20_), .A2(n545), .ZN(n565) );
  NAND2_X2 U1024 ( .A1(mem_24__1_), .A2(n545), .ZN(n566) );
  NAND2_X2 U1026 ( .A1(mem_24__19_), .A2(n545), .ZN(n567) );
  NAND2_X2 U1028 ( .A1(mem_24__18_), .A2(n545), .ZN(n568) );
  NAND2_X2 U1030 ( .A1(mem_24__17_), .A2(n545), .ZN(n569) );
  NAND2_X2 U1032 ( .A1(mem_24__16_), .A2(n3003), .ZN(n570) );
  NAND2_X2 U1034 ( .A1(mem_24__15_), .A2(n3003), .ZN(n571) );
  NAND2_X2 U1036 ( .A1(mem_24__14_), .A2(n545), .ZN(n572) );
  NAND2_X2 U1038 ( .A1(mem_24__13_), .A2(n3003), .ZN(n573) );
  NAND2_X2 U1040 ( .A1(mem_24__12_), .A2(n3003), .ZN(n574) );
  NAND2_X2 U1042 ( .A1(mem_24__11_), .A2(n545), .ZN(n575) );
  NAND2_X2 U1044 ( .A1(mem_24__10_), .A2(n3003), .ZN(n576) );
  NAND2_X2 U1046 ( .A1(mem_24__0_), .A2(n545), .ZN(n577) );
  NAND2_X2 U1047 ( .A1(n478), .A2(n105), .ZN(n545) );
  AND2_X2 U1048 ( .A1(n443), .A2(n578), .ZN(n478) );
  NAND2_X2 U1050 ( .A1(mem_23__9_), .A2(n3000), .ZN(n580) );
  NAND2_X2 U1052 ( .A1(mem_23__8_), .A2(n2999), .ZN(n581) );
  NAND2_X2 U1054 ( .A1(mem_23__7_), .A2(n2998), .ZN(n582) );
  NAND2_X2 U1056 ( .A1(mem_23__6_), .A2(n2999), .ZN(n583) );
  NAND2_X2 U1058 ( .A1(mem_23__5_), .A2(n2998), .ZN(n584) );
  NAND2_X2 U1060 ( .A1(mem_23__4_), .A2(n2999), .ZN(n585) );
  NAND2_X2 U1062 ( .A1(mem_23__3_), .A2(n2998), .ZN(n586) );
  NAND2_X2 U1068 ( .A1(mem_23__2_), .A2(n579), .ZN(n589) );
  NAND2_X2 U1084 ( .A1(mem_23__22_), .A2(n579), .ZN(n597) );
  NAND2_X2 U1086 ( .A1(mem_23__21_), .A2(n579), .ZN(n598) );
  NAND2_X2 U1088 ( .A1(mem_23__20_), .A2(n579), .ZN(n599) );
  NAND2_X2 U1090 ( .A1(mem_23__1_), .A2(n579), .ZN(n600) );
  NAND2_X2 U1092 ( .A1(mem_23__19_), .A2(n579), .ZN(n601) );
  NAND2_X2 U1094 ( .A1(mem_23__18_), .A2(n579), .ZN(n602) );
  NAND2_X2 U1096 ( .A1(mem_23__17_), .A2(n579), .ZN(n603) );
  NAND2_X2 U1098 ( .A1(mem_23__16_), .A2(n3000), .ZN(n604) );
  NAND2_X2 U1100 ( .A1(mem_23__15_), .A2(n3000), .ZN(n605) );
  NAND2_X2 U1102 ( .A1(mem_23__14_), .A2(n579), .ZN(n606) );
  NAND2_X2 U1104 ( .A1(mem_23__13_), .A2(n3000), .ZN(n607) );
  NAND2_X2 U1106 ( .A1(mem_23__12_), .A2(n3000), .ZN(n608) );
  NAND2_X2 U1108 ( .A1(mem_23__11_), .A2(n579), .ZN(n609) );
  NAND2_X2 U1110 ( .A1(mem_23__10_), .A2(n3000), .ZN(n610) );
  NAND2_X2 U1112 ( .A1(mem_23__0_), .A2(n579), .ZN(n611) );
  NAND2_X2 U1113 ( .A1(n612), .A2(n139), .ZN(n579) );
  NAND2_X2 U1115 ( .A1(mem_22__9_), .A2(n2996), .ZN(n614) );
  NAND2_X2 U1117 ( .A1(mem_22__8_), .A2(n2994), .ZN(n615) );
  NAND2_X2 U1119 ( .A1(mem_22__7_), .A2(n2994), .ZN(n616) );
  NAND2_X2 U1121 ( .A1(mem_22__6_), .A2(n2995), .ZN(n617) );
  NAND2_X2 U1123 ( .A1(mem_22__5_), .A2(n2994), .ZN(n618) );
  NAND2_X2 U1125 ( .A1(mem_22__4_), .A2(n2996), .ZN(n619) );
  NAND2_X2 U1127 ( .A1(mem_22__3_), .A2(n2995), .ZN(n620) );
  NAND2_X2 U1129 ( .A1(mem_22__31_), .A2(n2995), .ZN(n621) );
  NAND2_X2 U1131 ( .A1(mem_22__30_), .A2(n2996), .ZN(n622) );
  NAND2_X2 U1133 ( .A1(mem_22__2_), .A2(n2996), .ZN(n623) );
  NAND2_X2 U1135 ( .A1(mem_22__29_), .A2(n2996), .ZN(n624) );
  NAND2_X2 U1137 ( .A1(mem_22__28_), .A2(n2996), .ZN(n625) );
  NAND2_X2 U1139 ( .A1(mem_22__27_), .A2(n2994), .ZN(n626) );
  NAND2_X2 U1143 ( .A1(mem_22__25_), .A2(n2995), .ZN(n628) );
  NAND2_X2 U1145 ( .A1(mem_22__24_), .A2(n613), .ZN(n629) );
  NAND2_X2 U1147 ( .A1(mem_22__23_), .A2(n613), .ZN(n630) );
  NAND2_X2 U1149 ( .A1(mem_22__22_), .A2(n613), .ZN(n631) );
  NAND2_X2 U1151 ( .A1(mem_22__21_), .A2(n613), .ZN(n632) );
  NAND2_X2 U1153 ( .A1(mem_22__20_), .A2(n613), .ZN(n633) );
  NAND2_X2 U1155 ( .A1(mem_22__1_), .A2(n613), .ZN(n634) );
  NAND2_X2 U1157 ( .A1(mem_22__19_), .A2(n613), .ZN(n635) );
  NAND2_X2 U1159 ( .A1(mem_22__18_), .A2(n613), .ZN(n636) );
  NAND2_X2 U1161 ( .A1(mem_22__17_), .A2(n613), .ZN(n637) );
  NAND2_X2 U1163 ( .A1(mem_22__16_), .A2(n2996), .ZN(n638) );
  NAND2_X2 U1165 ( .A1(mem_22__15_), .A2(n2996), .ZN(n639) );
  NAND2_X2 U1167 ( .A1(mem_22__14_), .A2(n613), .ZN(n640) );
  NAND2_X2 U1169 ( .A1(mem_22__13_), .A2(n2996), .ZN(n641) );
  NAND2_X2 U1171 ( .A1(mem_22__12_), .A2(n2996), .ZN(n642) );
  NAND2_X2 U1173 ( .A1(mem_22__11_), .A2(n613), .ZN(n643) );
  NAND2_X2 U1175 ( .A1(mem_22__10_), .A2(n2996), .ZN(n644) );
  NAND2_X2 U1177 ( .A1(mem_22__0_), .A2(n613), .ZN(n645) );
  NAND2_X2 U1178 ( .A1(n612), .A2(n174), .ZN(n613) );
  NAND2_X2 U1180 ( .A1(mem_21__9_), .A2(n2991), .ZN(n647) );
  NAND2_X2 U1182 ( .A1(mem_21__8_), .A2(n2990), .ZN(n648) );
  NAND2_X2 U1184 ( .A1(mem_21__7_), .A2(n2990), .ZN(n649) );
  NAND2_X2 U1186 ( .A1(mem_21__6_), .A2(n2990), .ZN(n650) );
  NAND2_X2 U1188 ( .A1(mem_21__5_), .A2(n2989), .ZN(n651) );
  NAND2_X2 U1190 ( .A1(mem_21__4_), .A2(n2991), .ZN(n652) );
  NAND2_X2 U1192 ( .A1(mem_21__3_), .A2(n2990), .ZN(n653) );
  NAND2_X2 U1194 ( .A1(mem_21__31_), .A2(n2989), .ZN(n654) );
  NAND2_X2 U1196 ( .A1(mem_21__30_), .A2(n2991), .ZN(n655) );
  NAND2_X2 U1198 ( .A1(mem_21__2_), .A2(n2991), .ZN(n656) );
  NAND2_X2 U1200 ( .A1(mem_21__29_), .A2(n2989), .ZN(n657) );
  NAND2_X2 U1202 ( .A1(mem_21__28_), .A2(n2991), .ZN(n658) );
  NAND2_X2 U1204 ( .A1(mem_21__27_), .A2(n2989), .ZN(n659) );
  NAND2_X2 U1206 ( .A1(mem_21__26_), .A2(n2991), .ZN(n660) );
  NAND2_X2 U1208 ( .A1(mem_21__25_), .A2(n2989), .ZN(n661) );
  NAND2_X2 U1210 ( .A1(mem_21__24_), .A2(n2990), .ZN(n662) );
  NAND2_X2 U1212 ( .A1(mem_21__23_), .A2(n2991), .ZN(n663) );
  NAND2_X2 U1214 ( .A1(mem_21__22_), .A2(n646), .ZN(n664) );
  NAND2_X2 U1216 ( .A1(mem_21__21_), .A2(n646), .ZN(n665) );
  NAND2_X2 U1218 ( .A1(mem_21__20_), .A2(n646), .ZN(n666) );
  NAND2_X2 U1220 ( .A1(mem_21__1_), .A2(n646), .ZN(n667) );
  NAND2_X2 U1222 ( .A1(mem_21__19_), .A2(n646), .ZN(n668) );
  NAND2_X2 U1224 ( .A1(mem_21__18_), .A2(n646), .ZN(n669) );
  NAND2_X2 U1226 ( .A1(mem_21__17_), .A2(n646), .ZN(n670) );
  NAND2_X2 U1228 ( .A1(mem_21__16_), .A2(n2991), .ZN(n671) );
  NAND2_X2 U1230 ( .A1(mem_21__15_), .A2(n2991), .ZN(n672) );
  NAND2_X2 U1232 ( .A1(mem_21__14_), .A2(n646), .ZN(n673) );
  NAND2_X2 U1234 ( .A1(mem_21__13_), .A2(n2991), .ZN(n674) );
  NAND2_X2 U1236 ( .A1(mem_21__12_), .A2(n2991), .ZN(n675) );
  NAND2_X2 U1238 ( .A1(mem_21__11_), .A2(n646), .ZN(n676) );
  NAND2_X2 U1240 ( .A1(mem_21__10_), .A2(n2991), .ZN(n677) );
  NAND2_X2 U1242 ( .A1(mem_21__0_), .A2(n646), .ZN(n678) );
  NAND2_X2 U1243 ( .A1(n612), .A2(n70), .ZN(n646) );
  NAND2_X2 U1245 ( .A1(mem_20__9_), .A2(n2987), .ZN(n680) );
  NAND2_X2 U1247 ( .A1(mem_20__8_), .A2(n2986), .ZN(n681) );
  NAND2_X2 U1249 ( .A1(mem_20__7_), .A2(n2986), .ZN(n682) );
  NAND2_X2 U1251 ( .A1(mem_20__6_), .A2(n2985), .ZN(n683) );
  NAND2_X2 U1253 ( .A1(mem_20__5_), .A2(n2986), .ZN(n684) );
  NAND2_X2 U1255 ( .A1(mem_20__4_), .A2(n2987), .ZN(n685) );
  NAND2_X2 U1257 ( .A1(mem_20__3_), .A2(n2985), .ZN(n686) );
  NAND2_X2 U1259 ( .A1(mem_20__31_), .A2(n2985), .ZN(n687) );
  NAND2_X2 U1261 ( .A1(mem_20__30_), .A2(n2987), .ZN(n688) );
  NAND2_X2 U1263 ( .A1(mem_20__2_), .A2(n2987), .ZN(n689) );
  NAND2_X2 U1265 ( .A1(mem_20__29_), .A2(n2987), .ZN(n690) );
  NAND2_X2 U1267 ( .A1(mem_20__28_), .A2(n2986), .ZN(n691) );
  NAND2_X2 U1269 ( .A1(mem_20__27_), .A2(n2985), .ZN(n692) );
  NAND2_X2 U1271 ( .A1(mem_20__26_), .A2(n2987), .ZN(n693) );
  NAND2_X2 U1273 ( .A1(mem_20__25_), .A2(n679), .ZN(n694) );
  NAND2_X2 U1275 ( .A1(mem_20__24_), .A2(n679), .ZN(n695) );
  NAND2_X2 U1277 ( .A1(mem_20__23_), .A2(n679), .ZN(n696) );
  NAND2_X2 U1279 ( .A1(mem_20__22_), .A2(n679), .ZN(n697) );
  NAND2_X2 U1281 ( .A1(mem_20__21_), .A2(n679), .ZN(n698) );
  NAND2_X2 U1283 ( .A1(mem_20__20_), .A2(n679), .ZN(n699) );
  NAND2_X2 U1285 ( .A1(mem_20__1_), .A2(n679), .ZN(n700) );
  NAND2_X2 U1287 ( .A1(mem_20__19_), .A2(n679), .ZN(n701) );
  NAND2_X2 U1289 ( .A1(mem_20__18_), .A2(n679), .ZN(n702) );
  NAND2_X2 U1291 ( .A1(mem_20__17_), .A2(n679), .ZN(n703) );
  NAND2_X2 U1293 ( .A1(mem_20__16_), .A2(n2987), .ZN(n704) );
  NAND2_X2 U1295 ( .A1(mem_20__15_), .A2(n2987), .ZN(n705) );
  NAND2_X2 U1297 ( .A1(mem_20__14_), .A2(n679), .ZN(n706) );
  NAND2_X2 U1299 ( .A1(mem_20__13_), .A2(n2987), .ZN(n707) );
  NAND2_X2 U1301 ( .A1(mem_20__12_), .A2(n2987), .ZN(n708) );
  NAND2_X2 U1303 ( .A1(mem_20__11_), .A2(n679), .ZN(n709) );
  NAND2_X2 U1305 ( .A1(mem_20__10_), .A2(n2987), .ZN(n710) );
  NAND2_X2 U1307 ( .A1(mem_20__0_), .A2(n679), .ZN(n711) );
  NAND2_X2 U1308 ( .A1(n612), .A2(n105), .ZN(n679) );
  AND2_X2 U1309 ( .A1(n443), .A2(n241), .ZN(n612) );
  NAND2_X2 U1312 ( .A1(mem_1__9_), .A2(n2984), .ZN(n714) );
  NAND2_X2 U1314 ( .A1(mem_1__8_), .A2(n2983), .ZN(n715) );
  NAND2_X2 U1316 ( .A1(mem_1__7_), .A2(n2983), .ZN(n716) );
  NAND2_X2 U1318 ( .A1(mem_1__6_), .A2(n2983), .ZN(n717) );
  NAND2_X2 U1320 ( .A1(mem_1__5_), .A2(n2983), .ZN(n718) );
  NAND2_X2 U1322 ( .A1(mem_1__4_), .A2(n2982), .ZN(n719) );
  NAND2_X2 U1324 ( .A1(mem_1__3_), .A2(n2983), .ZN(n720) );
  NAND2_X2 U1326 ( .A1(mem_1__31_), .A2(n2982), .ZN(n721) );
  NAND2_X2 U1328 ( .A1(mem_1__30_), .A2(n2984), .ZN(n722) );
  NAND2_X2 U1330 ( .A1(mem_1__2_), .A2(n2984), .ZN(n723) );
  NAND2_X2 U1332 ( .A1(mem_1__29_), .A2(n2984), .ZN(n724) );
  NAND2_X2 U1334 ( .A1(mem_1__28_), .A2(n2984), .ZN(n725) );
  NAND2_X2 U1336 ( .A1(mem_1__27_), .A2(n2984), .ZN(n726) );
  NAND2_X2 U1338 ( .A1(mem_1__26_), .A2(n2984), .ZN(n727) );
  NAND2_X2 U1340 ( .A1(mem_1__25_), .A2(n2984), .ZN(n728) );
  NAND2_X2 U1342 ( .A1(mem_1__24_), .A2(n2984), .ZN(n729) );
  NAND2_X2 U1344 ( .A1(mem_1__23_), .A2(n2984), .ZN(n730) );
  NAND2_X2 U1346 ( .A1(mem_1__22_), .A2(n2984), .ZN(n731) );
  NAND2_X2 U1348 ( .A1(mem_1__21_), .A2(n2984), .ZN(n732) );
  NAND2_X2 U1350 ( .A1(mem_1__20_), .A2(n2984), .ZN(n733) );
  NAND2_X2 U1352 ( .A1(mem_1__1_), .A2(n2984), .ZN(n734) );
  NAND2_X2 U1354 ( .A1(mem_1__19_), .A2(n2984), .ZN(n735) );
  NAND2_X2 U1356 ( .A1(mem_1__18_), .A2(n2984), .ZN(n736) );
  NAND2_X2 U1358 ( .A1(mem_1__17_), .A2(n2984), .ZN(n737) );
  NAND2_X2 U1360 ( .A1(mem_1__16_), .A2(n2984), .ZN(n738) );
  NAND2_X2 U1362 ( .A1(mem_1__15_), .A2(n2984), .ZN(n739) );
  NAND2_X2 U1364 ( .A1(mem_1__14_), .A2(n2984), .ZN(n740) );
  NAND2_X2 U1366 ( .A1(mem_1__13_), .A2(n2984), .ZN(n741) );
  NAND2_X2 U1368 ( .A1(mem_1__12_), .A2(n2984), .ZN(n742) );
  NAND2_X2 U1370 ( .A1(mem_1__11_), .A2(n2984), .ZN(n743) );
  NAND2_X2 U1372 ( .A1(mem_1__10_), .A2(n2984), .ZN(n744) );
  NAND2_X2 U1374 ( .A1(mem_1__0_), .A2(n2984), .ZN(n745) );
  AND2_X2 U1376 ( .A1(n746), .A2(n242), .ZN(n276) );
  NAND2_X2 U1378 ( .A1(mem_19__9_), .A2(n2981), .ZN(n748) );
  NAND2_X2 U1380 ( .A1(mem_19__8_), .A2(n2980), .ZN(n749) );
  NAND2_X2 U1382 ( .A1(mem_19__7_), .A2(n2979), .ZN(n750) );
  NAND2_X2 U1384 ( .A1(mem_19__6_), .A2(n2980), .ZN(n751) );
  NAND2_X2 U1386 ( .A1(mem_19__5_), .A2(n2979), .ZN(n752) );
  NAND2_X2 U1388 ( .A1(mem_19__4_), .A2(n2980), .ZN(n753) );
  NAND2_X2 U1390 ( .A1(mem_19__3_), .A2(n2979), .ZN(n754) );
  NAND2_X2 U1396 ( .A1(mem_19__2_), .A2(n747), .ZN(n757) );
  NAND2_X2 U1412 ( .A1(mem_19__22_), .A2(n747), .ZN(n765) );
  NAND2_X2 U1414 ( .A1(mem_19__21_), .A2(n747), .ZN(n766) );
  NAND2_X2 U1416 ( .A1(mem_19__20_), .A2(n747), .ZN(n767) );
  NAND2_X2 U1418 ( .A1(mem_19__1_), .A2(n747), .ZN(n768) );
  NAND2_X2 U1420 ( .A1(mem_19__19_), .A2(n747), .ZN(n769) );
  NAND2_X2 U1422 ( .A1(mem_19__18_), .A2(n747), .ZN(n770) );
  NAND2_X2 U1424 ( .A1(mem_19__17_), .A2(n747), .ZN(n771) );
  NAND2_X2 U1426 ( .A1(mem_19__16_), .A2(n2981), .ZN(n772) );
  NAND2_X2 U1428 ( .A1(mem_19__15_), .A2(n2981), .ZN(n773) );
  NAND2_X2 U1430 ( .A1(mem_19__14_), .A2(n747), .ZN(n774) );
  NAND2_X2 U1432 ( .A1(mem_19__13_), .A2(n2981), .ZN(n775) );
  NAND2_X2 U1434 ( .A1(mem_19__12_), .A2(n2981), .ZN(n776) );
  NAND2_X2 U1436 ( .A1(mem_19__11_), .A2(n747), .ZN(n777) );
  NAND2_X2 U1438 ( .A1(mem_19__10_), .A2(n2981), .ZN(n778) );
  NAND2_X2 U1440 ( .A1(mem_19__0_), .A2(n747), .ZN(n779) );
  NAND2_X2 U1441 ( .A1(n780), .A2(n139), .ZN(n747) );
  NAND2_X2 U1443 ( .A1(mem_18__9_), .A2(n2977), .ZN(n782) );
  NAND2_X2 U1445 ( .A1(mem_18__8_), .A2(n2976), .ZN(n783) );
  NAND2_X2 U1447 ( .A1(mem_18__7_), .A2(n2975), .ZN(n784) );
  NAND2_X2 U1449 ( .A1(mem_18__6_), .A2(n2976), .ZN(n785) );
  NAND2_X2 U1451 ( .A1(mem_18__5_), .A2(n2975), .ZN(n786) );
  NAND2_X2 U1453 ( .A1(mem_18__4_), .A2(n2976), .ZN(n787) );
  NAND2_X2 U1455 ( .A1(mem_18__3_), .A2(n2975), .ZN(n788) );
  NAND2_X2 U1461 ( .A1(mem_18__2_), .A2(n781), .ZN(n791) );
  NAND2_X2 U1463 ( .A1(mem_18__29_), .A2(n781), .ZN(n792) );
  NAND2_X2 U1465 ( .A1(mem_18__28_), .A2(n781), .ZN(n793) );
  NAND2_X2 U1469 ( .A1(mem_18__26_), .A2(n781), .ZN(n795) );
  NAND2_X2 U1471 ( .A1(mem_18__25_), .A2(n781), .ZN(n796) );
  NAND2_X2 U1477 ( .A1(mem_18__22_), .A2(n781), .ZN(n799) );
  NAND2_X2 U1479 ( .A1(mem_18__21_), .A2(n781), .ZN(n800) );
  NAND2_X2 U1481 ( .A1(mem_18__20_), .A2(n781), .ZN(n801) );
  NAND2_X2 U1483 ( .A1(mem_18__1_), .A2(n781), .ZN(n802) );
  NAND2_X2 U1485 ( .A1(mem_18__19_), .A2(n781), .ZN(n803) );
  NAND2_X2 U1487 ( .A1(mem_18__18_), .A2(n781), .ZN(n804) );
  NAND2_X2 U1489 ( .A1(mem_18__17_), .A2(n781), .ZN(n805) );
  NAND2_X2 U1491 ( .A1(mem_18__16_), .A2(n2977), .ZN(n806) );
  NAND2_X2 U1493 ( .A1(mem_18__15_), .A2(n2977), .ZN(n807) );
  NAND2_X2 U1495 ( .A1(mem_18__14_), .A2(n781), .ZN(n808) );
  NAND2_X2 U1497 ( .A1(mem_18__13_), .A2(n2977), .ZN(n809) );
  NAND2_X2 U1499 ( .A1(mem_18__12_), .A2(n2977), .ZN(n810) );
  NAND2_X2 U1501 ( .A1(mem_18__11_), .A2(n781), .ZN(n811) );
  NAND2_X2 U1503 ( .A1(mem_18__10_), .A2(n2977), .ZN(n812) );
  NAND2_X2 U1505 ( .A1(mem_18__0_), .A2(n781), .ZN(n813) );
  NAND2_X2 U1506 ( .A1(n780), .A2(n174), .ZN(n781) );
  NAND2_X2 U1508 ( .A1(mem_17__9_), .A2(n2972), .ZN(n815) );
  NAND2_X2 U1510 ( .A1(mem_17__8_), .A2(n2971), .ZN(n816) );
  NAND2_X2 U1512 ( .A1(mem_17__7_), .A2(n2971), .ZN(n817) );
  NAND2_X2 U1514 ( .A1(mem_17__6_), .A2(n2971), .ZN(n818) );
  NAND2_X2 U1516 ( .A1(mem_17__5_), .A2(n2972), .ZN(n819) );
  NAND2_X2 U1518 ( .A1(mem_17__4_), .A2(n2971), .ZN(n820) );
  NAND2_X2 U1520 ( .A1(mem_17__3_), .A2(n2970), .ZN(n821) );
  NAND2_X2 U1522 ( .A1(mem_17__31_), .A2(n2970), .ZN(n822) );
  NAND2_X2 U1524 ( .A1(mem_17__30_), .A2(n2972), .ZN(n823) );
  NAND2_X2 U1526 ( .A1(mem_17__2_), .A2(n2972), .ZN(n824) );
  NAND2_X2 U1528 ( .A1(mem_17__29_), .A2(n2970), .ZN(n825) );
  NAND2_X2 U1530 ( .A1(mem_17__28_), .A2(n2972), .ZN(n826) );
  NAND2_X2 U1532 ( .A1(mem_17__27_), .A2(n2970), .ZN(n827) );
  NAND2_X2 U1534 ( .A1(mem_17__26_), .A2(n2972), .ZN(n828) );
  NAND2_X2 U1536 ( .A1(mem_17__25_), .A2(n2970), .ZN(n829) );
  NAND2_X2 U1538 ( .A1(mem_17__24_), .A2(n2971), .ZN(n830) );
  NAND2_X2 U1540 ( .A1(mem_17__23_), .A2(n814), .ZN(n831) );
  NAND2_X2 U1542 ( .A1(mem_17__22_), .A2(n814), .ZN(n832) );
  NAND2_X2 U1544 ( .A1(mem_17__21_), .A2(n2972), .ZN(n833) );
  NAND2_X2 U1546 ( .A1(mem_17__20_), .A2(n814), .ZN(n834) );
  NAND2_X2 U1548 ( .A1(mem_17__1_), .A2(n814), .ZN(n835) );
  NAND2_X2 U1550 ( .A1(mem_17__19_), .A2(n814), .ZN(n836) );
  NAND2_X2 U1552 ( .A1(mem_17__18_), .A2(n814), .ZN(n837) );
  NAND2_X2 U1554 ( .A1(mem_17__17_), .A2(n814), .ZN(n838) );
  NAND2_X2 U1556 ( .A1(mem_17__16_), .A2(n2972), .ZN(n839) );
  NAND2_X2 U1558 ( .A1(mem_17__15_), .A2(n2972), .ZN(n840) );
  NAND2_X2 U1560 ( .A1(mem_17__14_), .A2(n814), .ZN(n841) );
  NAND2_X2 U1562 ( .A1(mem_17__13_), .A2(n2972), .ZN(n842) );
  NAND2_X2 U1564 ( .A1(mem_17__12_), .A2(n2972), .ZN(n843) );
  NAND2_X2 U1566 ( .A1(mem_17__11_), .A2(n814), .ZN(n844) );
  NAND2_X2 U1568 ( .A1(mem_17__10_), .A2(n2972), .ZN(n845) );
  NAND2_X2 U1570 ( .A1(mem_17__0_), .A2(n814), .ZN(n846) );
  NAND2_X2 U1571 ( .A1(n780), .A2(n70), .ZN(n814) );
  NAND2_X2 U1573 ( .A1(mem_16__9_), .A2(n2968), .ZN(n848) );
  NAND2_X2 U1575 ( .A1(mem_16__8_), .A2(n2967), .ZN(n849) );
  NAND2_X2 U1577 ( .A1(mem_16__7_), .A2(n2967), .ZN(n850) );
  NAND2_X2 U1579 ( .A1(mem_16__6_), .A2(n2967), .ZN(n851) );
  NAND2_X2 U1581 ( .A1(mem_16__5_), .A2(n2968), .ZN(n852) );
  NAND2_X2 U1583 ( .A1(mem_16__4_), .A2(n2966), .ZN(n853) );
  NAND2_X2 U1585 ( .A1(mem_16__3_), .A2(n2967), .ZN(n854) );
  NAND2_X2 U1587 ( .A1(mem_16__31_), .A2(n2966), .ZN(n855) );
  NAND2_X2 U1589 ( .A1(mem_16__30_), .A2(n2968), .ZN(n856) );
  NAND2_X2 U1591 ( .A1(mem_16__2_), .A2(n2968), .ZN(n857) );
  NAND2_X2 U1593 ( .A1(mem_16__29_), .A2(n2966), .ZN(n858) );
  NAND2_X2 U1595 ( .A1(mem_16__28_), .A2(n2968), .ZN(n859) );
  NAND2_X2 U1597 ( .A1(mem_16__27_), .A2(n2966), .ZN(n860) );
  NAND2_X2 U1599 ( .A1(mem_16__26_), .A2(n2968), .ZN(n861) );
  NAND2_X2 U1601 ( .A1(mem_16__25_), .A2(n2966), .ZN(n862) );
  NAND2_X2 U1603 ( .A1(mem_16__24_), .A2(n2967), .ZN(n863) );
  NAND2_X2 U1605 ( .A1(mem_16__23_), .A2(n847), .ZN(n864) );
  NAND2_X2 U1607 ( .A1(mem_16__22_), .A2(n847), .ZN(n865) );
  NAND2_X2 U1609 ( .A1(mem_16__21_), .A2(n2968), .ZN(n866) );
  NAND2_X2 U1611 ( .A1(mem_16__20_), .A2(n847), .ZN(n867) );
  NAND2_X2 U1613 ( .A1(mem_16__1_), .A2(n847), .ZN(n868) );
  NAND2_X2 U1615 ( .A1(mem_16__19_), .A2(n847), .ZN(n869) );
  NAND2_X2 U1617 ( .A1(mem_16__18_), .A2(n847), .ZN(n870) );
  NAND2_X2 U1619 ( .A1(mem_16__17_), .A2(n847), .ZN(n871) );
  NAND2_X2 U1621 ( .A1(mem_16__16_), .A2(n2968), .ZN(n872) );
  NAND2_X2 U1623 ( .A1(mem_16__15_), .A2(n2968), .ZN(n873) );
  NAND2_X2 U1625 ( .A1(mem_16__14_), .A2(n847), .ZN(n874) );
  NAND2_X2 U1627 ( .A1(mem_16__13_), .A2(n2968), .ZN(n875) );
  NAND2_X2 U1629 ( .A1(mem_16__12_), .A2(n2968), .ZN(n876) );
  NAND2_X2 U1631 ( .A1(mem_16__11_), .A2(n847), .ZN(n877) );
  NAND2_X2 U1633 ( .A1(mem_16__10_), .A2(n2968), .ZN(n878) );
  NAND2_X2 U1635 ( .A1(mem_16__0_), .A2(n847), .ZN(n879) );
  NAND2_X2 U1636 ( .A1(n780), .A2(n105), .ZN(n847) );
  AND2_X2 U1637 ( .A1(n443), .A2(n746), .ZN(n780) );
  AND2_X2 U1638 ( .A1(rd[4]), .A2(regWr), .ZN(n443) );
  NAND2_X2 U1640 ( .A1(mem_15__9_), .A2(n2965), .ZN(n881) );
  NAND2_X2 U1642 ( .A1(mem_15__8_), .A2(n2964), .ZN(n882) );
  NAND2_X2 U1644 ( .A1(mem_15__7_), .A2(n2963), .ZN(n883) );
  NAND2_X2 U1646 ( .A1(mem_15__6_), .A2(n2964), .ZN(n884) );
  NAND2_X2 U1648 ( .A1(mem_15__5_), .A2(n2963), .ZN(n885) );
  NAND2_X2 U1650 ( .A1(mem_15__4_), .A2(n2964), .ZN(n886) );
  NAND2_X2 U1652 ( .A1(mem_15__3_), .A2(n2963), .ZN(n887) );
  NAND2_X2 U1658 ( .A1(mem_15__2_), .A2(n880), .ZN(n890) );
  NAND2_X2 U1674 ( .A1(mem_15__22_), .A2(n880), .ZN(n898) );
  NAND2_X2 U1676 ( .A1(mem_15__21_), .A2(n880), .ZN(n899) );
  NAND2_X2 U1678 ( .A1(mem_15__20_), .A2(n880), .ZN(n900) );
  NAND2_X2 U1680 ( .A1(mem_15__1_), .A2(n880), .ZN(n901) );
  NAND2_X2 U1682 ( .A1(mem_15__19_), .A2(n880), .ZN(n902) );
  NAND2_X2 U1684 ( .A1(mem_15__18_), .A2(n880), .ZN(n903) );
  NAND2_X2 U1686 ( .A1(mem_15__17_), .A2(n880), .ZN(n904) );
  NAND2_X2 U1688 ( .A1(mem_15__16_), .A2(n2965), .ZN(n905) );
  NAND2_X2 U1690 ( .A1(mem_15__15_), .A2(n2965), .ZN(n906) );
  NAND2_X2 U1692 ( .A1(mem_15__14_), .A2(n880), .ZN(n907) );
  NAND2_X2 U1694 ( .A1(mem_15__13_), .A2(n2965), .ZN(n908) );
  NAND2_X2 U1696 ( .A1(mem_15__12_), .A2(n2965), .ZN(n909) );
  NAND2_X2 U1698 ( .A1(mem_15__11_), .A2(n880), .ZN(n910) );
  NAND2_X2 U1700 ( .A1(mem_15__10_), .A2(n2965), .ZN(n911) );
  NAND2_X2 U1702 ( .A1(mem_15__0_), .A2(n880), .ZN(n912) );
  NAND2_X2 U1703 ( .A1(n913), .A2(n139), .ZN(n880) );
  NAND2_X2 U1705 ( .A1(mem_14__9_), .A2(n2961), .ZN(n915) );
  NAND2_X2 U1707 ( .A1(mem_14__8_), .A2(n2960), .ZN(n916) );
  NAND2_X2 U1709 ( .A1(mem_14__7_), .A2(n2959), .ZN(n917) );
  NAND2_X2 U1711 ( .A1(mem_14__6_), .A2(n2960), .ZN(n918) );
  NAND2_X2 U1713 ( .A1(mem_14__5_), .A2(n2959), .ZN(n919) );
  NAND2_X2 U1715 ( .A1(mem_14__4_), .A2(n2960), .ZN(n920) );
  NAND2_X2 U1717 ( .A1(mem_14__3_), .A2(n2959), .ZN(n921) );
  NAND2_X2 U1723 ( .A1(mem_14__2_), .A2(n914), .ZN(n924) );
  NAND2_X2 U1739 ( .A1(mem_14__22_), .A2(n914), .ZN(n932) );
  NAND2_X2 U1741 ( .A1(mem_14__21_), .A2(n914), .ZN(n933) );
  NAND2_X2 U1743 ( .A1(mem_14__20_), .A2(n914), .ZN(n934) );
  NAND2_X2 U1745 ( .A1(mem_14__1_), .A2(n914), .ZN(n935) );
  NAND2_X2 U1747 ( .A1(mem_14__19_), .A2(n914), .ZN(n936) );
  NAND2_X2 U1749 ( .A1(mem_14__18_), .A2(n914), .ZN(n937) );
  NAND2_X2 U1751 ( .A1(mem_14__17_), .A2(n914), .ZN(n938) );
  NAND2_X2 U1753 ( .A1(mem_14__16_), .A2(n2961), .ZN(n939) );
  NAND2_X2 U1755 ( .A1(mem_14__15_), .A2(n2961), .ZN(n940) );
  NAND2_X2 U1757 ( .A1(mem_14__14_), .A2(n914), .ZN(n941) );
  NAND2_X2 U1759 ( .A1(mem_14__13_), .A2(n2961), .ZN(n942) );
  NAND2_X2 U1761 ( .A1(mem_14__12_), .A2(n2961), .ZN(n943) );
  NAND2_X2 U1763 ( .A1(mem_14__11_), .A2(n914), .ZN(n944) );
  NAND2_X2 U1765 ( .A1(mem_14__10_), .A2(n2961), .ZN(n945) );
  NAND2_X2 U1767 ( .A1(mem_14__0_), .A2(n914), .ZN(n946) );
  NAND2_X2 U1768 ( .A1(n913), .A2(n174), .ZN(n914) );
  NAND2_X2 U1770 ( .A1(mem_13__9_), .A2(n2956), .ZN(n948) );
  NAND2_X2 U1772 ( .A1(mem_13__8_), .A2(n2955), .ZN(n949) );
  NAND2_X2 U1774 ( .A1(mem_13__7_), .A2(n2955), .ZN(n950) );
  NAND2_X2 U1776 ( .A1(mem_13__6_), .A2(n2955), .ZN(n951) );
  NAND2_X2 U1778 ( .A1(mem_13__5_), .A2(n2954), .ZN(n952) );
  NAND2_X2 U1780 ( .A1(mem_13__4_), .A2(n2956), .ZN(n953) );
  NAND2_X2 U1782 ( .A1(mem_13__3_), .A2(n2955), .ZN(n954) );
  NAND2_X2 U1784 ( .A1(mem_13__31_), .A2(n2954), .ZN(n955) );
  NAND2_X2 U1786 ( .A1(mem_13__30_), .A2(n2956), .ZN(n956) );
  NAND2_X2 U1788 ( .A1(mem_13__2_), .A2(n2956), .ZN(n957) );
  NAND2_X2 U1790 ( .A1(mem_13__29_), .A2(n2954), .ZN(n958) );
  NAND2_X2 U1792 ( .A1(mem_13__28_), .A2(n2956), .ZN(n959) );
  NAND2_X2 U1794 ( .A1(mem_13__27_), .A2(n2954), .ZN(n960) );
  NAND2_X2 U1796 ( .A1(mem_13__26_), .A2(n2956), .ZN(n961) );
  NAND2_X2 U1798 ( .A1(mem_13__25_), .A2(n2954), .ZN(n962) );
  NAND2_X2 U1800 ( .A1(mem_13__24_), .A2(n2955), .ZN(n963) );
  NAND2_X2 U1802 ( .A1(mem_13__23_), .A2(n947), .ZN(n964) );
  NAND2_X2 U1804 ( .A1(mem_13__22_), .A2(n947), .ZN(n965) );
  NAND2_X2 U1806 ( .A1(mem_13__21_), .A2(n2956), .ZN(n966) );
  NAND2_X2 U1808 ( .A1(mem_13__20_), .A2(n947), .ZN(n967) );
  NAND2_X2 U1810 ( .A1(mem_13__1_), .A2(n947), .ZN(n968) );
  NAND2_X2 U1812 ( .A1(mem_13__19_), .A2(n947), .ZN(n969) );
  NAND2_X2 U1814 ( .A1(mem_13__18_), .A2(n947), .ZN(n970) );
  NAND2_X2 U1816 ( .A1(mem_13__17_), .A2(n947), .ZN(n971) );
  NAND2_X2 U1818 ( .A1(mem_13__16_), .A2(n2956), .ZN(n972) );
  NAND2_X2 U1820 ( .A1(mem_13__15_), .A2(n2956), .ZN(n973) );
  NAND2_X2 U1822 ( .A1(mem_13__14_), .A2(n947), .ZN(n974) );
  NAND2_X2 U1824 ( .A1(mem_13__13_), .A2(n2956), .ZN(n975) );
  NAND2_X2 U1826 ( .A1(mem_13__12_), .A2(n2956), .ZN(n976) );
  NAND2_X2 U1828 ( .A1(mem_13__11_), .A2(n947), .ZN(n977) );
  NAND2_X2 U1830 ( .A1(mem_13__10_), .A2(n2956), .ZN(n978) );
  NAND2_X2 U1832 ( .A1(mem_13__0_), .A2(n947), .ZN(n979) );
  NAND2_X2 U1833 ( .A1(n913), .A2(n70), .ZN(n947) );
  NAND2_X2 U1836 ( .A1(mem_12__9_), .A2(n2953), .ZN(n982) );
  NAND2_X2 U1838 ( .A1(mem_12__8_), .A2(n2952), .ZN(n983) );
  NAND2_X2 U1840 ( .A1(mem_12__7_), .A2(n2951), .ZN(n984) );
  NAND2_X2 U1842 ( .A1(mem_12__6_), .A2(n2952), .ZN(n985) );
  NAND2_X2 U1844 ( .A1(mem_12__5_), .A2(n2951), .ZN(n986) );
  NAND2_X2 U1846 ( .A1(mem_12__4_), .A2(n2952), .ZN(n987) );
  NAND2_X2 U1848 ( .A1(mem_12__3_), .A2(n2951), .ZN(n988) );
  NAND2_X2 U1854 ( .A1(mem_12__2_), .A2(n981), .ZN(n991) );
  NAND2_X2 U1870 ( .A1(mem_12__22_), .A2(n981), .ZN(n999) );
  NAND2_X2 U1872 ( .A1(mem_12__21_), .A2(n981), .ZN(n1000) );
  NAND2_X2 U1874 ( .A1(mem_12__20_), .A2(n981), .ZN(n1001) );
  NAND2_X2 U1876 ( .A1(mem_12__1_), .A2(n981), .ZN(n1002) );
  NAND2_X2 U1878 ( .A1(mem_12__19_), .A2(n981), .ZN(n1003) );
  NAND2_X2 U1880 ( .A1(mem_12__18_), .A2(n981), .ZN(n1004) );
  NAND2_X2 U1882 ( .A1(mem_12__17_), .A2(n981), .ZN(n1005) );
  NAND2_X2 U1884 ( .A1(mem_12__16_), .A2(n2953), .ZN(n1006) );
  NAND2_X2 U1886 ( .A1(mem_12__15_), .A2(n2953), .ZN(n1007) );
  NAND2_X2 U1888 ( .A1(mem_12__14_), .A2(n981), .ZN(n1008) );
  NAND2_X2 U1890 ( .A1(mem_12__13_), .A2(n2953), .ZN(n1009) );
  NAND2_X2 U1892 ( .A1(mem_12__12_), .A2(n2953), .ZN(n1010) );
  NAND2_X2 U1894 ( .A1(mem_12__11_), .A2(n981), .ZN(n1011) );
  NAND2_X2 U1896 ( .A1(mem_12__10_), .A2(n2953), .ZN(n1012) );
  NAND2_X2 U1898 ( .A1(mem_12__0_), .A2(n981), .ZN(n1013) );
  NAND2_X2 U1899 ( .A1(n913), .A2(n105), .ZN(n981) );
  AND2_X2 U1900 ( .A1(n444), .A2(n242), .ZN(n913) );
  NAND2_X2 U1904 ( .A1(mem_11__9_), .A2(n2949), .ZN(n1016) );
  NAND2_X2 U1906 ( .A1(mem_11__8_), .A2(n2948), .ZN(n1017) );
  NAND2_X2 U1908 ( .A1(mem_11__7_), .A2(n2947), .ZN(n1018) );
  NAND2_X2 U1910 ( .A1(mem_11__6_), .A2(n2948), .ZN(n1019) );
  NAND2_X2 U1912 ( .A1(mem_11__5_), .A2(n2947), .ZN(n1020) );
  NAND2_X2 U1914 ( .A1(mem_11__4_), .A2(n2948), .ZN(n1021) );
  NAND2_X2 U1916 ( .A1(mem_11__3_), .A2(n2947), .ZN(n1022) );
  NAND2_X2 U1922 ( .A1(mem_11__2_), .A2(n1015), .ZN(n1025) );
  NAND2_X2 U1938 ( .A1(mem_11__22_), .A2(n1015), .ZN(n1033) );
  NAND2_X2 U1940 ( .A1(mem_11__21_), .A2(n1015), .ZN(n1034) );
  NAND2_X2 U1942 ( .A1(mem_11__20_), .A2(n1015), .ZN(n1035) );
  NAND2_X2 U1944 ( .A1(mem_11__1_), .A2(n1015), .ZN(n1036) );
  NAND2_X2 U1946 ( .A1(mem_11__19_), .A2(n1015), .ZN(n1037) );
  NAND2_X2 U1948 ( .A1(mem_11__18_), .A2(n1015), .ZN(n1038) );
  NAND2_X2 U1950 ( .A1(mem_11__17_), .A2(n1015), .ZN(n1039) );
  NAND2_X2 U1952 ( .A1(mem_11__16_), .A2(n2949), .ZN(n1040) );
  NAND2_X2 U1954 ( .A1(mem_11__15_), .A2(n2949), .ZN(n1041) );
  NAND2_X2 U1956 ( .A1(mem_11__14_), .A2(n1015), .ZN(n1042) );
  NAND2_X2 U1958 ( .A1(mem_11__13_), .A2(n2949), .ZN(n1043) );
  NAND2_X2 U1960 ( .A1(mem_11__12_), .A2(n2949), .ZN(n1044) );
  NAND2_X2 U1962 ( .A1(mem_11__11_), .A2(n1015), .ZN(n1045) );
  NAND2_X2 U1964 ( .A1(mem_11__10_), .A2(n2949), .ZN(n1046) );
  NAND2_X2 U1966 ( .A1(mem_11__0_), .A2(n1015), .ZN(n1047) );
  NAND2_X2 U1967 ( .A1(n139), .A2(n71), .ZN(n1015) );
  AND2_X2 U1968 ( .A1(rd[1]), .A2(rd[0]), .ZN(n139) );
  NAND2_X2 U1970 ( .A1(mem_10__9_), .A2(n2945), .ZN(n1049) );
  NAND2_X2 U1972 ( .A1(mem_10__8_), .A2(n2944), .ZN(n1050) );
  NAND2_X2 U1974 ( .A1(mem_10__7_), .A2(n2943), .ZN(n1051) );
  NAND2_X2 U1976 ( .A1(mem_10__6_), .A2(n2944), .ZN(n1052) );
  NAND2_X2 U1978 ( .A1(mem_10__5_), .A2(n2943), .ZN(n1053) );
  NAND2_X2 U1980 ( .A1(mem_10__4_), .A2(n2944), .ZN(n1054) );
  NAND2_X2 U1982 ( .A1(mem_10__3_), .A2(n2943), .ZN(n1055) );
  NAND2_X2 U1988 ( .A1(mem_10__2_), .A2(n1048), .ZN(n1058) );
  NAND2_X2 U2004 ( .A1(mem_10__22_), .A2(n1048), .ZN(n1066) );
  NAND2_X2 U2006 ( .A1(mem_10__21_), .A2(n1048), .ZN(n1067) );
  NAND2_X2 U2008 ( .A1(mem_10__20_), .A2(n1048), .ZN(n1068) );
  NAND2_X2 U2010 ( .A1(mem_10__1_), .A2(n1048), .ZN(n1069) );
  NAND2_X2 U2012 ( .A1(mem_10__19_), .A2(n1048), .ZN(n1070) );
  NAND2_X2 U2014 ( .A1(mem_10__18_), .A2(n1048), .ZN(n1071) );
  NAND2_X2 U2016 ( .A1(mem_10__17_), .A2(n1048), .ZN(n1072) );
  NAND2_X2 U2018 ( .A1(mem_10__16_), .A2(n2945), .ZN(n1073) );
  NAND2_X2 U2020 ( .A1(mem_10__15_), .A2(n2945), .ZN(n1074) );
  NAND2_X2 U2022 ( .A1(mem_10__14_), .A2(n1048), .ZN(n1075) );
  NAND2_X2 U2024 ( .A1(mem_10__13_), .A2(n2945), .ZN(n1076) );
  NAND2_X2 U2026 ( .A1(mem_10__12_), .A2(n2945), .ZN(n1077) );
  NAND2_X2 U2028 ( .A1(mem_10__11_), .A2(n1048), .ZN(n1078) );
  NAND2_X2 U2030 ( .A1(mem_10__10_), .A2(n2945), .ZN(n1079) );
  NAND2_X2 U2032 ( .A1(mem_10__0_), .A2(n1048), .ZN(n1080) );
  NAND2_X2 U2033 ( .A1(n174), .A2(n71), .ZN(n1048) );
  AND2_X2 U2034 ( .A1(n242), .A2(n578), .ZN(n71) );
  AND2_X2 U2037 ( .A1(regWr), .A2(n7227), .ZN(n242) );
  AND2_X2 U2038 ( .A1(rd[1]), .A2(n7230), .ZN(n174) );
  AND2_X2 U2040 ( .A1(mem_0__9_), .A2(n2940), .ZN(n1159) );
  AND2_X2 U2041 ( .A1(mem_0__8_), .A2(n2941), .ZN(n1158) );
  AND2_X2 U2042 ( .A1(mem_0__7_), .A2(n2940), .ZN(n1157) );
  AND2_X2 U2043 ( .A1(mem_0__6_), .A2(n2941), .ZN(n1156) );
  AND2_X2 U2044 ( .A1(mem_0__5_), .A2(n2940), .ZN(n1155) );
  AND2_X2 U2045 ( .A1(mem_0__4_), .A2(n2941), .ZN(n1154) );
  AND2_X2 U2046 ( .A1(mem_0__3_), .A2(n2940), .ZN(n1153) );
  AND2_X2 U2047 ( .A1(mem_0__31_), .A2(n2941), .ZN(n1181) );
  AND2_X2 U2048 ( .A1(mem_0__30_), .A2(n2940), .ZN(n1180) );
  AND2_X2 U2049 ( .A1(mem_0__2_), .A2(n2941), .ZN(n1152) );
  AND2_X2 U2050 ( .A1(mem_0__29_), .A2(n2941), .ZN(n1179) );
  AND2_X2 U2051 ( .A1(mem_0__28_), .A2(n2941), .ZN(n1178) );
  AND2_X2 U2052 ( .A1(mem_0__27_), .A2(n2941), .ZN(n1177) );
  AND2_X2 U2053 ( .A1(mem_0__26_), .A2(n2941), .ZN(n1176) );
  AND2_X2 U2054 ( .A1(mem_0__25_), .A2(n2941), .ZN(n1175) );
  AND2_X2 U2055 ( .A1(mem_0__24_), .A2(n2941), .ZN(n1174) );
  AND2_X2 U2056 ( .A1(mem_0__23_), .A2(n2941), .ZN(n1173) );
  AND2_X2 U2057 ( .A1(mem_0__22_), .A2(n2941), .ZN(n1172) );
  AND2_X2 U2058 ( .A1(mem_0__21_), .A2(n2941), .ZN(n1171) );
  AND2_X2 U2059 ( .A1(mem_0__20_), .A2(n2941), .ZN(n1170) );
  AND2_X2 U2060 ( .A1(mem_0__1_), .A2(n2941), .ZN(n1151) );
  AND2_X2 U2061 ( .A1(mem_0__19_), .A2(n2940), .ZN(n1169) );
  AND2_X2 U2062 ( .A1(mem_0__18_), .A2(n2940), .ZN(n1168) );
  AND2_X2 U2063 ( .A1(mem_0__17_), .A2(n2940), .ZN(n1167) );
  AND2_X2 U2064 ( .A1(mem_0__16_), .A2(n2940), .ZN(n1166) );
  AND2_X2 U2065 ( .A1(mem_0__15_), .A2(n2940), .ZN(n1165) );
  AND2_X2 U2066 ( .A1(mem_0__14_), .A2(n2940), .ZN(n1164) );
  AND2_X2 U2067 ( .A1(mem_0__13_), .A2(n2940), .ZN(n1163) );
  AND2_X2 U2068 ( .A1(mem_0__12_), .A2(n2940), .ZN(n1162) );
  AND2_X2 U2069 ( .A1(mem_0__11_), .A2(n2940), .ZN(n1161) );
  AND2_X2 U2070 ( .A1(mem_0__10_), .A2(n2940), .ZN(n1160) );
  AND2_X2 U2071 ( .A1(mem_0__0_), .A2(n2940), .ZN(n1150) );
  DFF_X1 rData2_reg_24_ ( .D(N217), .CK(n2238), .Q(rData2[24]) );
  DFF_X1 rData2_reg_27_ ( .D(N220), .CK(n2238), .Q(rData2[27]) );
  NOR2_X4 U2239 ( .A1(mem_23__23_), .A2(n2804), .ZN(n4140) );
  NOR2_X4 U2240 ( .A1(mem_23__24_), .A2(n2804), .ZN(n4203) );
  NAND2_X4 U2241 ( .A1(n4616), .A2(n4615), .ZN(n4625) );
  NAND2_X4 U2242 ( .A1(n4553), .A2(n4552), .ZN(n4562) );
  NOR2_X1 U2243 ( .A1(mem_6__31_), .A2(n2798), .ZN(n4612) );
  NOR2_X1 U2244 ( .A1(mem_6__30_), .A2(n2798), .ZN(n4549) );
  OAI21_X1 U2245 ( .B1(mem_7__2_), .B2(n2810), .A(n2757), .ZN(n3265) );
  NOR2_X2 U2246 ( .A1(n4468), .A2(n4467), .ZN(n4471) );
  MUX2_X1 U2247 ( .A(n4482), .B(n4481), .S(n3113), .Z(n4483) );
  INV_X16 U2248 ( .A(n2830), .ZN(n2839) );
  NAND2_X4 U2249 ( .A1(n4413), .A2(n4412), .ZN(n4416) );
  NAND3_X1 U2250 ( .A1(n2770), .A2(mem_1__26_), .A3(n3144), .ZN(n4307) );
  NAND3_X1 U2251 ( .A1(n2770), .A2(mem_1__23_), .A3(n3142), .ZN(n4118) );
  NAND3_X1 U2252 ( .A1(n2770), .A2(mem_17__23_), .A3(n3142), .ZN(n4148) );
  NAND3_X1 U2253 ( .A1(n2770), .A2(mem_1__25_), .A3(n3143), .ZN(n4244) );
  NAND3_X1 U2254 ( .A1(n2770), .A2(mem_17__24_), .A3(n3143), .ZN(n4211) );
  NAND3_X2 U2255 ( .A1(n2770), .A2(mem_17__28_), .A3(n3146), .ZN(n4463) );
  NAND3_X2 U2256 ( .A1(n2770), .A2(mem_17__25_), .A3(n3144), .ZN(n4274) );
  NAND3_X2 U2257 ( .A1(n2770), .A2(mem_17__29_), .A3(n3146), .ZN(n4526) );
  NAND3_X4 U2258 ( .A1(n2770), .A2(mem_25__25_), .A3(n3144), .ZN(n4288) );
  NOR2_X1 U2259 ( .A1(mem_4__2_), .A2(n2322), .ZN(n3261) );
  NOR2_X1 U2260 ( .A1(mem_4__3_), .A2(n2322), .ZN(n3301) );
  NOR2_X1 U2261 ( .A1(mem_4__19_), .A2(n2322), .ZN(n3942) );
  NOR2_X1 U2262 ( .A1(mem_4__4_), .A2(n2322), .ZN(n3341) );
  NOR2_X1 U2263 ( .A1(mem_20__15_), .A2(n2322), .ZN(n3800) );
  NOR2_X1 U2264 ( .A1(mem_20__18_), .A2(n2322), .ZN(n3920) );
  NOR2_X1 U2265 ( .A1(mem_12__15_), .A2(n2322), .ZN(n3790) );
  NOR2_X1 U2266 ( .A1(mem_20__11_), .A2(n2322), .ZN(n3639) );
  NOR2_X1 U2267 ( .A1(mem_20__10_), .A2(n2322), .ZN(n3599) );
  NOR2_X1 U2268 ( .A1(mem_20__19_), .A2(n2322), .ZN(n3960) );
  NOR2_X1 U2269 ( .A1(mem_12__20_), .A2(n2322), .ZN(n3990) );
  NOR2_X1 U2270 ( .A1(mem_12__5_), .A2(n2322), .ZN(n3389) );
  NOR2_X1 U2271 ( .A1(mem_28__16_), .A2(n2322), .ZN(n3848) );
  NOR2_X1 U2272 ( .A1(mem_28__3_), .A2(n2322), .ZN(n3327) );
  NOR2_X1 U2273 ( .A1(mem_28__10_), .A2(n2322), .ZN(n3607) );
  NOR2_X1 U2274 ( .A1(mem_28__18_), .A2(n2322), .ZN(n3928) );
  NOR2_X1 U2275 ( .A1(mem_28__2_), .A2(n2322), .ZN(n3287) );
  NOR2_X4 U2276 ( .A1(mem_12__25_), .A2(n2322), .ZN(n4254) );
  NOR2_X4 U2277 ( .A1(mem_28__26_), .A2(n2322), .ZN(n4347) );
  NOR2_X4 U2278 ( .A1(n2693), .A2(n2322), .ZN(n4410) );
  NAND2_X4 U2279 ( .A1(n5798), .A2(n3110), .ZN(n6146) );
  INV_X8 U2280 ( .A(rs1[0]), .ZN(n3110) );
  MUX2_X1 U2281 ( .A(n5951), .B(n5950), .S(n3063), .Z(n5952) );
  INV_X16 U2282 ( .A(n2865), .ZN(n2872) );
  INV_X8 U2283 ( .A(n2431), .ZN(n2865) );
  INV_X4 U2284 ( .A(n2829), .ZN(n2239) );
  INV_X4 U2285 ( .A(n2239), .ZN(n2240) );
  INV_X4 U2286 ( .A(n2239), .ZN(n2241) );
  INV_X4 U2287 ( .A(n2239), .ZN(n2242) );
  INV_X4 U2288 ( .A(n2239), .ZN(n2243) );
  INV_X4 U2289 ( .A(n2239), .ZN(n2244) );
  INV_X2 U2290 ( .A(n2827), .ZN(n2245) );
  INV_X2 U2291 ( .A(n2245), .ZN(n2246) );
  INV_X2 U2292 ( .A(n2245), .ZN(n2247) );
  INV_X2 U2293 ( .A(n2245), .ZN(n2248) );
  INV_X2 U2294 ( .A(n2245), .ZN(n2249) );
  INV_X2 U2295 ( .A(n2245), .ZN(n2250) );
  INV_X16 U2296 ( .A(n2826), .ZN(n2251) );
  INV_X4 U2297 ( .A(n2251), .ZN(n2252) );
  INV_X4 U2298 ( .A(n2251), .ZN(n2253) );
  INV_X2 U2299 ( .A(n2251), .ZN(n2254) );
  INV_X2 U2300 ( .A(n2251), .ZN(n2255) );
  INV_X2 U2301 ( .A(n2251), .ZN(n2256) );
  INV_X16 U2302 ( .A(n2821), .ZN(n2257) );
  INV_X4 U2303 ( .A(n2257), .ZN(n2258) );
  INV_X4 U2304 ( .A(n2257), .ZN(n2259) );
  INV_X2 U2305 ( .A(n2257), .ZN(n2260) );
  INV_X2 U2306 ( .A(n2257), .ZN(n2261) );
  INV_X2 U2307 ( .A(n2257), .ZN(n2262) );
  INV_X8 U2308 ( .A(n2820), .ZN(n2263) );
  INV_X4 U2309 ( .A(n2263), .ZN(n2264) );
  INV_X4 U2310 ( .A(n2263), .ZN(n2265) );
  INV_X4 U2311 ( .A(n2263), .ZN(n2266) );
  INV_X4 U2312 ( .A(n2263), .ZN(n2267) );
  INV_X4 U2313 ( .A(n2263), .ZN(n2268) );
  INV_X8 U2314 ( .A(n2814), .ZN(n2269) );
  INV_X4 U2315 ( .A(n2269), .ZN(n2270) );
  INV_X4 U2316 ( .A(n2269), .ZN(n2271) );
  INV_X2 U2317 ( .A(n2269), .ZN(n2272) );
  INV_X2 U2318 ( .A(n2269), .ZN(n2273) );
  INV_X2 U2319 ( .A(n2269), .ZN(n2274) );
  INV_X16 U2320 ( .A(n2815), .ZN(n2275) );
  INV_X4 U2321 ( .A(n2275), .ZN(n2276) );
  INV_X4 U2322 ( .A(n2275), .ZN(n2277) );
  INV_X4 U2323 ( .A(n2275), .ZN(n2278) );
  INV_X4 U2324 ( .A(n2275), .ZN(n2279) );
  INV_X4 U2325 ( .A(n2275), .ZN(n2280) );
  INV_X8 U2326 ( .A(n2817), .ZN(n2281) );
  INV_X2 U2327 ( .A(n2281), .ZN(n2282) );
  INV_X4 U2328 ( .A(n2281), .ZN(n2283) );
  INV_X4 U2329 ( .A(n2281), .ZN(n2284) );
  INV_X2 U2330 ( .A(n2281), .ZN(n2285) );
  INV_X2 U2331 ( .A(n2281), .ZN(n2286) );
  INV_X16 U2332 ( .A(n2816), .ZN(n2287) );
  INV_X4 U2333 ( .A(n2287), .ZN(n2288) );
  INV_X4 U2334 ( .A(n2287), .ZN(n2289) );
  INV_X4 U2335 ( .A(n2287), .ZN(n2290) );
  INV_X4 U2336 ( .A(n2287), .ZN(n2291) );
  INV_X4 U2337 ( .A(n2287), .ZN(n2292) );
  INV_X8 U2338 ( .A(n2818), .ZN(n2293) );
  INV_X4 U2339 ( .A(n2293), .ZN(n2294) );
  INV_X4 U2340 ( .A(n2293), .ZN(n2295) );
  INV_X2 U2341 ( .A(n2293), .ZN(n2296) );
  INV_X2 U2342 ( .A(n2293), .ZN(n2297) );
  INV_X4 U2343 ( .A(n2293), .ZN(n2298) );
  INV_X8 U2344 ( .A(n2813), .ZN(n2299) );
  INV_X4 U2345 ( .A(n2299), .ZN(n2300) );
  INV_X4 U2346 ( .A(n2299), .ZN(n2301) );
  INV_X4 U2347 ( .A(n2299), .ZN(n2302) );
  INV_X2 U2348 ( .A(n2299), .ZN(n2303) );
  INV_X2 U2349 ( .A(n2299), .ZN(n2304) );
  INV_X16 U2350 ( .A(n2822), .ZN(n2305) );
  INV_X2 U2351 ( .A(n2305), .ZN(n2306) );
  INV_X2 U2352 ( .A(n2305), .ZN(n2307) );
  INV_X2 U2353 ( .A(n2305), .ZN(n2308) );
  INV_X2 U2354 ( .A(n2305), .ZN(n2309) );
  INV_X2 U2355 ( .A(n2305), .ZN(n2310) );
  INV_X8 U2356 ( .A(n2819), .ZN(n2311) );
  INV_X2 U2357 ( .A(n2311), .ZN(n2312) );
  INV_X2 U2358 ( .A(n2311), .ZN(n2313) );
  INV_X2 U2359 ( .A(n2311), .ZN(n2314) );
  INV_X2 U2360 ( .A(n2311), .ZN(n2315) );
  INV_X2 U2361 ( .A(n2311), .ZN(n2316) );
  INV_X8 U2362 ( .A(n4664), .ZN(n2317) );
  INV_X16 U2363 ( .A(n2317), .ZN(n2318) );
  INV_X16 U2364 ( .A(n2317), .ZN(n2319) );
  INV_X16 U2365 ( .A(n2317), .ZN(n2320) );
  INV_X16 U2366 ( .A(n2317), .ZN(n2321) );
  INV_X8 U2367 ( .A(n2317), .ZN(n2322) );
  NAND2_X4 U2368 ( .A1(n3155), .A2(n3163), .ZN(n4664) );
  INV_X8 U2369 ( .A(n2829), .ZN(n2828) );
  INV_X8 U2370 ( .A(n2827), .ZN(n2823) );
  INV_X4 U2371 ( .A(n2826), .ZN(n2825) );
  INV_X4 U2372 ( .A(n2826), .ZN(n2824) );
  INV_X4 U2373 ( .A(n2828), .ZN(n2827) );
  INV_X4 U2374 ( .A(n2828), .ZN(n2826) );
  INV_X4 U2375 ( .A(n2828), .ZN(n2821) );
  INV_X4 U2376 ( .A(n2828), .ZN(n2820) );
  INV_X2 U2377 ( .A(n2823), .ZN(n2814) );
  INV_X2 U2378 ( .A(n2823), .ZN(n2817) );
  INV_X2 U2379 ( .A(n2823), .ZN(n2813) );
  INV_X4 U2380 ( .A(n2824), .ZN(n2822) );
  INV_X4 U2381 ( .A(n2760), .ZN(n2755) );
  INV_X16 U2382 ( .A(n2787), .ZN(n2783) );
  NAND2_X4 U2383 ( .A1(n4189), .A2(n4188), .ZN(n4198) );
  OAI211_X4 U2384 ( .C1(n4151), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4167)
         );
  OAI211_X4 U2385 ( .C1(n4214), .C2(n4213), .A(n4212), .B(n4211), .ZN(n4230)
         );
  NAND2_X4 U2386 ( .A1(n4147), .A2(n4146), .ZN(n4150) );
  NAND2_X4 U2387 ( .A1(n4210), .A2(n4209), .ZN(n4213) );
  NAND2_X4 U2388 ( .A1(n4399), .A2(n4398), .ZN(n4402) );
  NAND2_X4 U2389 ( .A1(n4194), .A2(n4193), .ZN(n4197) );
  NAND2_X4 U2390 ( .A1(n4635), .A2(n4634), .ZN(n4638) );
  NAND2_X4 U2391 ( .A1(n4630), .A2(n4629), .ZN(n4639) );
  NAND2_X4 U2392 ( .A1(n4572), .A2(n4571), .ZN(n4575) );
  NAND2_X4 U2393 ( .A1(n4567), .A2(n4566), .ZN(n4576) );
  NOR2_X4 U2394 ( .A1(mem_10__23_), .A2(n3132), .ZN(n4129) );
  NAND2_X4 U2395 ( .A1(n4255), .A2(n3162), .ZN(n4256) );
  NAND2_X4 U2396 ( .A1(n4131), .A2(n4130), .ZN(n4134) );
  NOR2_X2 U2397 ( .A1(mem_21__28_), .A2(n2781), .ZN(n4454) );
  OAI211_X4 U2398 ( .C1(n4466), .C2(n4465), .A(n4464), .B(n4463), .ZN(n4482)
         );
  INV_X4 U2399 ( .A(n3161), .ZN(n3158) );
  INV_X8 U2400 ( .A(n3144), .ZN(n3132) );
  INV_X8 U2401 ( .A(n3144), .ZN(n3133) );
  INV_X16 U2402 ( .A(n2801), .ZN(n2812) );
  INV_X8 U2403 ( .A(n2789), .ZN(n2799) );
  INV_X4 U2404 ( .A(rs2[2]), .ZN(n3136) );
  NAND3_X2 U2405 ( .A1(mem_9__1_), .A2(n3156), .A3(n3154), .ZN(n3235) );
  INV_X2 U2406 ( .A(n2765), .ZN(n2763) );
  INV_X8 U2407 ( .A(n2784), .ZN(n2775) );
  INV_X4 U2408 ( .A(n3153), .ZN(n3126) );
  INV_X4 U2409 ( .A(n2760), .ZN(n2754) );
  INV_X4 U2410 ( .A(n2790), .ZN(n2791) );
  INV_X8 U2411 ( .A(n2812), .ZN(n2808) );
  INV_X8 U2412 ( .A(n2784), .ZN(n2776) );
  INV_X4 U2413 ( .A(n3150), .ZN(n3127) );
  INV_X8 U2414 ( .A(n2800), .ZN(n2792) );
  INV_X4 U2415 ( .A(n3151), .ZN(n3128) );
  INV_X4 U2416 ( .A(n2765), .ZN(n2757) );
  INV_X8 U2417 ( .A(n2800), .ZN(n2793) );
  INV_X4 U2418 ( .A(n3138), .ZN(n3129) );
  INV_X8 U2419 ( .A(n2800), .ZN(n2794) );
  INV_X4 U2420 ( .A(n2760), .ZN(n2758) );
  INV_X8 U2421 ( .A(n2783), .ZN(n2778) );
  INV_X8 U2422 ( .A(n2783), .ZN(n2779) );
  INV_X4 U2423 ( .A(n2760), .ZN(n2759) );
  INV_X8 U2424 ( .A(n2800), .ZN(n2795) );
  INV_X8 U2425 ( .A(n2812), .ZN(n2805) );
  INV_X4 U2426 ( .A(n3152), .ZN(n3131) );
  INV_X4 U2427 ( .A(n2783), .ZN(n2780) );
  INV_X16 U2428 ( .A(n2812), .ZN(n2803) );
  INV_X4 U2429 ( .A(n2812), .ZN(n2810) );
  INV_X8 U2430 ( .A(n2799), .ZN(n2797) );
  INV_X8 U2431 ( .A(n2783), .ZN(n2781) );
  INV_X4 U2432 ( .A(n2799), .ZN(n2798) );
  INV_X4 U2433 ( .A(n3136), .ZN(n3122) );
  INV_X2 U2434 ( .A(n2783), .ZN(n2782) );
  INV_X4 U2435 ( .A(rs1[0]), .ZN(n3109) );
  INV_X4 U2436 ( .A(n2855), .ZN(n2853) );
  INV_X4 U2437 ( .A(n3106), .ZN(n3087) );
  INV_X4 U2438 ( .A(n2375), .ZN(n2856) );
  INV_X4 U2439 ( .A(n3108), .ZN(n3088) );
  INV_X4 U2440 ( .A(n2855), .ZN(n2852) );
  INV_X4 U2441 ( .A(n2378), .ZN(n2858) );
  INV_X4 U2442 ( .A(n2375), .ZN(n2857) );
  INV_X4 U2443 ( .A(n3105), .ZN(n3086) );
  INV_X4 U2444 ( .A(n2855), .ZN(n2854) );
  INV_X4 U2445 ( .A(n2378), .ZN(n2860) );
  INV_X8 U2446 ( .A(n2875), .ZN(n2874) );
  NOR2_X2 U2447 ( .A1(n4317), .A2(n4316), .ZN(n4320) );
  NOR2_X2 U2448 ( .A1(mem_12__26_), .A2(n2321), .ZN(n4317) );
  NOR2_X2 U2449 ( .A1(n4396), .A2(n4395), .ZN(n4399) );
  NOR2_X2 U2450 ( .A1(mem_19__27_), .A2(n2837), .ZN(n4395) );
  NOR2_X2 U2451 ( .A1(n4191), .A2(n4190), .ZN(n4194) );
  NOR2_X2 U2452 ( .A1(mem_12__24_), .A2(n2318), .ZN(n4191) );
  INV_X16 U2453 ( .A(rs2[0]), .ZN(n3163) );
  NOR3_X2 U2454 ( .A1(n3221), .A2(n3220), .A3(n3219), .ZN(n3227) );
  NOR3_X2 U2455 ( .A1(n3158), .A2(mem_26__1_), .A3(n3125), .ZN(n3220) );
  NOR2_X2 U2456 ( .A1(mem_29__1_), .A2(n2774), .ZN(n3219) );
  INV_X4 U2457 ( .A(n2774), .ZN(n2770) );
  INV_X4 U2458 ( .A(n2773), .ZN(n2771) );
  INV_X4 U2459 ( .A(n3109), .ZN(n3100) );
  INV_X4 U2460 ( .A(n2378), .ZN(n2859) );
  INV_X16 U2461 ( .A(n3068), .ZN(n3067) );
  INV_X16 U2462 ( .A(n2869), .ZN(n2866) );
  INV_X4 U2463 ( .A(n2853), .ZN(n2848) );
  NOR2_X2 U2464 ( .A1(mem_20__23_), .A2(n2321), .ZN(n4144) );
  NOR2_X2 U2465 ( .A1(mem_11__23_), .A2(n2835), .ZN(n4127) );
  NOR2_X2 U2466 ( .A1(mem_13__27_), .A2(n2780), .ZN(n4375) );
  NOR2_X2 U2467 ( .A1(mem_20__24_), .A2(n2321), .ZN(n4207) );
  INV_X8 U2468 ( .A(n2784), .ZN(n2777) );
  INV_X4 U2469 ( .A(n2760), .ZN(n2756) );
  INV_X4 U2470 ( .A(n2788), .ZN(n2786) );
  INV_X4 U2471 ( .A(n3139), .ZN(n3130) );
  INV_X8 U2472 ( .A(n2840), .ZN(n2835) );
  NOR2_X2 U2473 ( .A1(mem_22__28_), .A2(n2797), .ZN(n4453) );
  NOR2_X2 U2474 ( .A1(mem_22__29_), .A2(n2797), .ZN(n4516) );
  NOR2_X2 U2475 ( .A1(mem_13__30_), .A2(n2781), .ZN(n4564) );
  NOR2_X2 U2476 ( .A1(mem_7__30_), .A2(n2808), .ZN(n4551) );
  NOR2_X2 U2477 ( .A1(mem_22__30_), .A2(n2798), .ZN(n4579) );
  NOR2_X2 U2478 ( .A1(mem_7__31_), .A2(n2806), .ZN(n4614) );
  NOR2_X2 U2479 ( .A1(mem_22__31_), .A2(n2798), .ZN(n4642) );
  NOR2_X2 U2480 ( .A1(n2685), .A2(n3132), .ZN(n4159) );
  NOR2_X2 U2481 ( .A1(n4153), .A2(n4152), .ZN(n4156) );
  NOR2_X2 U2482 ( .A1(n2653), .A2(n2804), .ZN(n4154) );
  NOR2_X2 U2483 ( .A1(n4114), .A2(n4113), .ZN(n4117) );
  NOR2_X2 U2484 ( .A1(mem_4__23_), .A2(n2322), .ZN(n4114) );
  NOR2_X2 U2485 ( .A1(mem_3__23_), .A2(n2835), .ZN(n4113) );
  NOR2_X2 U2486 ( .A1(mem_2__23_), .A2(n3131), .ZN(n4115) );
  NOR2_X2 U2487 ( .A1(n4109), .A2(n4108), .ZN(n4112) );
  NOR2_X2 U2488 ( .A1(n2762), .A2(n4110), .ZN(n4111) );
  NOR2_X1 U2489 ( .A1(mem_5__23_), .A2(n2779), .ZN(n4109) );
  NOR2_X2 U2490 ( .A1(mem_2__26_), .A2(n3132), .ZN(n4304) );
  NOR2_X2 U2491 ( .A1(n4303), .A2(n4302), .ZN(n4306) );
  NOR2_X2 U2492 ( .A1(mem_4__26_), .A2(n2319), .ZN(n4303) );
  NOR2_X2 U2493 ( .A1(mem_3__26_), .A2(n2836), .ZN(n4302) );
  NOR2_X2 U2494 ( .A1(n4298), .A2(n4297), .ZN(n4301) );
  NOR2_X1 U2495 ( .A1(mem_5__26_), .A2(n2780), .ZN(n4298) );
  NOR2_X2 U2496 ( .A1(n4347), .A2(n4346), .ZN(n4350) );
  NOR2_X2 U2497 ( .A1(n2633), .A2(n2836), .ZN(n4346) );
  NOR2_X2 U2498 ( .A1(n2645), .A2(n3133), .ZN(n4348) );
  NOR2_X2 U2499 ( .A1(n4342), .A2(n4341), .ZN(n4345) );
  NOR2_X2 U2500 ( .A1(n2631), .A2(n2803), .ZN(n4343) );
  NOR2_X2 U2501 ( .A1(n2737), .A2(n3133), .ZN(n4334) );
  NOR2_X2 U2502 ( .A1(n4333), .A2(n4332), .ZN(n4336) );
  NOR2_X2 U2503 ( .A1(n2675), .A2(n2318), .ZN(n4333) );
  NOR2_X2 U2504 ( .A1(n2655), .A2(n2836), .ZN(n4332) );
  NOR2_X2 U2505 ( .A1(n4328), .A2(n4327), .ZN(n4331) );
  NOR2_X2 U2506 ( .A1(n2639), .A2(n2803), .ZN(n4329) );
  NOR2_X2 U2507 ( .A1(n4410), .A2(n4409), .ZN(n4413) );
  NOR2_X2 U2508 ( .A1(n2723), .A2(n2837), .ZN(n4409) );
  NOR2_X2 U2509 ( .A1(n2733), .A2(n3133), .ZN(n4411) );
  NOR2_X2 U2510 ( .A1(n4405), .A2(n4404), .ZN(n4408) );
  NOR2_X2 U2511 ( .A1(n2665), .A2(n2797), .ZN(n4404) );
  NOR2_X2 U2512 ( .A1(mem_2__27_), .A2(n3133), .ZN(n4367) );
  NOR2_X2 U2513 ( .A1(n4366), .A2(n4365), .ZN(n4369) );
  NOR2_X2 U2514 ( .A1(mem_4__27_), .A2(n2322), .ZN(n4366) );
  NOR2_X2 U2515 ( .A1(mem_3__27_), .A2(n2837), .ZN(n4365) );
  NOR2_X2 U2516 ( .A1(n4361), .A2(n4360), .ZN(n4364) );
  NOR2_X1 U2517 ( .A1(mem_5__27_), .A2(n2780), .ZN(n4361) );
  NOR2_X2 U2518 ( .A1(n4172), .A2(n4171), .ZN(n4175) );
  NOR2_X1 U2519 ( .A1(mem_5__24_), .A2(n2779), .ZN(n4172) );
  NOR2_X1 U2520 ( .A1(mem_6__24_), .A2(n2796), .ZN(n4171) );
  NOR2_X2 U2521 ( .A1(n4177), .A2(n4176), .ZN(n4180) );
  NOR2_X2 U2522 ( .A1(mem_4__24_), .A2(n2319), .ZN(n4177) );
  NOR2_X2 U2523 ( .A1(n4221), .A2(n4220), .ZN(n4224) );
  NOR2_X2 U2524 ( .A1(n2695), .A2(n2320), .ZN(n4221) );
  NOR2_X2 U2525 ( .A1(n2725), .A2(n2836), .ZN(n4220) );
  NOR2_X2 U2526 ( .A1(n2663), .A2(n3132), .ZN(n4222) );
  NOR2_X2 U2527 ( .A1(n4216), .A2(n4215), .ZN(n4219) );
  NOR2_X2 U2528 ( .A1(n2667), .A2(n2796), .ZN(n4215) );
  NOR2_X2 U2529 ( .A1(rd[0]), .A2(rd[1]), .ZN(n105) );
  NOR2_X2 U2530 ( .A1(n7230), .A2(rd[1]), .ZN(n70) );
  NOR2_X2 U2531 ( .A1(mem_12__0_), .A2(n2319), .ZN(n3174) );
  NOR2_X1 U2532 ( .A1(mem_11__0_), .A2(n2838), .ZN(n3173) );
  NOR3_X2 U2533 ( .A1(n3159), .A2(mem_10__0_), .A3(n3125), .ZN(n3175) );
  NOR3_X2 U2534 ( .A1(n3178), .A2(n3177), .A3(n3176), .ZN(n3179) );
  NOR2_X2 U2535 ( .A1(mem_13__0_), .A2(n2774), .ZN(n3177) );
  NOR2_X2 U2536 ( .A1(mem_14__0_), .A2(n2794), .ZN(n3176) );
  OAI21_X1 U2537 ( .B1(mem_15__0_), .B2(n2810), .A(n2754), .ZN(n3178) );
  OAI21_X1 U2538 ( .B1(mem_7__0_), .B2(n2810), .A(n2754), .ZN(n3170) );
  NOR2_X2 U2539 ( .A1(mem_6__0_), .A2(n2794), .ZN(n3168) );
  NOR2_X2 U2540 ( .A1(mem_5__0_), .A2(n2774), .ZN(n3169) );
  NOR2_X2 U2541 ( .A1(mem_4__0_), .A2(n2318), .ZN(n3166) );
  NOR2_X2 U2542 ( .A1(mem_3__0_), .A2(n2837), .ZN(n3165) );
  NOR3_X2 U2543 ( .A1(n3157), .A2(mem_2__0_), .A3(n3125), .ZN(n3167) );
  NOR3_X2 U2544 ( .A1(n3193), .A2(n3192), .A3(n3191), .ZN(n3198) );
  NOR3_X2 U2545 ( .A1(n3159), .A2(mem_26__0_), .A3(n3125), .ZN(n3193) );
  NOR2_X2 U2546 ( .A1(mem_27__0_), .A2(n2833), .ZN(n3191) );
  NOR2_X2 U2547 ( .A1(mem_28__0_), .A2(n2320), .ZN(n3192) );
  NOR3_X2 U2548 ( .A1(n3196), .A2(n3195), .A3(n3194), .ZN(n3197) );
  NOR2_X2 U2549 ( .A1(mem_30__0_), .A2(n2795), .ZN(n3194) );
  NOR2_X2 U2550 ( .A1(mem_29__0_), .A2(n2774), .ZN(n3195) );
  OAI21_X2 U2551 ( .B1(mem_31__0_), .B2(n2810), .A(n2759), .ZN(n3196) );
  NOR3_X2 U2552 ( .A1(n3188), .A2(n3187), .A3(n3186), .ZN(n3189) );
  NOR2_X2 U2553 ( .A1(mem_21__0_), .A2(n2774), .ZN(n3187) );
  NOR2_X2 U2554 ( .A1(mem_22__0_), .A2(n2793), .ZN(n3186) );
  OAI21_X1 U2555 ( .B1(mem_23__0_), .B2(n2810), .A(n2754), .ZN(n3188) );
  NOR3_X2 U2556 ( .A1(n3185), .A2(n3184), .A3(n3183), .ZN(n3190) );
  NOR3_X2 U2557 ( .A1(n3159), .A2(mem_18__0_), .A3(n3125), .ZN(n3185) );
  NOR2_X1 U2558 ( .A1(mem_19__0_), .A2(n2838), .ZN(n3183) );
  NOR2_X2 U2559 ( .A1(mem_20__0_), .A2(n2321), .ZN(n3184) );
  NOR2_X2 U2560 ( .A1(mem_12__2_), .A2(n2320), .ZN(n3269) );
  NOR2_X2 U2561 ( .A1(mem_11__2_), .A2(n2837), .ZN(n3268) );
  NOR3_X2 U2562 ( .A1(n3158), .A2(mem_10__2_), .A3(n3125), .ZN(n3270) );
  NOR3_X2 U2563 ( .A1(n3273), .A2(n3272), .A3(n3271), .ZN(n3274) );
  NOR2_X2 U2564 ( .A1(mem_13__2_), .A2(n2774), .ZN(n3272) );
  NOR2_X2 U2565 ( .A1(mem_14__2_), .A2(n2793), .ZN(n3271) );
  OAI21_X1 U2566 ( .B1(mem_15__2_), .B2(n2810), .A(n2758), .ZN(n3273) );
  NOR2_X2 U2567 ( .A1(mem_6__2_), .A2(n2793), .ZN(n3263) );
  NOR2_X2 U2568 ( .A1(mem_5__2_), .A2(n2774), .ZN(n3264) );
  NOR2_X2 U2569 ( .A1(mem_3__2_), .A2(n2837), .ZN(n3260) );
  NOR3_X2 U2570 ( .A1(n3159), .A2(mem_2__2_), .A3(n3125), .ZN(n3262) );
  NOR3_X2 U2571 ( .A1(n3291), .A2(n3290), .A3(n3289), .ZN(n3292) );
  NOR2_X2 U2572 ( .A1(mem_30__2_), .A2(n2791), .ZN(n3289) );
  NOR2_X2 U2573 ( .A1(mem_29__2_), .A2(n2775), .ZN(n3290) );
  OAI21_X2 U2574 ( .B1(mem_31__2_), .B2(n2810), .A(n2759), .ZN(n3291) );
  NOR3_X2 U2575 ( .A1(n3288), .A2(n3287), .A3(n3286), .ZN(n3293) );
  NOR3_X2 U2576 ( .A1(n3158), .A2(mem_26__2_), .A3(n3125), .ZN(n3288) );
  NOR2_X2 U2577 ( .A1(mem_27__2_), .A2(n2832), .ZN(n3286) );
  NOR3_X2 U2578 ( .A1(n3283), .A2(n3282), .A3(n3281), .ZN(n3284) );
  NOR2_X2 U2579 ( .A1(mem_21__2_), .A2(n2774), .ZN(n3282) );
  NOR2_X2 U2580 ( .A1(mem_22__2_), .A2(n2793), .ZN(n3281) );
  OAI21_X1 U2581 ( .B1(mem_23__2_), .B2(n2810), .A(n2758), .ZN(n3283) );
  NOR3_X2 U2582 ( .A1(n3280), .A2(n3279), .A3(n3278), .ZN(n3285) );
  NOR3_X2 U2583 ( .A1(n3159), .A2(mem_18__2_), .A3(n3125), .ZN(n3280) );
  NOR2_X2 U2584 ( .A1(mem_19__2_), .A2(n2837), .ZN(n3278) );
  NOR2_X2 U2585 ( .A1(mem_20__2_), .A2(n2320), .ZN(n3279) );
  NOR2_X2 U2586 ( .A1(mem_12__3_), .A2(n2318), .ZN(n3309) );
  NOR2_X2 U2587 ( .A1(mem_11__3_), .A2(n2837), .ZN(n3308) );
  NOR3_X2 U2588 ( .A1(n3158), .A2(mem_10__3_), .A3(n3125), .ZN(n3310) );
  NOR3_X2 U2589 ( .A1(n3313), .A2(n3312), .A3(n3311), .ZN(n3314) );
  NOR2_X2 U2590 ( .A1(mem_13__3_), .A2(n2775), .ZN(n3312) );
  NOR2_X2 U2591 ( .A1(mem_14__3_), .A2(n2794), .ZN(n3311) );
  OAI21_X2 U2592 ( .B1(mem_15__3_), .B2(n2809), .A(n2757), .ZN(n3313) );
  OAI21_X1 U2593 ( .B1(mem_7__3_), .B2(n2809), .A(n2759), .ZN(n3305) );
  NOR2_X2 U2594 ( .A1(mem_6__3_), .A2(n2794), .ZN(n3303) );
  NOR2_X2 U2595 ( .A1(mem_5__3_), .A2(n2775), .ZN(n3304) );
  NOR2_X2 U2596 ( .A1(mem_3__3_), .A2(n2836), .ZN(n3300) );
  NOR3_X2 U2597 ( .A1(n3159), .A2(mem_2__3_), .A3(n3125), .ZN(n3302) );
  NOR2_X2 U2598 ( .A1(mem_30__3_), .A2(n2792), .ZN(n3329) );
  NOR2_X2 U2599 ( .A1(mem_29__3_), .A2(n2775), .ZN(n3330) );
  OAI21_X2 U2600 ( .B1(mem_31__3_), .B2(n2809), .A(n2759), .ZN(n3331) );
  NOR3_X2 U2601 ( .A1(n3323), .A2(n3322), .A3(n3321), .ZN(n3324) );
  NOR2_X2 U2602 ( .A1(mem_21__3_), .A2(n2775), .ZN(n3322) );
  NOR2_X2 U2603 ( .A1(mem_22__3_), .A2(n2794), .ZN(n3321) );
  OAI21_X2 U2604 ( .B1(mem_23__3_), .B2(n2809), .A(n2757), .ZN(n3323) );
  NOR3_X2 U2605 ( .A1(n3320), .A2(n3319), .A3(n3318), .ZN(n3325) );
  NOR3_X2 U2606 ( .A1(n3159), .A2(mem_18__3_), .A3(n3126), .ZN(n3320) );
  NOR2_X1 U2607 ( .A1(mem_19__3_), .A2(n2832), .ZN(n3318) );
  NOR2_X2 U2608 ( .A1(mem_20__3_), .A2(n2319), .ZN(n3319) );
  NOR2_X2 U2609 ( .A1(mem_12__4_), .A2(n2321), .ZN(n3349) );
  NOR2_X1 U2610 ( .A1(mem_11__4_), .A2(n2832), .ZN(n3348) );
  NOR3_X2 U2611 ( .A1(n3158), .A2(mem_10__4_), .A3(n3126), .ZN(n3350) );
  NOR3_X2 U2612 ( .A1(n3353), .A2(n3352), .A3(n3351), .ZN(n3354) );
  NOR2_X2 U2613 ( .A1(mem_14__4_), .A2(n2791), .ZN(n3351) );
  NOR2_X2 U2614 ( .A1(mem_13__4_), .A2(n2775), .ZN(n3352) );
  OAI21_X1 U2615 ( .B1(mem_15__4_), .B2(n2809), .A(n2754), .ZN(n3353) );
  OAI21_X1 U2616 ( .B1(mem_7__4_), .B2(n2809), .A(n2754), .ZN(n3345) );
  NOR2_X2 U2617 ( .A1(mem_5__4_), .A2(n2775), .ZN(n3344) );
  NOR2_X2 U2618 ( .A1(mem_6__4_), .A2(n2791), .ZN(n3343) );
  NOR2_X1 U2619 ( .A1(mem_3__4_), .A2(n2832), .ZN(n3340) );
  NOR3_X2 U2620 ( .A1(n3159), .A2(mem_2__4_), .A3(n3126), .ZN(n3342) );
  NOR2_X2 U2621 ( .A1(mem_30__4_), .A2(n2791), .ZN(n3369) );
  NOR2_X2 U2622 ( .A1(mem_29__4_), .A2(n2775), .ZN(n3370) );
  OAI21_X2 U2623 ( .B1(mem_31__4_), .B2(n2809), .A(n2754), .ZN(n3371) );
  NOR3_X2 U2624 ( .A1(n3368), .A2(n3367), .A3(n3366), .ZN(n3373) );
  NOR3_X2 U2625 ( .A1(n3158), .A2(mem_26__4_), .A3(n3126), .ZN(n3368) );
  NOR2_X2 U2626 ( .A1(mem_28__4_), .A2(n2318), .ZN(n3367) );
  NOR3_X2 U2627 ( .A1(n3360), .A2(n3359), .A3(n3358), .ZN(n3365) );
  NOR3_X2 U2628 ( .A1(n3159), .A2(mem_18__4_), .A3(n3126), .ZN(n3360) );
  NOR2_X1 U2629 ( .A1(mem_19__4_), .A2(n2832), .ZN(n3358) );
  NOR2_X2 U2630 ( .A1(mem_20__4_), .A2(n2320), .ZN(n3359) );
  NOR2_X1 U2631 ( .A1(mem_11__5_), .A2(n2832), .ZN(n3388) );
  NOR3_X2 U2632 ( .A1(n3158), .A2(mem_10__5_), .A3(n3126), .ZN(n3390) );
  NOR3_X2 U2633 ( .A1(n3393), .A2(n3392), .A3(n3391), .ZN(n3394) );
  NOR2_X2 U2634 ( .A1(mem_14__5_), .A2(n2791), .ZN(n3391) );
  NOR2_X2 U2635 ( .A1(mem_13__5_), .A2(n2775), .ZN(n3392) );
  OAI21_X1 U2636 ( .B1(mem_15__5_), .B2(n2809), .A(n2754), .ZN(n3393) );
  OAI21_X2 U2637 ( .B1(mem_7__5_), .B2(n2809), .A(n2754), .ZN(n3385) );
  NOR2_X2 U2638 ( .A1(mem_5__5_), .A2(n2775), .ZN(n3384) );
  NOR2_X2 U2639 ( .A1(mem_6__5_), .A2(n2791), .ZN(n3383) );
  NOR2_X2 U2640 ( .A1(mem_4__5_), .A2(n2318), .ZN(n3381) );
  NOR2_X1 U2641 ( .A1(mem_3__5_), .A2(n2832), .ZN(n3380) );
  NOR3_X2 U2642 ( .A1(n3159), .A2(mem_2__5_), .A3(n3126), .ZN(n3382) );
  NOR2_X2 U2643 ( .A1(mem_30__5_), .A2(n2791), .ZN(n3409) );
  NOR2_X2 U2644 ( .A1(mem_29__5_), .A2(n2775), .ZN(n3410) );
  OAI21_X2 U2645 ( .B1(mem_31__5_), .B2(n2809), .A(n2754), .ZN(n3411) );
  NOR2_X2 U2646 ( .A1(mem_22__5_), .A2(n2791), .ZN(n3401) );
  NOR2_X2 U2647 ( .A1(mem_21__5_), .A2(n2775), .ZN(n3402) );
  OAI21_X2 U2648 ( .B1(mem_23__5_), .B2(n2809), .A(n2754), .ZN(n3403) );
  NOR3_X2 U2649 ( .A1(n3400), .A2(n3399), .A3(n3398), .ZN(n3405) );
  NOR3_X2 U2650 ( .A1(n3159), .A2(mem_18__5_), .A3(n3126), .ZN(n3400) );
  NOR2_X1 U2651 ( .A1(mem_19__5_), .A2(n2832), .ZN(n3398) );
  NOR2_X2 U2652 ( .A1(mem_20__5_), .A2(n2318), .ZN(n3399) );
  NOR2_X2 U2653 ( .A1(mem_12__6_), .A2(n2320), .ZN(n3429) );
  NOR2_X1 U2654 ( .A1(mem_11__6_), .A2(n2832), .ZN(n3428) );
  NOR3_X2 U2655 ( .A1(n3158), .A2(mem_10__6_), .A3(n3126), .ZN(n3430) );
  NOR2_X2 U2656 ( .A1(mem_14__6_), .A2(n2791), .ZN(n3431) );
  NOR2_X2 U2657 ( .A1(mem_13__6_), .A2(n2776), .ZN(n3432) );
  OAI21_X2 U2658 ( .B1(mem_15__6_), .B2(n2808), .A(n2754), .ZN(n3433) );
  OAI21_X2 U2659 ( .B1(mem_7__6_), .B2(n2808), .A(n2754), .ZN(n3425) );
  NOR2_X2 U2660 ( .A1(mem_5__6_), .A2(n2776), .ZN(n3424) );
  NOR2_X2 U2661 ( .A1(mem_6__6_), .A2(n2791), .ZN(n3423) );
  NOR2_X2 U2662 ( .A1(mem_4__6_), .A2(n2320), .ZN(n3421) );
  NOR2_X1 U2663 ( .A1(mem_3__6_), .A2(n2832), .ZN(n3420) );
  NOR3_X2 U2664 ( .A1(n3157), .A2(mem_2__6_), .A3(n3126), .ZN(n3422) );
  NOR2_X2 U2665 ( .A1(mem_30__6_), .A2(n2791), .ZN(n3449) );
  NOR2_X2 U2666 ( .A1(mem_29__6_), .A2(n2776), .ZN(n3450) );
  NOR3_X2 U2667 ( .A1(n3158), .A2(mem_26__6_), .A3(n3127), .ZN(n3448) );
  NOR2_X2 U2668 ( .A1(mem_28__6_), .A2(n2320), .ZN(n3447) );
  NOR2_X2 U2669 ( .A1(mem_22__6_), .A2(n2791), .ZN(n3441) );
  NOR2_X2 U2670 ( .A1(mem_21__6_), .A2(n2776), .ZN(n3442) );
  OAI21_X2 U2671 ( .B1(mem_23__6_), .B2(n2808), .A(n2754), .ZN(n3443) );
  NOR2_X2 U2672 ( .A1(mem_13__7_), .A2(n2776), .ZN(n3472) );
  NOR2_X2 U2673 ( .A1(mem_14__7_), .A2(n2792), .ZN(n3471) );
  OAI21_X2 U2674 ( .B1(mem_15__7_), .B2(n2808), .A(n2755), .ZN(n3473) );
  NOR3_X2 U2675 ( .A1(n3470), .A2(n3469), .A3(n3468), .ZN(n3475) );
  NOR3_X2 U2676 ( .A1(n3158), .A2(mem_10__7_), .A3(n3127), .ZN(n3470) );
  NOR2_X1 U2677 ( .A1(mem_11__7_), .A2(n2833), .ZN(n3468) );
  NOR2_X2 U2678 ( .A1(mem_12__7_), .A2(n2320), .ZN(n3469) );
  NOR2_X2 U2679 ( .A1(mem_4__7_), .A2(n2318), .ZN(n3461) );
  NOR2_X1 U2680 ( .A1(mem_3__7_), .A2(n2833), .ZN(n3460) );
  NOR3_X2 U2681 ( .A1(n3158), .A2(mem_2__7_), .A3(n3127), .ZN(n3462) );
  NOR2_X2 U2682 ( .A1(mem_5__7_), .A2(n2776), .ZN(n3464) );
  NOR2_X2 U2683 ( .A1(mem_6__7_), .A2(n2795), .ZN(n3463) );
  OAI21_X2 U2684 ( .B1(mem_7__7_), .B2(n2808), .A(n2755), .ZN(n3465) );
  NOR3_X2 U2685 ( .A1(n3488), .A2(n3487), .A3(n3486), .ZN(n3493) );
  NOR3_X2 U2686 ( .A1(n3157), .A2(mem_26__7_), .A3(n3127), .ZN(n3488) );
  NOR2_X2 U2687 ( .A1(mem_28__7_), .A2(n2320), .ZN(n3487) );
  NOR3_X2 U2688 ( .A1(n3491), .A2(n3490), .A3(n3489), .ZN(n3492) );
  OAI21_X2 U2689 ( .B1(mem_31__7_), .B2(n2808), .A(n2755), .ZN(n3491) );
  NOR2_X2 U2690 ( .A1(mem_30__7_), .A2(n2795), .ZN(n3489) );
  NOR2_X2 U2691 ( .A1(mem_29__7_), .A2(n2776), .ZN(n3490) );
  NOR3_X2 U2692 ( .A1(n3480), .A2(n3479), .A3(n3478), .ZN(n3485) );
  NOR3_X2 U2693 ( .A1(n3158), .A2(mem_18__7_), .A3(n3127), .ZN(n3480) );
  NOR2_X1 U2694 ( .A1(mem_19__7_), .A2(n2833), .ZN(n3478) );
  NOR2_X2 U2695 ( .A1(mem_20__7_), .A2(n2319), .ZN(n3479) );
  NOR3_X2 U2696 ( .A1(n3483), .A2(n3482), .A3(n3481), .ZN(n3484) );
  OAI21_X2 U2697 ( .B1(mem_23__7_), .B2(n2808), .A(n2755), .ZN(n3483) );
  NOR2_X2 U2698 ( .A1(mem_22__7_), .A2(n2792), .ZN(n3481) );
  NOR2_X2 U2699 ( .A1(mem_21__7_), .A2(n2776), .ZN(n3482) );
  NOR2_X2 U2700 ( .A1(mem_12__8_), .A2(n2319), .ZN(n3509) );
  NOR2_X1 U2701 ( .A1(mem_11__8_), .A2(n2833), .ZN(n3508) );
  NOR3_X2 U2702 ( .A1(n3157), .A2(mem_10__8_), .A3(n3127), .ZN(n3510) );
  NOR2_X2 U2703 ( .A1(mem_13__8_), .A2(n2776), .ZN(n3512) );
  NOR2_X2 U2704 ( .A1(mem_14__8_), .A2(n2793), .ZN(n3511) );
  OAI21_X2 U2705 ( .B1(mem_15__8_), .B2(n2808), .A(n2755), .ZN(n3513) );
  NOR2_X2 U2706 ( .A1(mem_4__8_), .A2(n2320), .ZN(n3501) );
  NOR2_X1 U2707 ( .A1(mem_3__8_), .A2(n2833), .ZN(n3500) );
  NOR3_X2 U2708 ( .A1(n3157), .A2(mem_2__8_), .A3(n3127), .ZN(n3502) );
  NOR2_X2 U2709 ( .A1(mem_5__8_), .A2(n2776), .ZN(n3504) );
  NOR2_X2 U2710 ( .A1(mem_6__8_), .A2(n2794), .ZN(n3503) );
  OAI21_X2 U2711 ( .B1(mem_7__8_), .B2(n2808), .A(n2755), .ZN(n3505) );
  INV_X4 U2712 ( .A(n2823), .ZN(n2815) );
  NOR3_X2 U2713 ( .A1(n3531), .A2(n3530), .A3(n3529), .ZN(n3532) );
  OAI21_X2 U2714 ( .B1(mem_31__8_), .B2(n2808), .A(n2755), .ZN(n3531) );
  NOR2_X2 U2715 ( .A1(mem_30__8_), .A2(n2792), .ZN(n3529) );
  NOR2_X2 U2716 ( .A1(mem_29__8_), .A2(n2776), .ZN(n3530) );
  NOR3_X2 U2717 ( .A1(n3520), .A2(n3519), .A3(n3518), .ZN(n3525) );
  NOR3_X2 U2718 ( .A1(n3157), .A2(mem_18__8_), .A3(n3127), .ZN(n3520) );
  NOR2_X1 U2719 ( .A1(mem_19__8_), .A2(n2833), .ZN(n3518) );
  NOR2_X2 U2720 ( .A1(mem_20__8_), .A2(n2321), .ZN(n3519) );
  NOR3_X2 U2721 ( .A1(n3523), .A2(n3522), .A3(n3521), .ZN(n3524) );
  OAI21_X2 U2722 ( .B1(mem_23__8_), .B2(n2808), .A(n2755), .ZN(n3523) );
  NOR2_X2 U2723 ( .A1(mem_22__8_), .A2(n2795), .ZN(n3521) );
  NOR2_X2 U2724 ( .A1(mem_21__8_), .A2(n2776), .ZN(n3522) );
  NOR2_X2 U2725 ( .A1(mem_12__9_), .A2(n2321), .ZN(n3549) );
  NOR2_X1 U2726 ( .A1(mem_11__9_), .A2(n2833), .ZN(n3548) );
  NOR3_X2 U2727 ( .A1(n3157), .A2(mem_10__9_), .A3(n3127), .ZN(n3550) );
  NOR3_X2 U2728 ( .A1(n3553), .A2(n3552), .A3(n3551), .ZN(n3554) );
  NOR2_X2 U2729 ( .A1(mem_14__9_), .A2(n2793), .ZN(n3551) );
  NOR2_X2 U2730 ( .A1(mem_13__9_), .A2(n2777), .ZN(n3552) );
  OAI21_X2 U2731 ( .B1(mem_15__9_), .B2(n2807), .A(n2755), .ZN(n3553) );
  OAI21_X2 U2732 ( .B1(mem_7__9_), .B2(n2807), .A(n2755), .ZN(n3545) );
  NOR2_X2 U2733 ( .A1(mem_5__9_), .A2(n2776), .ZN(n3544) );
  NOR2_X2 U2734 ( .A1(mem_6__9_), .A2(n2791), .ZN(n3543) );
  NOR2_X2 U2735 ( .A1(mem_4__9_), .A2(n2319), .ZN(n3541) );
  NOR2_X1 U2736 ( .A1(mem_3__9_), .A2(n2833), .ZN(n3540) );
  NOR3_X2 U2737 ( .A1(n3157), .A2(mem_2__9_), .A3(n3127), .ZN(n3542) );
  NOR3_X2 U2738 ( .A1(n3571), .A2(n3570), .A3(n3569), .ZN(n3572) );
  NOR2_X2 U2739 ( .A1(mem_30__9_), .A2(n2791), .ZN(n3569) );
  NOR2_X2 U2740 ( .A1(mem_29__9_), .A2(n2777), .ZN(n3570) );
  OAI21_X2 U2741 ( .B1(mem_31__9_), .B2(n2807), .A(n2755), .ZN(n3571) );
  NOR3_X2 U2742 ( .A1(n3157), .A2(mem_26__9_), .A3(n3128), .ZN(n3568) );
  NOR2_X2 U2743 ( .A1(mem_28__9_), .A2(n2318), .ZN(n3567) );
  NOR3_X2 U2744 ( .A1(n3563), .A2(n3562), .A3(n3561), .ZN(n3564) );
  NOR2_X2 U2745 ( .A1(mem_22__9_), .A2(n2793), .ZN(n3561) );
  NOR2_X2 U2746 ( .A1(mem_21__9_), .A2(n2777), .ZN(n3562) );
  OAI21_X2 U2747 ( .B1(mem_23__9_), .B2(n2807), .A(n2755), .ZN(n3563) );
  NOR2_X2 U2748 ( .A1(mem_12__10_), .A2(n2318), .ZN(n3589) );
  NOR2_X1 U2749 ( .A1(mem_11__10_), .A2(n2834), .ZN(n3588) );
  NOR3_X2 U2750 ( .A1(n3157), .A2(mem_10__10_), .A3(n3128), .ZN(n3590) );
  NOR3_X2 U2751 ( .A1(n3593), .A2(n3592), .A3(n3591), .ZN(n3594) );
  NOR2_X2 U2752 ( .A1(mem_14__10_), .A2(n2792), .ZN(n3591) );
  NOR2_X2 U2753 ( .A1(mem_13__10_), .A2(n2777), .ZN(n3592) );
  OAI21_X2 U2754 ( .B1(mem_15__10_), .B2(n2807), .A(n2756), .ZN(n3593) );
  NOR2_X2 U2755 ( .A1(mem_4__10_), .A2(n2321), .ZN(n3581) );
  NOR2_X1 U2756 ( .A1(mem_3__10_), .A2(n2834), .ZN(n3580) );
  NOR3_X2 U2757 ( .A1(n3157), .A2(mem_2__10_), .A3(n3128), .ZN(n3582) );
  NOR3_X2 U2758 ( .A1(n3585), .A2(n3584), .A3(n3583), .ZN(n3586) );
  NOR2_X2 U2759 ( .A1(mem_6__10_), .A2(n2792), .ZN(n3583) );
  NOR2_X2 U2760 ( .A1(mem_5__10_), .A2(n2777), .ZN(n3584) );
  OAI21_X2 U2761 ( .B1(mem_7__10_), .B2(n2807), .A(n2756), .ZN(n3585) );
  NOR3_X2 U2762 ( .A1(n3611), .A2(n3610), .A3(n3609), .ZN(n3612) );
  NOR2_X2 U2763 ( .A1(mem_30__10_), .A2(n2792), .ZN(n3609) );
  NOR2_X2 U2764 ( .A1(mem_29__10_), .A2(n2777), .ZN(n3610) );
  OAI21_X2 U2765 ( .B1(mem_31__10_), .B2(n2807), .A(n2756), .ZN(n3611) );
  NOR3_X2 U2766 ( .A1(n3157), .A2(mem_26__10_), .A3(n3128), .ZN(n3608) );
  NOR2_X2 U2767 ( .A1(mem_27__10_), .A2(n2834), .ZN(n3606) );
  NOR3_X2 U2768 ( .A1(n3603), .A2(n3602), .A3(n3601), .ZN(n3604) );
  NOR2_X2 U2769 ( .A1(mem_22__10_), .A2(n2792), .ZN(n3601) );
  NOR2_X2 U2770 ( .A1(mem_21__10_), .A2(n2777), .ZN(n3602) );
  OAI21_X2 U2771 ( .B1(mem_23__10_), .B2(n2807), .A(n2756), .ZN(n3603) );
  NOR3_X2 U2772 ( .A1(n3600), .A2(n3599), .A3(n3598), .ZN(n3605) );
  NOR3_X2 U2773 ( .A1(n3157), .A2(mem_18__10_), .A3(n3128), .ZN(n3600) );
  NOR2_X1 U2774 ( .A1(mem_19__10_), .A2(n2834), .ZN(n3598) );
  NOR2_X2 U2775 ( .A1(mem_12__11_), .A2(n2321), .ZN(n3629) );
  NOR2_X1 U2776 ( .A1(mem_11__11_), .A2(n2834), .ZN(n3628) );
  NOR3_X2 U2777 ( .A1(n3158), .A2(mem_10__11_), .A3(n3128), .ZN(n3630) );
  NOR3_X2 U2778 ( .A1(n3633), .A2(n3632), .A3(n3631), .ZN(n3634) );
  NOR2_X2 U2779 ( .A1(mem_14__11_), .A2(n2792), .ZN(n3631) );
  NOR2_X2 U2780 ( .A1(mem_13__11_), .A2(n2777), .ZN(n3632) );
  OAI21_X2 U2781 ( .B1(mem_15__11_), .B2(n2807), .A(n2756), .ZN(n3633) );
  OAI21_X2 U2782 ( .B1(mem_7__11_), .B2(n2807), .A(n2756), .ZN(n3625) );
  NOR2_X2 U2783 ( .A1(mem_5__11_), .A2(n2777), .ZN(n3624) );
  NOR2_X2 U2784 ( .A1(mem_6__11_), .A2(n2792), .ZN(n3623) );
  NOR2_X2 U2785 ( .A1(mem_4__11_), .A2(n2319), .ZN(n3621) );
  NOR2_X1 U2786 ( .A1(mem_3__11_), .A2(n2834), .ZN(n3620) );
  NOR3_X2 U2787 ( .A1(n3157), .A2(mem_2__11_), .A3(n3128), .ZN(n3622) );
  NOR3_X2 U2788 ( .A1(n3157), .A2(mem_26__11_), .A3(n3128), .ZN(n3648) );
  NOR2_X2 U2789 ( .A1(mem_27__11_), .A2(n2834), .ZN(n3646) );
  NOR2_X2 U2790 ( .A1(mem_28__11_), .A2(n2319), .ZN(n3647) );
  NOR3_X2 U2791 ( .A1(n3643), .A2(n3642), .A3(n3641), .ZN(n3644) );
  NOR2_X2 U2792 ( .A1(mem_22__11_), .A2(n2792), .ZN(n3641) );
  NOR2_X2 U2793 ( .A1(mem_21__11_), .A2(n2777), .ZN(n3642) );
  OAI21_X2 U2794 ( .B1(mem_23__11_), .B2(n2807), .A(n2756), .ZN(n3643) );
  NOR3_X2 U2795 ( .A1(n3640), .A2(n3639), .A3(n3638), .ZN(n3645) );
  NOR3_X2 U2796 ( .A1(n3157), .A2(mem_18__11_), .A3(n3128), .ZN(n3640) );
  NOR2_X1 U2797 ( .A1(mem_19__11_), .A2(n2834), .ZN(n3638) );
  NOR2_X2 U2798 ( .A1(mem_12__13_), .A2(n2320), .ZN(n3710) );
  NOR2_X1 U2799 ( .A1(mem_11__13_), .A2(n2834), .ZN(n3709) );
  NOR3_X2 U2800 ( .A1(n3157), .A2(mem_10__13_), .A3(n3128), .ZN(n3711) );
  NOR3_X2 U2801 ( .A1(n3714), .A2(n3713), .A3(n3712), .ZN(n3715) );
  NOR2_X2 U2802 ( .A1(mem_14__13_), .A2(n2792), .ZN(n3712) );
  NOR2_X2 U2803 ( .A1(mem_13__13_), .A2(n2777), .ZN(n3713) );
  OAI21_X2 U2804 ( .B1(mem_15__13_), .B2(n2806), .A(n2756), .ZN(n3714) );
  NOR2_X2 U2805 ( .A1(mem_4__13_), .A2(n2321), .ZN(n3702) );
  NOR2_X1 U2806 ( .A1(mem_3__13_), .A2(n2834), .ZN(n3701) );
  NOR3_X2 U2807 ( .A1(n3158), .A2(mem_2__13_), .A3(n3129), .ZN(n3703) );
  NOR3_X2 U2808 ( .A1(n3706), .A2(n3705), .A3(n3704), .ZN(n3707) );
  NOR2_X2 U2809 ( .A1(mem_6__13_), .A2(n2792), .ZN(n3704) );
  NOR2_X2 U2810 ( .A1(mem_5__13_), .A2(n2777), .ZN(n3705) );
  OAI21_X2 U2811 ( .B1(mem_7__13_), .B2(n2806), .A(n2756), .ZN(n3706) );
  NOR3_X2 U2812 ( .A1(n3732), .A2(n3731), .A3(n3730), .ZN(n3733) );
  NOR2_X2 U2813 ( .A1(mem_30__13_), .A2(n2792), .ZN(n3730) );
  NOR2_X2 U2814 ( .A1(mem_29__13_), .A2(n2778), .ZN(n3731) );
  OAI21_X2 U2815 ( .B1(mem_31__13_), .B2(n2806), .A(n2756), .ZN(n3732) );
  NOR3_X2 U2816 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3725) );
  NOR2_X2 U2817 ( .A1(mem_22__13_), .A2(n2792), .ZN(n3722) );
  NOR2_X2 U2818 ( .A1(mem_21__13_), .A2(n2778), .ZN(n3723) );
  OAI21_X2 U2819 ( .B1(mem_23__13_), .B2(n2806), .A(n2756), .ZN(n3724) );
  NOR3_X2 U2820 ( .A1(n3721), .A2(n3720), .A3(n3719), .ZN(n3726) );
  NOR3_X2 U2821 ( .A1(n3157), .A2(mem_18__13_), .A3(n3128), .ZN(n3721) );
  NOR2_X1 U2822 ( .A1(mem_19__13_), .A2(n2834), .ZN(n3719) );
  NOR2_X2 U2823 ( .A1(mem_20__13_), .A2(n2318), .ZN(n3720) );
  NOR2_X2 U2824 ( .A1(mem_12__14_), .A2(n2319), .ZN(n3750) );
  NOR2_X2 U2825 ( .A1(mem_11__14_), .A2(n2837), .ZN(n3749) );
  NOR3_X2 U2826 ( .A1(n3157), .A2(mem_10__14_), .A3(n3129), .ZN(n3751) );
  NOR3_X2 U2827 ( .A1(n3754), .A2(n3753), .A3(n3752), .ZN(n3755) );
  NOR2_X2 U2828 ( .A1(mem_13__14_), .A2(n2778), .ZN(n3753) );
  NOR2_X2 U2829 ( .A1(mem_14__14_), .A2(n2793), .ZN(n3752) );
  OAI21_X2 U2830 ( .B1(mem_15__14_), .B2(n2806), .A(n2757), .ZN(n3754) );
  OAI21_X2 U2831 ( .B1(mem_7__14_), .B2(n2806), .A(n2757), .ZN(n3746) );
  NOR2_X2 U2832 ( .A1(mem_6__14_), .A2(n2793), .ZN(n3744) );
  NOR2_X2 U2833 ( .A1(mem_5__14_), .A2(n2776), .ZN(n3745) );
  NOR2_X2 U2834 ( .A1(mem_4__14_), .A2(n2320), .ZN(n3742) );
  NOR2_X2 U2835 ( .A1(mem_3__14_), .A2(n2837), .ZN(n3741) );
  NOR3_X2 U2836 ( .A1(n3158), .A2(mem_2__14_), .A3(n3129), .ZN(n3743) );
  NOR3_X2 U2837 ( .A1(n3772), .A2(n3771), .A3(n3770), .ZN(n3773) );
  NOR2_X2 U2838 ( .A1(mem_29__14_), .A2(n2778), .ZN(n3771) );
  NOR2_X2 U2839 ( .A1(mem_30__14_), .A2(n2793), .ZN(n3770) );
  OAI21_X2 U2840 ( .B1(mem_31__14_), .B2(n2806), .A(n2757), .ZN(n3772) );
  NOR3_X2 U2841 ( .A1(n3157), .A2(mem_26__14_), .A3(n3129), .ZN(n3769) );
  NOR2_X2 U2842 ( .A1(mem_28__14_), .A2(n2318), .ZN(n3768) );
  NOR3_X2 U2843 ( .A1(n3764), .A2(n3763), .A3(n3762), .ZN(n3765) );
  NOR2_X2 U2844 ( .A1(mem_21__14_), .A2(n2775), .ZN(n3763) );
  NOR2_X2 U2845 ( .A1(mem_22__14_), .A2(n2793), .ZN(n3762) );
  OAI21_X2 U2846 ( .B1(mem_23__14_), .B2(n2806), .A(n2757), .ZN(n3764) );
  NOR3_X2 U2847 ( .A1(n3761), .A2(n3760), .A3(n3759), .ZN(n3766) );
  NOR3_X2 U2848 ( .A1(n3158), .A2(mem_18__14_), .A3(n3129), .ZN(n3761) );
  NOR2_X1 U2849 ( .A1(mem_19__14_), .A2(n2834), .ZN(n3759) );
  NOR2_X2 U2850 ( .A1(mem_20__14_), .A2(n2318), .ZN(n3760) );
  NOR2_X1 U2851 ( .A1(mem_11__15_), .A2(n2838), .ZN(n3789) );
  NOR3_X2 U2852 ( .A1(n3157), .A2(mem_10__15_), .A3(n3129), .ZN(n3791) );
  NOR3_X2 U2853 ( .A1(n3794), .A2(n3793), .A3(n3792), .ZN(n3795) );
  NOR2_X2 U2854 ( .A1(mem_13__15_), .A2(n2775), .ZN(n3793) );
  NOR2_X2 U2855 ( .A1(mem_14__15_), .A2(n2793), .ZN(n3792) );
  OAI21_X2 U2856 ( .B1(mem_15__15_), .B2(n2806), .A(n2757), .ZN(n3794) );
  OAI21_X2 U2857 ( .B1(mem_7__15_), .B2(n2806), .A(n2757), .ZN(n3786) );
  NOR2_X2 U2858 ( .A1(mem_6__15_), .A2(n2793), .ZN(n3784) );
  NOR2_X2 U2859 ( .A1(mem_5__15_), .A2(n2777), .ZN(n3785) );
  NOR2_X2 U2860 ( .A1(mem_4__15_), .A2(n2319), .ZN(n3782) );
  NOR2_X1 U2861 ( .A1(mem_3__15_), .A2(n2834), .ZN(n3781) );
  NOR3_X2 U2862 ( .A1(n3157), .A2(mem_2__15_), .A3(n3129), .ZN(n3783) );
  NOR3_X2 U2863 ( .A1(n3812), .A2(n3811), .A3(n3810), .ZN(n3813) );
  NOR2_X2 U2864 ( .A1(mem_29__15_), .A2(n2778), .ZN(n3811) );
  NOR2_X2 U2865 ( .A1(mem_30__15_), .A2(n2793), .ZN(n3810) );
  OAI21_X2 U2866 ( .B1(mem_31__15_), .B2(n2806), .A(n2757), .ZN(n3812) );
  NOR3_X2 U2867 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3805) );
  NOR2_X2 U2868 ( .A1(mem_21__15_), .A2(n2776), .ZN(n3803) );
  NOR2_X2 U2869 ( .A1(mem_22__15_), .A2(n2793), .ZN(n3802) );
  OAI21_X2 U2870 ( .B1(mem_23__15_), .B2(n2806), .A(n2757), .ZN(n3804) );
  NOR2_X2 U2871 ( .A1(mem_12__16_), .A2(n2321), .ZN(n3830) );
  NOR3_X2 U2872 ( .A1(n3156), .A2(mem_10__16_), .A3(n3130), .ZN(n3831) );
  NOR2_X2 U2873 ( .A1(mem_11__16_), .A2(n2836), .ZN(n3829) );
  NOR3_X2 U2874 ( .A1(n3834), .A2(n3833), .A3(n3832), .ZN(n3835) );
  NOR2_X2 U2875 ( .A1(mem_13__16_), .A2(n2776), .ZN(n3833) );
  NOR2_X2 U2876 ( .A1(mem_14__16_), .A2(n2793), .ZN(n3832) );
  OAI21_X2 U2877 ( .B1(mem_15__16_), .B2(n2806), .A(n2757), .ZN(n3834) );
  INV_X4 U2878 ( .A(n2774), .ZN(n2768) );
  NOR2_X2 U2879 ( .A1(mem_4__16_), .A2(n2321), .ZN(n3822) );
  NOR3_X2 U2880 ( .A1(n3156), .A2(mem_2__16_), .A3(n3129), .ZN(n3823) );
  NOR2_X1 U2881 ( .A1(mem_3__16_), .A2(n2834), .ZN(n3821) );
  INV_X4 U2882 ( .A(n2823), .ZN(n2816) );
  NOR3_X2 U2883 ( .A1(n3826), .A2(n3825), .A3(n3824), .ZN(n3827) );
  NOR2_X2 U2884 ( .A1(mem_5__16_), .A2(n2778), .ZN(n3825) );
  NOR2_X2 U2885 ( .A1(mem_6__16_), .A2(n2793), .ZN(n3824) );
  OAI21_X2 U2886 ( .B1(mem_7__16_), .B2(n2806), .A(n2757), .ZN(n3826) );
  NOR3_X2 U2887 ( .A1(n3852), .A2(n3851), .A3(n3850), .ZN(n3853) );
  NOR2_X2 U2888 ( .A1(mem_29__16_), .A2(n2778), .ZN(n3851) );
  NOR2_X2 U2889 ( .A1(mem_30__16_), .A2(n2793), .ZN(n3850) );
  NOR3_X2 U2890 ( .A1(n3844), .A2(n3843), .A3(n3842), .ZN(n3845) );
  NOR2_X2 U2891 ( .A1(mem_21__16_), .A2(n2777), .ZN(n3843) );
  NOR2_X2 U2892 ( .A1(mem_22__16_), .A2(n2793), .ZN(n3842) );
  OAI21_X2 U2893 ( .B1(mem_23__16_), .B2(n2806), .A(n2757), .ZN(n3844) );
  NOR2_X2 U2894 ( .A1(mem_12__17_), .A2(n2318), .ZN(n3870) );
  NOR3_X2 U2895 ( .A1(n3156), .A2(mem_10__17_), .A3(n3130), .ZN(n3871) );
  NOR2_X2 U2896 ( .A1(mem_11__17_), .A2(n2836), .ZN(n3869) );
  NOR3_X2 U2897 ( .A1(n3874), .A2(n3873), .A3(n3872), .ZN(n3875) );
  NOR2_X2 U2898 ( .A1(mem_13__17_), .A2(n2778), .ZN(n3873) );
  NOR2_X2 U2899 ( .A1(mem_14__17_), .A2(n2794), .ZN(n3872) );
  OAI21_X1 U2900 ( .B1(mem_15__17_), .B2(n2806), .A(n2758), .ZN(n3874) );
  NOR2_X2 U2901 ( .A1(mem_4__17_), .A2(n2318), .ZN(n3862) );
  NOR3_X2 U2902 ( .A1(n3156), .A2(mem_2__17_), .A3(n3130), .ZN(n3863) );
  NOR2_X2 U2903 ( .A1(mem_3__17_), .A2(n2836), .ZN(n3861) );
  NOR3_X2 U2904 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3867) );
  NOR2_X2 U2905 ( .A1(mem_5__17_), .A2(n2778), .ZN(n3865) );
  NOR2_X2 U2906 ( .A1(mem_6__17_), .A2(n2794), .ZN(n3864) );
  OAI21_X2 U2907 ( .B1(mem_7__17_), .B2(n2806), .A(n2758), .ZN(n3866) );
  NOR2_X2 U2908 ( .A1(mem_29__17_), .A2(n2778), .ZN(n3891) );
  NOR2_X2 U2909 ( .A1(mem_30__17_), .A2(n2794), .ZN(n3890) );
  NOR3_X2 U2910 ( .A1(n3881), .A2(n3880), .A3(n3879), .ZN(n3886) );
  NOR2_X2 U2911 ( .A1(mem_19__17_), .A2(n2836), .ZN(n3879) );
  NOR3_X2 U2912 ( .A1(n3156), .A2(mem_18__17_), .A3(n3130), .ZN(n3881) );
  NOR2_X2 U2913 ( .A1(mem_20__17_), .A2(n2320), .ZN(n3880) );
  NOR2_X2 U2914 ( .A1(mem_12__18_), .A2(n2321), .ZN(n3910) );
  NOR3_X2 U2915 ( .A1(n3156), .A2(mem_10__18_), .A3(n3130), .ZN(n3911) );
  NOR2_X2 U2916 ( .A1(mem_11__18_), .A2(n2836), .ZN(n3909) );
  INV_X4 U2917 ( .A(n2823), .ZN(n2818) );
  NOR2_X2 U2918 ( .A1(mem_4__18_), .A2(n2321), .ZN(n3902) );
  NOR3_X2 U2919 ( .A1(n3156), .A2(mem_2__18_), .A3(n3130), .ZN(n3903) );
  NOR2_X1 U2920 ( .A1(mem_3__18_), .A2(n2838), .ZN(n3901) );
  NOR3_X2 U2921 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3907) );
  NOR2_X2 U2922 ( .A1(mem_5__18_), .A2(n2778), .ZN(n3905) );
  NOR2_X2 U2923 ( .A1(mem_6__18_), .A2(n2794), .ZN(n3904) );
  OAI21_X2 U2924 ( .B1(mem_7__18_), .B2(n2806), .A(n2758), .ZN(n3906) );
  INV_X4 U2925 ( .A(n2825), .ZN(n2819) );
  NOR2_X2 U2926 ( .A1(mem_29__18_), .A2(n2778), .ZN(n3931) );
  NOR2_X2 U2927 ( .A1(mem_30__18_), .A2(n2794), .ZN(n3930) );
  NOR3_X2 U2928 ( .A1(n3929), .A2(n3928), .A3(n3927), .ZN(n3934) );
  NOR2_X2 U2929 ( .A1(mem_27__18_), .A2(n2838), .ZN(n3927) );
  NOR3_X2 U2930 ( .A1(n3156), .A2(mem_26__18_), .A3(n3130), .ZN(n3929) );
  NOR3_X2 U2931 ( .A1(n3921), .A2(n3920), .A3(n3919), .ZN(n3926) );
  NOR2_X1 U2932 ( .A1(mem_19__18_), .A2(n2838), .ZN(n3919) );
  NOR3_X2 U2933 ( .A1(n3156), .A2(mem_18__18_), .A3(n3130), .ZN(n3921) );
  NOR2_X2 U2934 ( .A1(mem_12__19_), .A2(n2320), .ZN(n3950) );
  NOR3_X2 U2935 ( .A1(n3156), .A2(mem_10__19_), .A3(n3131), .ZN(n3951) );
  NOR2_X1 U2936 ( .A1(mem_11__19_), .A2(n2838), .ZN(n3949) );
  NOR2_X2 U2937 ( .A1(mem_6__19_), .A2(n2794), .ZN(n3944) );
  OAI21_X2 U2938 ( .B1(mem_7__19_), .B2(n2805), .A(n2758), .ZN(n3946) );
  NOR2_X2 U2939 ( .A1(mem_5__19_), .A2(n2778), .ZN(n3945) );
  NOR3_X2 U2940 ( .A1(n3156), .A2(mem_2__19_), .A3(n3130), .ZN(n3943) );
  NOR2_X1 U2941 ( .A1(mem_3__19_), .A2(n2838), .ZN(n3941) );
  INV_X4 U2942 ( .A(n3123), .ZN(n3140) );
  NOR2_X2 U2943 ( .A1(mem_29__19_), .A2(n2778), .ZN(n3971) );
  NOR2_X2 U2944 ( .A1(mem_30__19_), .A2(n2794), .ZN(n3970) );
  NOR3_X2 U2945 ( .A1(n3969), .A2(n3968), .A3(n3967), .ZN(n3974) );
  NOR2_X2 U2946 ( .A1(mem_27__19_), .A2(n2838), .ZN(n3967) );
  NOR3_X2 U2947 ( .A1(n3156), .A2(mem_26__19_), .A3(n3131), .ZN(n3969) );
  NOR2_X2 U2948 ( .A1(mem_28__19_), .A2(n2318), .ZN(n3968) );
  NOR3_X2 U2949 ( .A1(n3964), .A2(n3963), .A3(n3962), .ZN(n3965) );
  NOR2_X2 U2950 ( .A1(mem_21__19_), .A2(n2778), .ZN(n3963) );
  OAI21_X2 U2951 ( .B1(mem_23__19_), .B2(n2805), .A(n2758), .ZN(n3964) );
  NOR2_X2 U2952 ( .A1(mem_22__19_), .A2(n2794), .ZN(n3962) );
  NOR3_X2 U2953 ( .A1(n3961), .A2(n3960), .A3(n3959), .ZN(n3966) );
  NOR2_X2 U2954 ( .A1(mem_19__19_), .A2(n2836), .ZN(n3959) );
  NOR3_X2 U2955 ( .A1(n3156), .A2(mem_18__19_), .A3(n3130), .ZN(n3961) );
  NOR2_X1 U2956 ( .A1(mem_13__20_), .A2(n2779), .ZN(n3993) );
  OAI21_X1 U2957 ( .B1(mem_15__20_), .B2(n2805), .A(n2759), .ZN(n3994) );
  NOR2_X2 U2958 ( .A1(mem_14__20_), .A2(n2795), .ZN(n3992) );
  NOR3_X2 U2959 ( .A1(n3156), .A2(mem_10__20_), .A3(n3131), .ZN(n3991) );
  NOR2_X2 U2960 ( .A1(mem_11__20_), .A2(n2835), .ZN(n3989) );
  NOR2_X1 U2961 ( .A1(mem_5__20_), .A2(n2779), .ZN(n3985) );
  OAI21_X2 U2962 ( .B1(mem_7__20_), .B2(n2805), .A(n2759), .ZN(n3986) );
  NOR2_X2 U2963 ( .A1(mem_6__20_), .A2(n2795), .ZN(n3984) );
  NOR3_X2 U2964 ( .A1(n3156), .A2(mem_2__20_), .A3(n3131), .ZN(n3983) );
  NOR2_X2 U2965 ( .A1(mem_4__20_), .A2(n2320), .ZN(n3982) );
  NOR2_X2 U2966 ( .A1(mem_3__20_), .A2(n2835), .ZN(n3981) );
  NOR2_X2 U2967 ( .A1(mem_30__20_), .A2(n2795), .ZN(n4010) );
  OAI21_X2 U2968 ( .B1(mem_31__20_), .B2(n2805), .A(n2759), .ZN(n4012) );
  NOR2_X1 U2969 ( .A1(mem_29__20_), .A2(n2779), .ZN(n4011) );
  NOR3_X2 U2970 ( .A1(n4009), .A2(n4008), .A3(n4007), .ZN(n4014) );
  NOR2_X2 U2971 ( .A1(mem_27__20_), .A2(n2835), .ZN(n4007) );
  NOR2_X2 U2972 ( .A1(mem_28__20_), .A2(n2321), .ZN(n4008) );
  NOR3_X2 U2973 ( .A1(n3156), .A2(mem_26__20_), .A3(n3131), .ZN(n4009) );
  NOR3_X2 U2974 ( .A1(n4001), .A2(n4000), .A3(n3999), .ZN(n4006) );
  NOR2_X2 U2975 ( .A1(mem_19__20_), .A2(n2835), .ZN(n3999) );
  NOR2_X2 U2976 ( .A1(mem_20__20_), .A2(n2319), .ZN(n4000) );
  NOR3_X2 U2977 ( .A1(n3156), .A2(mem_18__20_), .A3(n3131), .ZN(n4001) );
  NOR2_X1 U2978 ( .A1(mem_13__21_), .A2(n2779), .ZN(n4033) );
  OAI21_X1 U2979 ( .B1(mem_15__21_), .B2(n2805), .A(n2759), .ZN(n4034) );
  NOR2_X2 U2980 ( .A1(mem_14__21_), .A2(n2795), .ZN(n4032) );
  NOR3_X2 U2981 ( .A1(n3156), .A2(mem_10__21_), .A3(n3131), .ZN(n4031) );
  NOR2_X2 U2982 ( .A1(mem_12__21_), .A2(n2321), .ZN(n4030) );
  NOR2_X2 U2983 ( .A1(mem_11__21_), .A2(n2835), .ZN(n4029) );
  NOR2_X1 U2984 ( .A1(mem_5__21_), .A2(n2779), .ZN(n4025) );
  OAI21_X2 U2985 ( .B1(mem_7__21_), .B2(n2805), .A(n2759), .ZN(n4026) );
  NOR2_X2 U2986 ( .A1(mem_6__21_), .A2(n2795), .ZN(n4024) );
  NOR3_X2 U2987 ( .A1(n3156), .A2(mem_2__21_), .A3(n3131), .ZN(n4023) );
  NOR2_X2 U2988 ( .A1(mem_4__21_), .A2(n2319), .ZN(n4022) );
  NOR2_X2 U2989 ( .A1(mem_3__21_), .A2(n2835), .ZN(n4021) );
  INV_X4 U2990 ( .A(n3123), .ZN(n3141) );
  INV_X4 U2991 ( .A(n3123), .ZN(n3142) );
  NOR2_X2 U2992 ( .A1(mem_30__21_), .A2(n2795), .ZN(n4051) );
  NOR2_X1 U2993 ( .A1(mem_29__21_), .A2(n2779), .ZN(n4052) );
  NOR3_X2 U2994 ( .A1(n4049), .A2(n4048), .A3(n4047), .ZN(n4055) );
  NOR2_X2 U2995 ( .A1(mem_27__21_), .A2(n2835), .ZN(n4047) );
  NOR2_X2 U2996 ( .A1(mem_28__21_), .A2(n2318), .ZN(n4048) );
  NOR3_X2 U2997 ( .A1(n3156), .A2(mem_26__21_), .A3(n3131), .ZN(n4049) );
  NOR3_X2 U2998 ( .A1(n4044), .A2(n4043), .A3(n4042), .ZN(n4045) );
  NOR2_X2 U2999 ( .A1(mem_22__21_), .A2(n2795), .ZN(n4042) );
  OAI21_X2 U3000 ( .B1(mem_23__21_), .B2(n2805), .A(n2759), .ZN(n4044) );
  NOR2_X1 U3001 ( .A1(mem_21__21_), .A2(n2779), .ZN(n4043) );
  NOR3_X2 U3002 ( .A1(n4041), .A2(n4040), .A3(n4039), .ZN(n4046) );
  NOR2_X2 U3003 ( .A1(mem_19__21_), .A2(n2835), .ZN(n4039) );
  NOR2_X2 U3004 ( .A1(mem_20__21_), .A2(n2318), .ZN(n4040) );
  NOR3_X2 U3005 ( .A1(n3156), .A2(mem_18__21_), .A3(n3131), .ZN(n4041) );
  NOR2_X2 U3006 ( .A1(n3111), .A2(n3131), .ZN(n4083) );
  NOR2_X2 U3007 ( .A1(n4254), .A2(n4253), .ZN(n4257) );
  NOR2_X2 U3008 ( .A1(mem_11__25_), .A2(n2836), .ZN(n4253) );
  NOR2_X2 U3009 ( .A1(n4249), .A2(n4248), .ZN(n4252) );
  NOR2_X2 U3010 ( .A1(mem_14__25_), .A2(n2796), .ZN(n4248) );
  NOR2_X2 U3011 ( .A1(mem_2__25_), .A2(n3132), .ZN(n4241) );
  NOR2_X2 U3012 ( .A1(n4240), .A2(n4239), .ZN(n4243) );
  NOR2_X2 U3013 ( .A1(mem_4__25_), .A2(n2321), .ZN(n4240) );
  NOR2_X2 U3014 ( .A1(mem_3__25_), .A2(n2836), .ZN(n4239) );
  NOR2_X2 U3015 ( .A1(n4235), .A2(n4234), .ZN(n4238) );
  NOR2_X2 U3016 ( .A1(n2762), .A2(n4236), .ZN(n4237) );
  NOR2_X1 U3017 ( .A1(mem_5__25_), .A2(n2780), .ZN(n4235) );
  NOR2_X2 U3018 ( .A1(n2739), .A2(n3132), .ZN(n4285) );
  NOR2_X2 U3019 ( .A1(n4284), .A2(n4283), .ZN(n4287) );
  NOR2_X2 U3020 ( .A1(n2671), .A2(n2319), .ZN(n4284) );
  NOR2_X2 U3021 ( .A1(n4438), .A2(n4437), .ZN(n4441) );
  NOR2_X2 U3022 ( .A1(mem_14__28_), .A2(n2797), .ZN(n4437) );
  NOR2_X2 U3023 ( .A1(mem_13__28_), .A2(n2781), .ZN(n4438) );
  NOR2_X2 U3024 ( .A1(n4443), .A2(n4442), .ZN(n4446) );
  NOR2_X2 U3025 ( .A1(mem_12__28_), .A2(n2319), .ZN(n4443) );
  NOR2_X2 U3026 ( .A1(mem_7__28_), .A2(n2803), .ZN(n4425) );
  NOR2_X2 U3027 ( .A1(n4424), .A2(n4423), .ZN(n4427) );
  NOR2_X1 U3028 ( .A1(mem_5__28_), .A2(n2781), .ZN(n4424) );
  NOR2_X2 U3029 ( .A1(mem_6__28_), .A2(n2797), .ZN(n4423) );
  NOR2_X2 U3030 ( .A1(n4429), .A2(n4428), .ZN(n4432) );
  NOR2_X2 U3031 ( .A1(mem_4__28_), .A2(n2318), .ZN(n4429) );
  NOR2_X2 U3032 ( .A1(n2735), .A2(n3133), .ZN(n4474) );
  NOR2_X2 U3033 ( .A1(n4473), .A2(n4472), .ZN(n4476) );
  NOR2_X2 U3034 ( .A1(n2669), .A2(n2320), .ZN(n4473) );
  NOR2_X2 U3035 ( .A1(n4501), .A2(n4500), .ZN(n4504) );
  NOR2_X2 U3036 ( .A1(mem_14__29_), .A2(n2797), .ZN(n4500) );
  NOR2_X2 U3037 ( .A1(mem_13__29_), .A2(n2781), .ZN(n4501) );
  NOR2_X2 U3038 ( .A1(n4506), .A2(n4505), .ZN(n4509) );
  NOR2_X2 U3039 ( .A1(mem_12__29_), .A2(n2318), .ZN(n4506) );
  NOR2_X2 U3040 ( .A1(n4492), .A2(n4491), .ZN(n4495) );
  NOR2_X2 U3041 ( .A1(mem_4__29_), .A2(n2319), .ZN(n4492) );
  NOR2_X2 U3042 ( .A1(mem_3__29_), .A2(n2837), .ZN(n4491) );
  NOR2_X2 U3043 ( .A1(mem_2__29_), .A2(n3133), .ZN(n4493) );
  NOR2_X2 U3044 ( .A1(n4487), .A2(n4486), .ZN(n4490) );
  NOR2_X2 U3045 ( .A1(n2762), .A2(n4488), .ZN(n4489) );
  NOR2_X1 U3046 ( .A1(mem_5__29_), .A2(n2781), .ZN(n4487) );
  NOR2_X2 U3047 ( .A1(n4536), .A2(n4535), .ZN(n4539) );
  NOR2_X2 U3048 ( .A1(n2673), .A2(n2321), .ZN(n4536) );
  NOR2_X2 U3049 ( .A1(n2741), .A2(n3134), .ZN(n4537) );
  NOR2_X2 U3050 ( .A1(n4531), .A2(n4530), .ZN(n4534) );
  NOR2_X1 U3051 ( .A1(n2743), .A2(n2801), .ZN(n4532) );
  NOR2_X2 U3052 ( .A1(n4632), .A2(n4631), .ZN(n4635) );
  NOR2_X2 U3053 ( .A1(mem_12__31_), .A2(n2320), .ZN(n4632) );
  NOR2_X2 U3054 ( .A1(mem_11__31_), .A2(n2838), .ZN(n4631) );
  NOR2_X2 U3055 ( .A1(n4627), .A2(n4626), .ZN(n4630) );
  NOR2_X2 U3056 ( .A1(mem_14__31_), .A2(n2798), .ZN(n4626) );
  INV_X4 U3057 ( .A(n2774), .ZN(n2772) );
  INV_X4 U3058 ( .A(n3121), .ZN(n3146) );
  NOR2_X2 U3059 ( .A1(n4667), .A2(n4666), .ZN(n4670) );
  NOR2_X2 U3060 ( .A1(n2729), .A2(n2838), .ZN(n4666) );
  NOR2_X2 U3061 ( .A1(n2701), .A2(n2319), .ZN(n4667) );
  NOR2_X2 U3062 ( .A1(n2677), .A2(n3134), .ZN(n4668) );
  NOR2_X2 U3063 ( .A1(n4659), .A2(n4658), .ZN(n4663) );
  NOR2_X1 U3064 ( .A1(n2747), .A2(n2801), .ZN(n4661) );
  NOR2_X2 U3065 ( .A1(wData[0]), .A2(n2336), .ZN(n4692) );
  NOR2_X2 U3066 ( .A1(wData[1]), .A2(n2341), .ZN(n4740) );
  NOR2_X2 U3067 ( .A1(wData[2]), .A2(n2327), .ZN(n4788) );
  NOR2_X2 U3068 ( .A1(wData[3]), .A2(n2333), .ZN(n4836) );
  NOR2_X2 U3069 ( .A1(wData[4]), .A2(n2332), .ZN(n4884) );
  NOR2_X2 U3070 ( .A1(wData[5]), .A2(n2334), .ZN(n4932) );
  NOR2_X2 U3071 ( .A1(wData[6]), .A2(n2328), .ZN(n4980) );
  NOR2_X2 U3072 ( .A1(wData[7]), .A2(n2334), .ZN(n5028) );
  NOR2_X2 U3073 ( .A1(wData[8]), .A2(n2342), .ZN(n5076) );
  NOR2_X2 U3074 ( .A1(wData[9]), .A2(n2333), .ZN(n5124) );
  NOR2_X2 U3075 ( .A1(wData[11]), .A2(n2329), .ZN(n5223) );
  NOR2_X2 U3076 ( .A1(wData[12]), .A2(n2333), .ZN(n5271) );
  NOR2_X2 U3077 ( .A1(wData[13]), .A2(n2335), .ZN(n5319) );
  NOR2_X2 U3078 ( .A1(wData[14]), .A2(n2337), .ZN(n5367) );
  NOR2_X2 U3079 ( .A1(wData[15]), .A2(n2330), .ZN(n5415) );
  NOR2_X2 U3080 ( .A1(wData[16]), .A2(n2332), .ZN(n5463) );
  NOR2_X2 U3081 ( .A1(wData[17]), .A2(n2327), .ZN(n5511) );
  NOR2_X2 U3082 ( .A1(wData[18]), .A2(n2335), .ZN(n5559) );
  NOR2_X2 U3083 ( .A1(wData[19]), .A2(n2336), .ZN(n5607) );
  NOR2_X2 U3084 ( .A1(wData[20]), .A2(n2328), .ZN(n5655) );
  INV_X8 U3085 ( .A(n4691), .ZN(n5704) );
  NOR2_X2 U3086 ( .A1(wData[21]), .A2(n2334), .ZN(n5703) );
  NOR2_X2 U3087 ( .A1(mem_22__23_), .A2(n2873), .ZN(n5817) );
  NOR2_X1 U3088 ( .A1(mem_21__23_), .A2(n2869), .ZN(n5818) );
  NOR2_X2 U3089 ( .A1(mem_20__23_), .A2(n2853), .ZN(n5815) );
  NOR2_X2 U3090 ( .A1(mem_30__23_), .A2(n2873), .ZN(n5825) );
  NOR2_X2 U3091 ( .A1(mem_27__23_), .A2(n2856), .ZN(n5822) );
  NOR2_X2 U3092 ( .A1(mem_28__23_), .A2(n2853), .ZN(n5823) );
  NOR3_X2 U3093 ( .A1(n5801), .A2(n5800), .A3(n5799), .ZN(n5802) );
  OAI21_X2 U3094 ( .B1(mem_7__23_), .B2(n2862), .A(n2859), .ZN(n5801) );
  NOR2_X1 U3095 ( .A1(mem_5__23_), .A2(n2869), .ZN(n5800) );
  NOR2_X1 U3096 ( .A1(mem_6__23_), .A2(n2873), .ZN(n5799) );
  NOR3_X2 U3097 ( .A1(n5797), .A2(n5796), .A3(n5795), .ZN(n5803) );
  NOR2_X2 U3098 ( .A1(mem_4__23_), .A2(n2853), .ZN(n5796) );
  NOR2_X2 U3099 ( .A1(mem_3__23_), .A2(n2856), .ZN(n5795) );
  NOR2_X2 U3100 ( .A1(mem_13__23_), .A2(n2869), .ZN(n5808) );
  NOR2_X2 U3101 ( .A1(mem_27__24_), .A2(n2856), .ZN(n5862) );
  NOR2_X2 U3102 ( .A1(mem_28__24_), .A2(n2853), .ZN(n5863) );
  NOR2_X2 U3103 ( .A1(mem_29__24_), .A2(n2869), .ZN(n5866) );
  NOR2_X1 U3104 ( .A1(mem_30__24_), .A2(n2873), .ZN(n5865) );
  NOR2_X2 U3105 ( .A1(mem_20__24_), .A2(n2853), .ZN(n5855) );
  NOR2_X2 U3106 ( .A1(mem_21__24_), .A2(n2869), .ZN(n5858) );
  NOR2_X1 U3107 ( .A1(mem_22__24_), .A2(n2873), .ZN(n5857) );
  OAI21_X2 U3108 ( .B1(mem_7__24_), .B2(n2863), .A(n2859), .ZN(n5841) );
  NOR2_X1 U3109 ( .A1(mem_5__24_), .A2(n2869), .ZN(n5840) );
  NOR2_X1 U3110 ( .A1(mem_6__24_), .A2(n2873), .ZN(n5839) );
  NOR3_X2 U3111 ( .A1(n5838), .A2(n5837), .A3(n5836), .ZN(n5843) );
  NOR2_X2 U3112 ( .A1(mem_4__24_), .A2(n2853), .ZN(n5837) );
  NOR3_X2 U3113 ( .A1(n3088), .A2(n3066), .A3(mem_2__24_), .ZN(n5838) );
  NOR2_X2 U3114 ( .A1(mem_3__24_), .A2(n2856), .ZN(n5836) );
  NOR2_X2 U3115 ( .A1(mem_13__24_), .A2(n2869), .ZN(n5848) );
  NOR2_X2 U3116 ( .A1(mem_13__25_), .A2(n2870), .ZN(n5888) );
  NOR2_X2 U3117 ( .A1(mem_3__25_), .A2(n2856), .ZN(n5876) );
  NOR2_X2 U3118 ( .A1(mem_4__25_), .A2(n2853), .ZN(n5877) );
  NOR3_X2 U3119 ( .A1(n5881), .A2(n5880), .A3(n5879), .ZN(n5882) );
  OAI21_X2 U3120 ( .B1(mem_7__25_), .B2(n2862), .A(n2859), .ZN(n5881) );
  NOR2_X1 U3121 ( .A1(mem_5__25_), .A2(n2870), .ZN(n5880) );
  NOR2_X1 U3122 ( .A1(mem_6__25_), .A2(n2873), .ZN(n5879) );
  NOR2_X2 U3123 ( .A1(mem_29__25_), .A2(n2870), .ZN(n5906) );
  NOR2_X2 U3124 ( .A1(mem_30__25_), .A2(n2873), .ZN(n5905) );
  NOR3_X2 U3125 ( .A1(n5904), .A2(n5903), .A3(n5902), .ZN(n5909) );
  NOR2_X2 U3126 ( .A1(mem_28__25_), .A2(n2853), .ZN(n5903) );
  NOR2_X2 U3127 ( .A1(mem_27__25_), .A2(n2856), .ZN(n5902) );
  NOR2_X2 U3128 ( .A1(mem_21__25_), .A2(n2870), .ZN(n5898) );
  NOR2_X1 U3129 ( .A1(mem_22__25_), .A2(n2873), .ZN(n5897) );
  NOR3_X2 U3130 ( .A1(n5896), .A2(n5895), .A3(n5894), .ZN(n5901) );
  NOR2_X2 U3131 ( .A1(mem_20__25_), .A2(n2852), .ZN(n5895) );
  NOR2_X1 U3132 ( .A1(mem_13__26_), .A2(n2870), .ZN(n5928) );
  NOR2_X1 U3133 ( .A1(mem_6__26_), .A2(n2873), .ZN(n5919) );
  NOR2_X1 U3134 ( .A1(mem_5__26_), .A2(n2870), .ZN(n5920) );
  OAI21_X2 U3135 ( .B1(mem_7__26_), .B2(n2862), .A(n2860), .ZN(n5921) );
  NOR2_X2 U3136 ( .A1(mem_3__26_), .A2(n2857), .ZN(n5916) );
  NOR2_X2 U3137 ( .A1(mem_4__26_), .A2(n2852), .ZN(n5917) );
  NOR2_X2 U3138 ( .A1(mem_27__26_), .A2(n2857), .ZN(n5942) );
  NOR2_X2 U3139 ( .A1(mem_21__26_), .A2(n2870), .ZN(n5938) );
  NOR3_X2 U3140 ( .A1(n5936), .A2(n5935), .A3(n5934), .ZN(n5941) );
  NOR2_X2 U3141 ( .A1(mem_20__26_), .A2(n2853), .ZN(n5935) );
  NOR2_X2 U3142 ( .A1(mem_29__26_), .A2(n2870), .ZN(n5946) );
  NOR2_X2 U3143 ( .A1(mem_27__27_), .A2(n2857), .ZN(n5982) );
  NOR2_X2 U3144 ( .A1(mem_28__27_), .A2(n2852), .ZN(n5983) );
  NOR3_X2 U3145 ( .A1(n3086), .A2(n3066), .A3(mem_26__27_), .ZN(n5984) );
  NOR2_X2 U3146 ( .A1(mem_30__27_), .A2(n2874), .ZN(n5985) );
  NOR2_X2 U3147 ( .A1(mem_29__27_), .A2(n2870), .ZN(n5986) );
  NOR2_X2 U3148 ( .A1(mem_20__27_), .A2(n2853), .ZN(n5975) );
  NOR2_X2 U3149 ( .A1(mem_22__27_), .A2(n2874), .ZN(n5977) );
  NOR2_X2 U3150 ( .A1(mem_21__27_), .A2(n2870), .ZN(n5978) );
  OAI21_X2 U3151 ( .B1(mem_7__27_), .B2(n2862), .A(n2860), .ZN(n5961) );
  NOR2_X2 U3152 ( .A1(mem_6__27_), .A2(n2874), .ZN(n5959) );
  NOR2_X2 U3153 ( .A1(mem_5__27_), .A2(n2870), .ZN(n5960) );
  NOR3_X2 U3154 ( .A1(n5958), .A2(n5957), .A3(n5956), .ZN(n5963) );
  NOR2_X2 U3155 ( .A1(mem_4__27_), .A2(n2852), .ZN(n5957) );
  NOR2_X2 U3156 ( .A1(mem_3__27_), .A2(n2857), .ZN(n5956) );
  NOR2_X2 U3157 ( .A1(mem_13__27_), .A2(n2870), .ZN(n5968) );
  NOR3_X2 U3158 ( .A1(n5966), .A2(n5965), .A3(n5964), .ZN(n5971) );
  NOR2_X1 U3159 ( .A1(mem_13__28_), .A2(n2871), .ZN(n6008) );
  NOR3_X2 U3160 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(n6011) );
  NOR2_X1 U3161 ( .A1(mem_6__28_), .A2(n2873), .ZN(n5999) );
  NOR2_X2 U3162 ( .A1(mem_5__28_), .A2(n2870), .ZN(n6000) );
  OAI21_X2 U3163 ( .B1(mem_7__28_), .B2(n2862), .A(n2860), .ZN(n6001) );
  NOR2_X2 U3164 ( .A1(mem_3__28_), .A2(n2857), .ZN(n5996) );
  NOR2_X2 U3165 ( .A1(mem_4__28_), .A2(n2852), .ZN(n5997) );
  NOR3_X2 U3166 ( .A1(n3087), .A2(n3066), .A3(mem_2__28_), .ZN(n5998) );
  INV_X4 U3167 ( .A(n2852), .ZN(n2849) );
  NOR2_X2 U3168 ( .A1(mem_29__28_), .A2(n2871), .ZN(n6026) );
  NOR2_X2 U3169 ( .A1(mem_30__28_), .A2(n2873), .ZN(n6025) );
  NOR3_X2 U3170 ( .A1(n6024), .A2(n6023), .A3(n6022), .ZN(n6029) );
  NOR3_X2 U3171 ( .A1(n3086), .A2(n3066), .A3(mem_26__28_), .ZN(n6024) );
  NOR2_X2 U3172 ( .A1(mem_28__28_), .A2(n2854), .ZN(n6023) );
  NOR2_X2 U3173 ( .A1(mem_27__28_), .A2(n2857), .ZN(n6022) );
  NOR2_X1 U3174 ( .A1(mem_21__28_), .A2(n2871), .ZN(n6018) );
  NOR2_X1 U3175 ( .A1(mem_22__28_), .A2(n2873), .ZN(n6017) );
  NOR3_X2 U3176 ( .A1(n6016), .A2(n6015), .A3(n6014), .ZN(n6021) );
  NOR3_X2 U3177 ( .A1(n3087), .A2(n3066), .A3(mem_18__28_), .ZN(n6016) );
  NOR2_X2 U3178 ( .A1(mem_20__28_), .A2(n2854), .ZN(n6015) );
  NOR2_X2 U3179 ( .A1(mem_27__29_), .A2(n2857), .ZN(n6062) );
  NOR2_X2 U3180 ( .A1(mem_28__29_), .A2(n2854), .ZN(n6063) );
  NOR3_X2 U3181 ( .A1(n3086), .A2(n3066), .A3(mem_26__29_), .ZN(n6064) );
  OAI21_X2 U3182 ( .B1(mem_31__29_), .B2(n2863), .A(n2858), .ZN(n6067) );
  NOR2_X2 U3183 ( .A1(mem_29__29_), .A2(n2871), .ZN(n6066) );
  NOR2_X2 U3184 ( .A1(mem_30__29_), .A2(n2874), .ZN(n6065) );
  NOR2_X2 U3185 ( .A1(mem_22__29_), .A2(n2874), .ZN(n6057) );
  NOR2_X1 U3186 ( .A1(mem_21__29_), .A2(n2871), .ZN(n6058) );
  NOR2_X2 U3187 ( .A1(mem_20__29_), .A2(n2854), .ZN(n6055) );
  NOR3_X2 U3188 ( .A1(n3086), .A2(n3066), .A3(mem_18__29_), .ZN(n6056) );
  NOR3_X2 U3189 ( .A1(n6038), .A2(n6037), .A3(n6036), .ZN(n6043) );
  NOR2_X2 U3190 ( .A1(mem_4__29_), .A2(n2854), .ZN(n6037) );
  NOR2_X2 U3191 ( .A1(mem_3__29_), .A2(n2857), .ZN(n6036) );
  NOR3_X2 U3192 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(n6042) );
  OAI21_X2 U3193 ( .B1(mem_7__29_), .B2(n2863), .A(n2858), .ZN(n6041) );
  NOR2_X1 U3194 ( .A1(mem_5__29_), .A2(n2871), .ZN(n6040) );
  NOR2_X2 U3195 ( .A1(mem_6__29_), .A2(n2874), .ZN(n6039) );
  NOR3_X2 U3196 ( .A1(n6046), .A2(n6045), .A3(n6044), .ZN(n6051) );
  NOR2_X2 U3197 ( .A1(mem_13__29_), .A2(n2871), .ZN(n6048) );
  NOR2_X2 U3198 ( .A1(mem_27__30_), .A2(n2856), .ZN(n6102) );
  NOR2_X2 U3199 ( .A1(mem_28__30_), .A2(n2854), .ZN(n6103) );
  NOR3_X2 U3200 ( .A1(n3086), .A2(n3066), .A3(mem_26__30_), .ZN(n6104) );
  OAI21_X2 U3201 ( .B1(mem_31__30_), .B2(n2863), .A(n2858), .ZN(n6107) );
  NOR2_X2 U3202 ( .A1(mem_29__30_), .A2(n2871), .ZN(n6106) );
  NOR2_X2 U3203 ( .A1(mem_30__30_), .A2(n2874), .ZN(n6105) );
  NOR2_X2 U3204 ( .A1(mem_22__30_), .A2(n2874), .ZN(n6097) );
  NOR2_X1 U3205 ( .A1(mem_21__30_), .A2(n2871), .ZN(n6098) );
  NOR2_X2 U3206 ( .A1(mem_20__30_), .A2(n2854), .ZN(n6095) );
  NOR3_X2 U3207 ( .A1(n6081), .A2(n6080), .A3(n6079), .ZN(n6082) );
  OAI21_X2 U3208 ( .B1(mem_7__30_), .B2(n2863), .A(n2858), .ZN(n6081) );
  NOR2_X1 U3209 ( .A1(mem_5__30_), .A2(n2869), .ZN(n6080) );
  NOR2_X2 U3210 ( .A1(mem_6__30_), .A2(n2874), .ZN(n6079) );
  NOR3_X2 U3211 ( .A1(n6078), .A2(n6077), .A3(n6076), .ZN(n6083) );
  NOR2_X2 U3212 ( .A1(mem_4__30_), .A2(n2854), .ZN(n6077) );
  NOR3_X2 U3213 ( .A1(n3086), .A2(n3066), .A3(mem_2__30_), .ZN(n6078) );
  NOR2_X2 U3214 ( .A1(mem_3__30_), .A2(n2856), .ZN(n6076) );
  NOR3_X2 U3215 ( .A1(n6086), .A2(n6085), .A3(n6084), .ZN(n6091) );
  NOR2_X2 U3216 ( .A1(mem_13__30_), .A2(n2871), .ZN(n6088) );
  NOR2_X2 U3217 ( .A1(mem_27__31_), .A2(n2857), .ZN(n6142) );
  NOR2_X2 U3218 ( .A1(mem_28__31_), .A2(n2854), .ZN(n6143) );
  INV_X4 U3219 ( .A(n2852), .ZN(n2851) );
  OAI21_X2 U3220 ( .B1(mem_31__31_), .B2(n2863), .A(n2858), .ZN(n6149) );
  NOR2_X2 U3221 ( .A1(mem_30__31_), .A2(n2874), .ZN(n6147) );
  NOR2_X2 U3222 ( .A1(mem_20__31_), .A2(n2854), .ZN(n6135) );
  INV_X16 U3223 ( .A(n2870), .ZN(n2868) );
  NOR2_X2 U3224 ( .A1(mem_21__31_), .A2(n2871), .ZN(n6138) );
  NOR2_X2 U3225 ( .A1(mem_22__31_), .A2(n2874), .ZN(n6137) );
  INV_X4 U3226 ( .A(n2852), .ZN(n2850) );
  NOR3_X2 U3227 ( .A1(n6121), .A2(n6120), .A3(n6119), .ZN(n6122) );
  OAI21_X2 U3228 ( .B1(mem_7__31_), .B2(n2863), .A(n2858), .ZN(n6121) );
  NOR2_X1 U3229 ( .A1(mem_5__31_), .A2(n2871), .ZN(n6120) );
  NOR2_X2 U3230 ( .A1(mem_6__31_), .A2(n2874), .ZN(n6119) );
  NOR3_X2 U3231 ( .A1(n6118), .A2(n6117), .A3(n6116), .ZN(n6123) );
  NOR2_X2 U3232 ( .A1(mem_4__31_), .A2(n2854), .ZN(n6117) );
  NOR3_X1 U3233 ( .A1(n3086), .A2(n3067), .A3(mem_2__31_), .ZN(n6118) );
  NOR2_X2 U3234 ( .A1(mem_3__31_), .A2(n2857), .ZN(n6116) );
  NOR3_X2 U3235 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(n6131) );
  NOR2_X2 U3236 ( .A1(mem_13__31_), .A2(n2871), .ZN(n6128) );
  NAND3_X2 U3237 ( .A1(n2249), .A2(mem_8__26_), .A3(n3144), .ZN(n4322) );
  NAND3_X2 U3238 ( .A1(n2770), .A2(mem_9__26_), .A3(n3144), .ZN(n4321) );
  NAND3_X2 U3239 ( .A1(n2252), .A2(mem_16__27_), .A3(n3145), .ZN(n4401) );
  NAND3_X2 U3240 ( .A1(n2771), .A2(mem_17__27_), .A3(n3145), .ZN(n4400) );
  NAND3_X2 U3241 ( .A1(n2250), .A2(mem_8__24_), .A3(n3143), .ZN(n4196) );
  NAND3_X2 U3242 ( .A1(n2771), .A2(mem_9__24_), .A3(n3143), .ZN(n4195) );
  NOR3_X2 U3243 ( .A1(n3212), .A2(n3211), .A3(n3210), .ZN(n3216) );
  NOR3_X2 U3244 ( .A1(n3159), .A2(mem_18__1_), .A3(n3125), .ZN(n3211) );
  NOR2_X2 U3245 ( .A1(mem_21__1_), .A2(n2774), .ZN(n3210) );
  NOR3_X2 U3246 ( .A1(n3222), .A2(mem_23__1_), .A3(n3153), .ZN(n3214) );
  NOR3_X2 U3247 ( .A1(n3223), .A2(mem_22__1_), .A3(n3153), .ZN(n3213) );
  NOR2_X2 U3248 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  NOR2_X2 U3249 ( .A1(wData[1]), .A2(n2356), .ZN(n3251) );
  NOR2_X2 U3250 ( .A1(n2623), .A2(n3233), .ZN(n3234) );
  OAI21_X2 U3251 ( .B1(n3232), .B2(n3231), .A(n3230), .ZN(n3233) );
  NOR2_X2 U3252 ( .A1(n2622), .A2(n2499), .ZN(n3249) );
  NAND3_X2 U3253 ( .A1(n3246), .A2(n3245), .A3(n3244), .ZN(n3247) );
  AOI211_X2 U3254 ( .C1(n3227), .C2(n3226), .A(n2557), .B(n2436), .ZN(n3228)
         );
  NOR2_X2 U3255 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  NOR2_X2 U3256 ( .A1(n3673), .A2(n3672), .ZN(n3675) );
  OAI21_X2 U3257 ( .B1(wData[12]), .B2(n2355), .A(n4076), .ZN(n3674) );
  NOR2_X2 U3258 ( .A1(n3669), .A2(n3668), .ZN(n3677) );
  NOR2_X2 U3259 ( .A1(n3663), .A2(n3662), .ZN(n3669) );
  NOR2_X2 U3260 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  NOR2_X2 U3261 ( .A1(n4098), .A2(n2351), .ZN(n3695) );
  NOR2_X2 U3262 ( .A1(n4094), .A2(n2351), .ZN(n3697) );
  NOR2_X2 U3263 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  NOR2_X2 U3264 ( .A1(n4075), .A2(n4074), .ZN(n4078) );
  OAI21_X2 U3265 ( .B1(wData[22]), .B2(n2356), .A(n4076), .ZN(n4077) );
  NOR2_X2 U3266 ( .A1(n4071), .A2(n4070), .ZN(n4080) );
  NOR2_X2 U3267 ( .A1(n4065), .A2(n4064), .ZN(n4071) );
  NOR2_X2 U3268 ( .A1(n4069), .A2(n4068), .ZN(n4070) );
  NOR2_X2 U3269 ( .A1(n4098), .A2(n2349), .ZN(n4102) );
  NOR2_X2 U3270 ( .A1(n4094), .A2(n2350), .ZN(n4104) );
  INV_X4 U3271 ( .A(n2843), .ZN(n2346) );
  NOR2_X2 U3272 ( .A1(n5166), .A2(n5746), .ZN(n5167) );
  NOR2_X2 U3273 ( .A1(n5162), .A2(n2859), .ZN(n5163) );
  NAND3_X1 U3274 ( .A1(mem_1__10_), .A2(n2866), .A3(n3072), .ZN(n5205) );
  NAND3_X2 U3275 ( .A1(mem_0__10_), .A2(n2848), .A3(n3073), .ZN(n5207) );
  NOR2_X2 U3276 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  INV_X4 U3277 ( .A(n2843), .ZN(n2344) );
  NOR2_X2 U3278 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  NOR2_X2 U3279 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  NAND3_X2 U3280 ( .A1(mem_0__22_), .A2(n3106), .A3(n3084), .ZN(n5781) );
  INV_X4 U3281 ( .A(n2831), .ZN(n2830) );
  INV_X4 U3282 ( .A(n3107), .ZN(n3104) );
  INV_X4 U3283 ( .A(n4656), .ZN(n2788) );
  INV_X4 U3284 ( .A(n2764), .ZN(n2760) );
  NOR2_X2 U3285 ( .A1(mem_7__23_), .A2(n2804), .ZN(n4110) );
  NOR2_X2 U3286 ( .A1(mem_6__23_), .A2(n2795), .ZN(n4108) );
  NOR2_X2 U3287 ( .A1(mem_11__26_), .A2(n2836), .ZN(n4316) );
  NOR2_X2 U3288 ( .A1(mem_7__26_), .A2(n2803), .ZN(n4299) );
  NOR2_X2 U3289 ( .A1(mem_6__26_), .A2(n2796), .ZN(n4297) );
  NOR2_X2 U3290 ( .A1(n2657), .A2(n2796), .ZN(n4327) );
  NOR2_X2 U3291 ( .A1(n2659), .A2(n2803), .ZN(n4406) );
  NOR2_X2 U3292 ( .A1(n2649), .A2(n2781), .ZN(n4405) );
  NOR2_X2 U3293 ( .A1(mem_7__27_), .A2(n2803), .ZN(n4362) );
  NOR2_X2 U3294 ( .A1(mem_6__27_), .A2(n2797), .ZN(n4360) );
  NOR2_X2 U3295 ( .A1(mem_2__24_), .A2(n3132), .ZN(n4178) );
  NOR2_X2 U3296 ( .A1(mem_3__24_), .A2(n2836), .ZN(n4176) );
  NOR2_X2 U3297 ( .A1(n2661), .A2(n2804), .ZN(n4217) );
  NOR2_X2 U3298 ( .A1(n2651), .A2(n2780), .ZN(n4216) );
  NOR2_X2 U3299 ( .A1(rd[2]), .A2(rd[3]), .ZN(n746) );
  NOR2_X2 U3300 ( .A1(n7229), .A2(rd[3]), .ZN(n241) );
  NOR2_X2 U3301 ( .A1(n7228), .A2(rd[2]), .ZN(n578) );
  NOR2_X2 U3302 ( .A1(n7229), .A2(n7228), .ZN(n444) );
  INV_X4 U3303 ( .A(rs2[2]), .ZN(n3135) );
  NOR2_X2 U3304 ( .A1(mem_27__1_), .A2(n3163), .ZN(n3217) );
  INV_X16 U3305 ( .A(n2799), .ZN(n2796) );
  NOR2_X2 U3306 ( .A1(mem_7__25_), .A2(n2804), .ZN(n4236) );
  NOR2_X2 U3307 ( .A1(mem_6__25_), .A2(n2796), .ZN(n4234) );
  NOR2_X2 U3308 ( .A1(mem_21__25_), .A2(n2780), .ZN(n4265) );
  INV_X16 U3309 ( .A(n2812), .ZN(n2804) );
  NOR2_X2 U3310 ( .A1(mem_2__28_), .A2(n3133), .ZN(n4430) );
  NOR2_X2 U3311 ( .A1(mem_3__28_), .A2(n2837), .ZN(n4428) );
  NOR2_X2 U3312 ( .A1(n2719), .A2(n2797), .ZN(n4467) );
  NOR2_X2 U3313 ( .A1(mem_7__29_), .A2(n2806), .ZN(n4488) );
  NOR2_X2 U3314 ( .A1(mem_6__29_), .A2(n2797), .ZN(n4486) );
  NOR2_X2 U3315 ( .A1(n2709), .A2(n2797), .ZN(n4530) );
  NOR2_X2 U3316 ( .A1(n2713), .A2(n2798), .ZN(n4658) );
  NOR2_X2 U3317 ( .A1(n2681), .A2(n2782), .ZN(n4659) );
  INV_X4 U3318 ( .A(n2847), .ZN(n2846) );
  INV_X16 U3319 ( .A(rs1[2]), .ZN(n3068) );
  INV_X4 U3320 ( .A(n5749), .ZN(n5798) );
  NOR2_X2 U3321 ( .A1(n3063), .A2(n3076), .ZN(n5765) );
  INV_X4 U3322 ( .A(n2858), .ZN(n2861) );
  NOR2_X2 U3323 ( .A1(n4139), .A2(n4138), .ZN(n4142) );
  NOR2_X2 U3324 ( .A1(mem_21__23_), .A2(n2779), .ZN(n4139) );
  NOR2_X2 U3325 ( .A1(mem_22__23_), .A2(n2795), .ZN(n4138) );
  NOR2_X2 U3326 ( .A1(n2762), .A2(n4140), .ZN(n4141) );
  NOR2_X2 U3327 ( .A1(n4144), .A2(n4143), .ZN(n4147) );
  NOR2_X2 U3328 ( .A1(mem_19__23_), .A2(n2835), .ZN(n4143) );
  NOR2_X2 U3329 ( .A1(n4123), .A2(n4122), .ZN(n4126) );
  NOR2_X2 U3330 ( .A1(mem_14__23_), .A2(n2795), .ZN(n4122) );
  NOR2_X2 U3331 ( .A1(mem_13__23_), .A2(n2779), .ZN(n4123) );
  NOR2_X2 U3332 ( .A1(n4128), .A2(n4127), .ZN(n4131) );
  NOR2_X2 U3333 ( .A1(mem_12__23_), .A2(n2319), .ZN(n4128) );
  NOR2_X2 U3334 ( .A1(n4391), .A2(n4390), .ZN(n4394) );
  NOR2_X2 U3335 ( .A1(mem_21__27_), .A2(n2781), .ZN(n4391) );
  NOR2_X2 U3336 ( .A1(mem_22__27_), .A2(n2797), .ZN(n4390) );
  NAND2_X2 U3337 ( .A1(n4381), .A2(n3161), .ZN(n4382) );
  NOR2_X2 U3338 ( .A1(n4380), .A2(n4379), .ZN(n4383) );
  NOR2_X2 U3339 ( .A1(mem_12__27_), .A2(n2319), .ZN(n4380) );
  NOR2_X2 U3340 ( .A1(mem_11__27_), .A2(n2837), .ZN(n4379) );
  NOR2_X2 U3341 ( .A1(n4375), .A2(n4374), .ZN(n4378) );
  NOR2_X2 U3342 ( .A1(mem_14__27_), .A2(n2797), .ZN(n4374) );
  NOR2_X2 U3343 ( .A1(n4202), .A2(n4201), .ZN(n4205) );
  NOR2_X2 U3344 ( .A1(mem_21__24_), .A2(n2780), .ZN(n4202) );
  NOR2_X2 U3345 ( .A1(mem_22__24_), .A2(n2796), .ZN(n4201) );
  NOR2_X2 U3346 ( .A1(n2762), .A2(n4203), .ZN(n4204) );
  NOR2_X2 U3347 ( .A1(n4207), .A2(n4206), .ZN(n4210) );
  NOR2_X2 U3348 ( .A1(mem_19__24_), .A2(n2836), .ZN(n4206) );
  NOR2_X2 U3349 ( .A1(mem_19__1_), .A2(n3163), .ZN(n3208) );
  OAI21_X2 U3350 ( .B1(mem_3__1_), .B2(n3163), .A(rs2[1]), .ZN(n3231) );
  NOR2_X2 U3351 ( .A1(mem_2__1_), .A2(n3159), .ZN(n3232) );
  NAND3_X2 U3352 ( .A1(mem_0__1_), .A2(n3162), .A3(n3155), .ZN(n3230) );
  NOR2_X2 U3353 ( .A1(mem_14__1_), .A2(n3155), .ZN(n3242) );
  NOR2_X2 U3354 ( .A1(mem_10__1_), .A2(n3159), .ZN(n3238) );
  NAND3_X2 U3355 ( .A1(mem_8__1_), .A2(n3162), .A3(n3154), .ZN(n3236) );
  OAI21_X2 U3356 ( .B1(mem_11__1_), .B2(n3163), .A(rs2[1]), .ZN(n3237) );
  NOR2_X2 U3357 ( .A1(n3241), .A2(n3240), .ZN(n3246) );
  NOR3_X2 U3358 ( .A1(rs2[1]), .A2(mem_13__1_), .A3(n3162), .ZN(n3240) );
  NOR3_X2 U3359 ( .A1(rs2[1]), .A2(mem_12__1_), .A3(n3156), .ZN(n3241) );
  AOI21_X2 U3360 ( .B1(n3243), .B2(n3159), .A(n3153), .ZN(n3244) );
  NOR2_X2 U3361 ( .A1(mem_15__1_), .A2(n3155), .ZN(n3243) );
  NOR3_X2 U3362 ( .A1(n3223), .A2(mem_30__1_), .A3(n3153), .ZN(n3224) );
  NOR3_X2 U3363 ( .A1(n3222), .A2(mem_31__1_), .A3(n3153), .ZN(n3225) );
  NOR2_X2 U3364 ( .A1(n4270), .A2(n4269), .ZN(n4273) );
  NOR2_X2 U3365 ( .A1(mem_19__25_), .A2(n2836), .ZN(n4269) );
  NOR2_X2 U3366 ( .A1(n2647), .A2(n3132), .ZN(n4271) );
  NOR2_X2 U3367 ( .A1(n2643), .A2(n3133), .ZN(n4460) );
  NOR2_X2 U3368 ( .A1(n2762), .A2(n4455), .ZN(n4456) );
  NOR2_X2 U3369 ( .A1(n4454), .A2(n4453), .ZN(n4457) );
  NOR2_X2 U3370 ( .A1(n2641), .A2(n3133), .ZN(n4523) );
  NOR2_X2 U3371 ( .A1(n4517), .A2(n4516), .ZN(n4520) );
  NOR2_X2 U3372 ( .A1(mem_21__29_), .A2(n2781), .ZN(n4517) );
  NOR2_X2 U3373 ( .A1(n4569), .A2(n4568), .ZN(n4572) );
  NOR2_X2 U3374 ( .A1(mem_12__30_), .A2(n2320), .ZN(n4569) );
  NOR2_X2 U3375 ( .A1(mem_11__30_), .A2(n2838), .ZN(n4568) );
  NOR2_X2 U3376 ( .A1(n4564), .A2(n4563), .ZN(n4567) );
  NOR2_X2 U3377 ( .A1(mem_14__30_), .A2(n2798), .ZN(n4563) );
  NOR2_X2 U3378 ( .A1(mem_2__30_), .A2(n3133), .ZN(n4556) );
  NOR2_X2 U3379 ( .A1(n4555), .A2(n4554), .ZN(n4558) );
  NOR2_X2 U3380 ( .A1(mem_4__30_), .A2(n2320), .ZN(n4555) );
  NOR2_X2 U3381 ( .A1(mem_3__30_), .A2(n2838), .ZN(n4554) );
  NOR2_X2 U3382 ( .A1(n4550), .A2(n4549), .ZN(n4553) );
  NOR2_X2 U3383 ( .A1(mem_5__30_), .A2(n2781), .ZN(n4550) );
  NOR2_X2 U3384 ( .A1(n4585), .A2(n4584), .ZN(n4588) );
  NOR2_X2 U3385 ( .A1(mem_19__30_), .A2(n2838), .ZN(n4584) );
  NOR2_X2 U3386 ( .A1(n4580), .A2(n4579), .ZN(n4583) );
  NOR2_X2 U3387 ( .A1(mem_21__30_), .A2(n2781), .ZN(n4580) );
  NOR2_X2 U3388 ( .A1(n4594), .A2(n4593), .ZN(n4597) );
  NOR2_X2 U3389 ( .A1(n2683), .A2(n2782), .ZN(n4594) );
  NOR2_X2 U3390 ( .A1(n2711), .A2(n2798), .ZN(n4593) );
  NOR2_X2 U3391 ( .A1(n2745), .A2(n2801), .ZN(n4595) );
  NOR2_X2 U3392 ( .A1(n4599), .A2(n4598), .ZN(n4602) );
  NOR2_X2 U3393 ( .A1(n2727), .A2(n2838), .ZN(n4598) );
  NOR2_X2 U3394 ( .A1(n2699), .A2(n2318), .ZN(n4599) );
  NOR2_X2 U3395 ( .A1(n2749), .A2(n3134), .ZN(n4600) );
  NOR2_X2 U3396 ( .A1(n6163), .A2(n6164), .ZN(n3205) );
  AOI21_X2 U3397 ( .B1(n4684), .B2(n2365), .A(n3204), .ZN(n3206) );
  NOR2_X2 U3398 ( .A1(mem_2__31_), .A2(n3134), .ZN(n4619) );
  NOR2_X2 U3399 ( .A1(n4618), .A2(n4617), .ZN(n4621) );
  NOR2_X2 U3400 ( .A1(mem_4__31_), .A2(n2321), .ZN(n4618) );
  NOR2_X2 U3401 ( .A1(mem_3__31_), .A2(n2838), .ZN(n4617) );
  NOR2_X2 U3402 ( .A1(n4613), .A2(n4612), .ZN(n4616) );
  NOR2_X2 U3403 ( .A1(mem_5__31_), .A2(n2782), .ZN(n4613) );
  NOR2_X2 U3404 ( .A1(n4643), .A2(n4642), .ZN(n4646) );
  NOR2_X2 U3405 ( .A1(mem_21__31_), .A2(n2782), .ZN(n4643) );
  INV_X4 U3406 ( .A(n3108), .ZN(n3097) );
  INV_X4 U3407 ( .A(n3108), .ZN(n3096) );
  INV_X4 U3408 ( .A(n3108), .ZN(n3095) );
  INV_X16 U3409 ( .A(n3110), .ZN(n3103) );
  AOI21_X2 U3410 ( .B1(n5196), .B2(n3106), .A(n5195), .ZN(n5203) );
  NOR2_X2 U3411 ( .A1(mem_5__10_), .A2(n2869), .ZN(n5195) );
  NOR2_X2 U3412 ( .A1(n3067), .A2(mem_2__10_), .ZN(n5196) );
  AOI21_X2 U3413 ( .B1(n5198), .B2(n5197), .A(n2861), .ZN(n5202) );
  NOR2_X2 U3414 ( .A1(n3088), .A2(n3084), .ZN(n5197) );
  NOR2_X2 U3415 ( .A1(mem_6__10_), .A2(n3071), .ZN(n5198) );
  NOR2_X2 U3416 ( .A1(n3108), .A2(n3084), .ZN(n5199) );
  NOR2_X2 U3417 ( .A1(mem_7__10_), .A2(n3072), .ZN(n5200) );
  AOI21_X2 U3418 ( .B1(n5194), .B2(n3070), .A(n5193), .ZN(n5204) );
  NOR2_X2 U3419 ( .A1(mem_3__10_), .A2(n3105), .ZN(n5194) );
  NOR2_X2 U3420 ( .A1(mem_4__10_), .A2(n2853), .ZN(n5193) );
  NOR3_X2 U3421 ( .A1(n3059), .A2(n5186), .A3(n5743), .ZN(n5187) );
  NOR3_X2 U3422 ( .A1(n3063), .A2(n5185), .A3(n5746), .ZN(n5188) );
  NOR2_X2 U3423 ( .A1(n5183), .A2(n2859), .ZN(n5184) );
  INV_X4 U3424 ( .A(n3105), .ZN(n3091) );
  INV_X4 U3425 ( .A(n3105), .ZN(n3090) );
  INV_X4 U3426 ( .A(n3105), .ZN(n3089) );
  INV_X4 U3427 ( .A(n3106), .ZN(n3092) );
  INV_X4 U3428 ( .A(n3106), .ZN(n3093) );
  INV_X4 U3429 ( .A(n3106), .ZN(n3094) );
  OAI21_X2 U3430 ( .B1(mem_7__22_), .B2(n3106), .A(n3074), .ZN(n5786) );
  NAND3_X2 U3431 ( .A1(mem_4__22_), .A2(n3105), .A3(n3084), .ZN(n5785) );
  NOR2_X2 U3432 ( .A1(n3088), .A2(mem_6__22_), .ZN(n5787) );
  NAND3_X2 U3433 ( .A1(mem_5__22_), .A2(n3086), .A3(n3084), .ZN(n5784) );
  OAI21_X2 U3434 ( .B1(mem_3__22_), .B2(n3108), .A(n3075), .ZN(n5782) );
  NOR2_X2 U3435 ( .A1(n3088), .A2(mem_2__22_), .ZN(n5783) );
  NAND3_X2 U3436 ( .A1(mem_1__22_), .A2(n3086), .A3(n3084), .ZN(n5780) );
  NOR2_X2 U3437 ( .A1(n5774), .A2(n2859), .ZN(n5775) );
  NAND3_X2 U3438 ( .A1(mem_8__22_), .A2(n3108), .A3(n3084), .ZN(n5771) );
  NAND3_X2 U3439 ( .A1(mem_9__22_), .A2(n3086), .A3(n3084), .ZN(n5772) );
  NAND3_X2 U3440 ( .A1(n2258), .A2(mem_24__23_), .A3(n3142), .ZN(n4163) );
  NAND3_X2 U3441 ( .A1(n2771), .A2(mem_25__23_), .A3(n3143), .ZN(n4162) );
  NAND3_X2 U3442 ( .A1(n2301), .A2(mem_0__23_), .A3(n3142), .ZN(n4119) );
  NAND3_X2 U3443 ( .A1(n2302), .A2(mem_0__26_), .A3(n3144), .ZN(n4308) );
  NAND3_X2 U3444 ( .A1(n2255), .A2(mem_24__26_), .A3(n3145), .ZN(n4352) );
  NAND3_X2 U3445 ( .A1(n2772), .A2(mem_25__26_), .A3(n3145), .ZN(n4351) );
  NAND2_X2 U3446 ( .A1(n4336), .A2(n4335), .ZN(n4339) );
  NAND3_X2 U3447 ( .A1(n2259), .A2(mem_16__26_), .A3(n3144), .ZN(n4338) );
  NAND3_X2 U3448 ( .A1(n2784), .A2(mem_17__26_), .A3(n3144), .ZN(n4337) );
  NAND3_X2 U3449 ( .A1(n2276), .A2(mem_24__27_), .A3(n3145), .ZN(n4415) );
  NAND3_X2 U3450 ( .A1(n2772), .A2(mem_25__27_), .A3(n3145), .ZN(n4414) );
  NAND3_X2 U3451 ( .A1(n2304), .A2(mem_0__27_), .A3(n3145), .ZN(n4371) );
  NAND3_X2 U3452 ( .A1(n2771), .A2(mem_1__27_), .A3(n3145), .ZN(n4370) );
  NAND3_X2 U3453 ( .A1(n2255), .A2(mem_0__24_), .A3(n3143), .ZN(n4182) );
  NAND3_X2 U3454 ( .A1(n2772), .A2(mem_1__24_), .A3(n3143), .ZN(n4181) );
  NAND3_X2 U3455 ( .A1(n2253), .A2(mem_24__24_), .A3(n3143), .ZN(n4226) );
  NAND3_X2 U3456 ( .A1(n2770), .A2(mem_25__24_), .A3(n3143), .ZN(n4225) );
  AOI211_X2 U3457 ( .C1(n3180), .C2(n3179), .A(n2553), .B(n2432), .ZN(n3181)
         );
  NOR3_X2 U3458 ( .A1(n3175), .A2(n3174), .A3(n3173), .ZN(n3180) );
  AOI211_X2 U3459 ( .C1(n3172), .C2(n3171), .A(n2483), .B(n2604), .ZN(n3182)
         );
  NOR3_X2 U3460 ( .A1(n3167), .A2(n3166), .A3(n3165), .ZN(n3172) );
  NOR3_X2 U3461 ( .A1(n3170), .A2(n3169), .A3(n3168), .ZN(n3171) );
  AOI211_X2 U3462 ( .C1(n3190), .C2(n3189), .A(n2554), .B(n2433), .ZN(n3200)
         );
  AOI211_X2 U3463 ( .C1(n3198), .C2(n3197), .A(n2555), .B(n2434), .ZN(n3199)
         );
  AOI211_X2 U3464 ( .C1(n3275), .C2(n3274), .A(n2558), .B(n2437), .ZN(n3276)
         );
  NOR3_X2 U3465 ( .A1(n3270), .A2(n3269), .A3(n3268), .ZN(n3275) );
  AOI211_X2 U3466 ( .C1(n3267), .C2(n3266), .A(n2372), .B(n2605), .ZN(n3277)
         );
  NOR3_X2 U3467 ( .A1(n3262), .A2(n3261), .A3(n3260), .ZN(n3267) );
  NOR3_X2 U3468 ( .A1(n3265), .A2(n3264), .A3(n3263), .ZN(n3266) );
  AOI211_X2 U3469 ( .C1(n3285), .C2(n3284), .A(n2559), .B(n2438), .ZN(n3295)
         );
  AOI211_X2 U3470 ( .C1(n3293), .C2(n3292), .A(n2560), .B(n2439), .ZN(n3294)
         );
  AOI211_X2 U3471 ( .C1(n3315), .C2(n3314), .A(n2561), .B(n2440), .ZN(n3316)
         );
  NOR3_X2 U3472 ( .A1(n3310), .A2(n3309), .A3(n3308), .ZN(n3315) );
  AOI211_X2 U3473 ( .C1(n3307), .C2(n3306), .A(n2484), .B(n2606), .ZN(n3317)
         );
  NOR3_X2 U3474 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(n3307) );
  NOR3_X2 U3475 ( .A1(n3305), .A2(n3304), .A3(n3303), .ZN(n3306) );
  AOI211_X2 U3476 ( .C1(n3325), .C2(n3324), .A(n2562), .B(n2441), .ZN(n3335)
         );
  AOI211_X2 U3477 ( .C1(n3333), .C2(n3332), .A(n2563), .B(n2442), .ZN(n3334)
         );
  AOI211_X2 U3478 ( .C1(n3355), .C2(n3354), .A(n2564), .B(n2443), .ZN(n3356)
         );
  NOR3_X2 U3479 ( .A1(n3350), .A2(n3349), .A3(n3348), .ZN(n3355) );
  AOI211_X2 U3480 ( .C1(n3347), .C2(n3346), .A(n2485), .B(n2607), .ZN(n3357)
         );
  NOR3_X2 U3481 ( .A1(n3342), .A2(n3341), .A3(n3340), .ZN(n3347) );
  NOR3_X2 U3482 ( .A1(n3345), .A2(n3344), .A3(n3343), .ZN(n3346) );
  AOI211_X2 U3483 ( .C1(n3365), .C2(n3364), .A(n2565), .B(n2444), .ZN(n3375)
         );
  AOI211_X2 U3484 ( .C1(n3395), .C2(n3394), .A(n2566), .B(n2445), .ZN(n3396)
         );
  NOR3_X2 U3485 ( .A1(n3390), .A2(n3389), .A3(n3388), .ZN(n3395) );
  AOI211_X2 U3486 ( .C1(n3387), .C2(n3386), .A(n2486), .B(n2608), .ZN(n3397)
         );
  NOR3_X2 U3487 ( .A1(n3382), .A2(n3381), .A3(n3380), .ZN(n3387) );
  NOR3_X2 U3488 ( .A1(n3385), .A2(n3384), .A3(n3383), .ZN(n3386) );
  AOI211_X2 U3489 ( .C1(n3405), .C2(n3404), .A(n2567), .B(n2446), .ZN(n3415)
         );
  AOI211_X2 U3490 ( .C1(n3435), .C2(n3434), .A(n2568), .B(n2447), .ZN(n3436)
         );
  NOR3_X2 U3491 ( .A1(n3430), .A2(n3429), .A3(n3428), .ZN(n3435) );
  AOI211_X2 U3492 ( .C1(n3427), .C2(n3426), .A(n2487), .B(n2609), .ZN(n3437)
         );
  NOR3_X2 U3493 ( .A1(n3422), .A2(n3421), .A3(n3420), .ZN(n3427) );
  NOR3_X2 U3494 ( .A1(n3425), .A2(n3424), .A3(n3423), .ZN(n3426) );
  AOI211_X2 U3495 ( .C1(n3445), .C2(n3444), .A(n2569), .B(n2448), .ZN(n3455)
         );
  AOI211_X2 U3496 ( .C1(n3453), .C2(n3452), .A(n2570), .B(n2449), .ZN(n3454)
         );
  AOI211_X2 U3497 ( .C1(n3475), .C2(n3474), .A(n2571), .B(n2450), .ZN(n3476)
         );
  NOR3_X2 U3498 ( .A1(n3473), .A2(n3472), .A3(n3471), .ZN(n3474) );
  AOI211_X2 U3499 ( .C1(n3467), .C2(n3466), .A(n2488), .B(n2610), .ZN(n3477)
         );
  NOR3_X2 U3500 ( .A1(n3465), .A2(n3464), .A3(n3463), .ZN(n3466) );
  NOR3_X2 U3501 ( .A1(n3462), .A2(n3461), .A3(n3460), .ZN(n3467) );
  AOI211_X2 U3502 ( .C1(n3485), .C2(n3484), .A(n2572), .B(n2451), .ZN(n3495)
         );
  AOI211_X2 U3503 ( .C1(n3493), .C2(n3492), .A(n2573), .B(n2452), .ZN(n3494)
         );
  AOI211_X2 U3504 ( .C1(n3515), .C2(n3514), .A(n2574), .B(n2453), .ZN(n3516)
         );
  NOR3_X2 U3505 ( .A1(n3513), .A2(n3512), .A3(n3511), .ZN(n3514) );
  NOR3_X2 U3506 ( .A1(n3510), .A2(n3509), .A3(n3508), .ZN(n3515) );
  AOI211_X2 U3507 ( .C1(n3507), .C2(n3506), .A(n2489), .B(n2611), .ZN(n3517)
         );
  NOR3_X2 U3508 ( .A1(n3505), .A2(n3504), .A3(n3503), .ZN(n3506) );
  NOR3_X2 U3509 ( .A1(n3502), .A2(n3501), .A3(n3500), .ZN(n3507) );
  AOI211_X2 U3510 ( .C1(n3525), .C2(n3524), .A(n2575), .B(n2454), .ZN(n3535)
         );
  AOI211_X2 U3511 ( .C1(n3533), .C2(n3532), .A(n2576), .B(n2455), .ZN(n3534)
         );
  AOI211_X2 U3512 ( .C1(n3555), .C2(n3554), .A(n2577), .B(n2456), .ZN(n3556)
         );
  NOR3_X2 U3513 ( .A1(n3550), .A2(n3549), .A3(n3548), .ZN(n3555) );
  AOI211_X2 U3514 ( .C1(n3547), .C2(n3546), .A(n2490), .B(n2612), .ZN(n3557)
         );
  NOR3_X2 U3515 ( .A1(n3542), .A2(n3541), .A3(n3540), .ZN(n3547) );
  NOR3_X2 U3516 ( .A1(n3545), .A2(n3544), .A3(n3543), .ZN(n3546) );
  AOI211_X2 U3517 ( .C1(n3565), .C2(n3564), .A(n2578), .B(n2457), .ZN(n3575)
         );
  AOI211_X2 U3518 ( .C1(n3573), .C2(n3572), .A(n2579), .B(n2458), .ZN(n3574)
         );
  AOI211_X2 U3519 ( .C1(n3595), .C2(n3594), .A(n2580), .B(n2459), .ZN(n3596)
         );
  NOR3_X2 U3520 ( .A1(n3590), .A2(n3589), .A3(n3588), .ZN(n3595) );
  AOI211_X2 U3521 ( .C1(n3587), .C2(n3586), .A(n2498), .B(n2620), .ZN(n3597)
         );
  NOR3_X2 U3522 ( .A1(n3582), .A2(n3581), .A3(n3580), .ZN(n3587) );
  AOI211_X2 U3523 ( .C1(n3605), .C2(n3604), .A(n2581), .B(n2460), .ZN(n3615)
         );
  AOI211_X2 U3524 ( .C1(n3613), .C2(n3612), .A(n2582), .B(n2461), .ZN(n3614)
         );
  AOI211_X2 U3525 ( .C1(n3635), .C2(n3634), .A(n2583), .B(n2462), .ZN(n3636)
         );
  NOR3_X2 U3526 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n3635) );
  AOI211_X2 U3527 ( .C1(n3627), .C2(n3626), .A(n2491), .B(n2613), .ZN(n3637)
         );
  NOR3_X2 U3528 ( .A1(n3622), .A2(n3621), .A3(n3620), .ZN(n3627) );
  NOR3_X2 U3529 ( .A1(n3625), .A2(n3624), .A3(n3623), .ZN(n3626) );
  AOI211_X2 U3530 ( .C1(n3645), .C2(n3644), .A(n2584), .B(n2463), .ZN(n3655)
         );
  AOI211_X2 U3531 ( .C1(n3653), .C2(n3652), .A(n2585), .B(n2464), .ZN(n3654)
         );
  AOI211_X2 U3532 ( .C1(n3716), .C2(n3715), .A(n2586), .B(n2465), .ZN(n3717)
         );
  NOR3_X2 U3533 ( .A1(n3711), .A2(n3710), .A3(n3709), .ZN(n3716) );
  AOI211_X2 U3534 ( .C1(n3708), .C2(n3707), .A(n2492), .B(n2614), .ZN(n3718)
         );
  NOR3_X2 U3535 ( .A1(n3703), .A2(n3702), .A3(n3701), .ZN(n3708) );
  AOI211_X2 U3536 ( .C1(n3726), .C2(n3725), .A(n2587), .B(n2466), .ZN(n3736)
         );
  AOI211_X2 U3537 ( .C1(n3734), .C2(n3733), .A(n2588), .B(n2467), .ZN(n3735)
         );
  AOI211_X2 U3538 ( .C1(n3756), .C2(n3755), .A(n2589), .B(n2468), .ZN(n3757)
         );
  NOR3_X2 U3539 ( .A1(n3751), .A2(n3750), .A3(n3749), .ZN(n3756) );
  AOI211_X2 U3540 ( .C1(n3748), .C2(n3747), .A(n2493), .B(n2615), .ZN(n3758)
         );
  NOR3_X2 U3541 ( .A1(n3743), .A2(n3742), .A3(n3741), .ZN(n3748) );
  NOR3_X2 U3542 ( .A1(n3746), .A2(n3745), .A3(n3744), .ZN(n3747) );
  AOI211_X2 U3543 ( .C1(n3766), .C2(n3765), .A(n2590), .B(n2469), .ZN(n3776)
         );
  AOI211_X2 U3544 ( .C1(n3774), .C2(n3773), .A(n2591), .B(n2470), .ZN(n3775)
         );
  AOI211_X2 U3545 ( .C1(n3796), .C2(n3795), .A(n2592), .B(n2471), .ZN(n3797)
         );
  NOR3_X2 U3546 ( .A1(n3791), .A2(n3790), .A3(n3789), .ZN(n3796) );
  AOI211_X2 U3547 ( .C1(n3788), .C2(n3787), .A(n2494), .B(n2616), .ZN(n3798)
         );
  NOR3_X2 U3548 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n3788) );
  NOR3_X2 U3549 ( .A1(n3786), .A2(n3785), .A3(n3784), .ZN(n3787) );
  AOI211_X2 U3550 ( .C1(n3806), .C2(n3805), .A(n2419), .B(n2506), .ZN(n3816)
         );
  AOI211_X2 U3551 ( .C1(n3814), .C2(n3813), .A(n2420), .B(n2507), .ZN(n3815)
         );
  AOI211_X2 U3552 ( .C1(n3836), .C2(n3835), .A(n2422), .B(n2509), .ZN(n3837)
         );
  NOR3_X2 U3553 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(n3836) );
  AOI211_X2 U3554 ( .C1(n3828), .C2(n3827), .A(n2421), .B(n2508), .ZN(n3838)
         );
  NOR3_X2 U3555 ( .A1(n3823), .A2(n3822), .A3(n3821), .ZN(n3828) );
  AOI211_X2 U3556 ( .C1(n3846), .C2(n3845), .A(n2423), .B(n2510), .ZN(n3856)
         );
  AOI211_X2 U3557 ( .C1(n3854), .C2(n3853), .A(n2424), .B(n2511), .ZN(n3855)
         );
  AOI211_X2 U3558 ( .C1(n3876), .C2(n3875), .A(n2426), .B(n2513), .ZN(n3877)
         );
  NOR3_X2 U3559 ( .A1(n3871), .A2(n3870), .A3(n3869), .ZN(n3876) );
  AOI211_X2 U3560 ( .C1(n3868), .C2(n3867), .A(n2425), .B(n2512), .ZN(n3878)
         );
  NOR3_X2 U3561 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3868) );
  AOI211_X2 U3562 ( .C1(n3886), .C2(n3885), .A(n2427), .B(n2514), .ZN(n3896)
         );
  AOI211_X2 U3563 ( .C1(n3894), .C2(n3893), .A(n2428), .B(n2515), .ZN(n3895)
         );
  AOI211_X2 U3564 ( .C1(n3916), .C2(n3915), .A(n2430), .B(n2552), .ZN(n3917)
         );
  NOR3_X2 U3565 ( .A1(n3911), .A2(n3910), .A3(n3909), .ZN(n3916) );
  AOI211_X2 U3566 ( .C1(n3908), .C2(n3907), .A(n2429), .B(n2516), .ZN(n3918)
         );
  NOR3_X2 U3567 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3908) );
  AOI211_X2 U3568 ( .C1(n3926), .C2(n3925), .A(n2593), .B(n2472), .ZN(n3936)
         );
  AOI211_X2 U3569 ( .C1(n3934), .C2(n3933), .A(n2594), .B(n2473), .ZN(n3935)
         );
  AOI211_X2 U3570 ( .C1(n3956), .C2(n3955), .A(n2595), .B(n2474), .ZN(n3957)
         );
  NOR3_X2 U3571 ( .A1(n3951), .A2(n3950), .A3(n3949), .ZN(n3956) );
  AOI211_X2 U3572 ( .C1(n3948), .C2(n3947), .A(n2495), .B(n2617), .ZN(n3958)
         );
  NOR3_X2 U3573 ( .A1(n3943), .A2(n3942), .A3(n3941), .ZN(n3948) );
  NOR3_X2 U3574 ( .A1(n3946), .A2(n3945), .A3(n3944), .ZN(n3947) );
  AOI211_X2 U3575 ( .C1(n3966), .C2(n3965), .A(n2596), .B(n2475), .ZN(n3976)
         );
  AOI211_X2 U3576 ( .C1(n3974), .C2(n3973), .A(n2597), .B(n2476), .ZN(n3975)
         );
  AOI211_X2 U3577 ( .C1(n3996), .C2(n3995), .A(n2598), .B(n2477), .ZN(n3997)
         );
  NOR3_X2 U3578 ( .A1(n3991), .A2(n3990), .A3(n3989), .ZN(n3996) );
  NOR3_X2 U3579 ( .A1(n3994), .A2(n3993), .A3(n3992), .ZN(n3995) );
  AOI211_X2 U3580 ( .C1(n3988), .C2(n3987), .A(n2496), .B(n2618), .ZN(n3998)
         );
  NOR3_X2 U3581 ( .A1(n3983), .A2(n3982), .A3(n3981), .ZN(n3988) );
  NOR3_X2 U3582 ( .A1(n3986), .A2(n3985), .A3(n3984), .ZN(n3987) );
  AOI211_X2 U3583 ( .C1(n4006), .C2(n4005), .A(n2599), .B(n2478), .ZN(n4016)
         );
  AOI211_X2 U3584 ( .C1(n4014), .C2(n4013), .A(n2600), .B(n2479), .ZN(n4015)
         );
  AOI211_X2 U3585 ( .C1(n4036), .C2(n4035), .A(n2601), .B(n2480), .ZN(n4037)
         );
  NOR3_X2 U3586 ( .A1(n4031), .A2(n4030), .A3(n4029), .ZN(n4036) );
  NOR3_X2 U3587 ( .A1(n4034), .A2(n4033), .A3(n4032), .ZN(n4035) );
  AOI211_X2 U3588 ( .C1(n4028), .C2(n4027), .A(n2497), .B(n2619), .ZN(n4038)
         );
  NOR3_X2 U3589 ( .A1(n4023), .A2(n4022), .A3(n4021), .ZN(n4028) );
  NOR3_X2 U3590 ( .A1(n4026), .A2(n4025), .A3(n4024), .ZN(n4027) );
  AOI211_X2 U3591 ( .C1(n4046), .C2(n4045), .A(n2602), .B(n2481), .ZN(n4057)
         );
  AOI211_X2 U3592 ( .C1(n4055), .C2(n4054), .A(n2603), .B(n2482), .ZN(n4056)
         );
  NAND3_X2 U3593 ( .A1(n2247), .A2(mem_8__25_), .A3(n3144), .ZN(n4259) );
  NAND3_X2 U3594 ( .A1(n2770), .A2(mem_9__25_), .A3(n3144), .ZN(n4258) );
  NAND3_X2 U3595 ( .A1(n2286), .A2(mem_0__25_), .A3(n3143), .ZN(n4245) );
  NAND2_X2 U3596 ( .A1(n4287), .A2(n4286), .ZN(n4290) );
  NAND3_X2 U3597 ( .A1(n2290), .A2(mem_24__25_), .A3(n3144), .ZN(n4289) );
  NAND3_X2 U3598 ( .A1(n2244), .A2(mem_8__28_), .A3(n3146), .ZN(n4448) );
  NAND3_X2 U3599 ( .A1(n2771), .A2(mem_9__28_), .A3(n3146), .ZN(n4447) );
  NAND3_X2 U3600 ( .A1(n2288), .A2(mem_0__28_), .A3(n3145), .ZN(n4434) );
  NAND3_X2 U3601 ( .A1(n2771), .A2(mem_1__28_), .A3(n3145), .ZN(n4433) );
  NAND2_X2 U3602 ( .A1(n4476), .A2(n4475), .ZN(n4479) );
  NAND3_X2 U3603 ( .A1(n2289), .A2(mem_24__28_), .A3(n3146), .ZN(n4478) );
  NAND3_X2 U3604 ( .A1(n2771), .A2(mem_25__28_), .A3(n3146), .ZN(n4477) );
  NAND3_X2 U3605 ( .A1(n2246), .A2(mem_8__29_), .A3(n3146), .ZN(n4511) );
  NAND3_X2 U3606 ( .A1(n2771), .A2(mem_9__29_), .A3(n3146), .ZN(n4510) );
  NAND3_X2 U3607 ( .A1(n2285), .A2(mem_0__29_), .A3(n3146), .ZN(n4497) );
  NAND3_X2 U3608 ( .A1(n2770), .A2(mem_1__29_), .A3(n3146), .ZN(n4496) );
  NAND2_X2 U3609 ( .A1(n4539), .A2(n4538), .ZN(n4542) );
  NAND3_X2 U3610 ( .A1(n2248), .A2(mem_8__31_), .A3(n3144), .ZN(n4637) );
  NAND3_X2 U3611 ( .A1(n2771), .A2(mem_9__31_), .A3(n3146), .ZN(n4636) );
  NAND2_X2 U3612 ( .A1(n4670), .A2(n4669), .ZN(n4673) );
  NAND3_X2 U3613 ( .A1(n2294), .A2(mem_24__31_), .A3(n3138), .ZN(n4672) );
  NAND3_X2 U3614 ( .A1(n2771), .A2(mem_25__31_), .A3(n3151), .ZN(n4671) );
  NOR2_X2 U3615 ( .A1(n5704), .A2(n4692), .ZN(n4693) );
  NOR2_X2 U3616 ( .A1(n5704), .A2(n4740), .ZN(n4741) );
  NOR2_X2 U3617 ( .A1(n5704), .A2(n4788), .ZN(n4789) );
  NOR2_X2 U3618 ( .A1(n5704), .A2(n4836), .ZN(n4837) );
  NOR2_X2 U3619 ( .A1(n5704), .A2(n4884), .ZN(n4885) );
  NOR2_X2 U3620 ( .A1(n5704), .A2(n4932), .ZN(n4933) );
  NOR2_X2 U3621 ( .A1(n5704), .A2(n4980), .ZN(n4981) );
  NOR2_X2 U3622 ( .A1(n5704), .A2(n5028), .ZN(n5029) );
  NOR2_X2 U3623 ( .A1(n5704), .A2(n5076), .ZN(n5077) );
  NOR2_X2 U3624 ( .A1(n5704), .A2(n5124), .ZN(n5125) );
  NOR2_X2 U3625 ( .A1(n5704), .A2(n5223), .ZN(n5224) );
  NOR2_X2 U3626 ( .A1(n5704), .A2(n5271), .ZN(n5272) );
  NOR2_X2 U3627 ( .A1(n5704), .A2(n5319), .ZN(n5320) );
  NOR2_X2 U3628 ( .A1(n5704), .A2(n5367), .ZN(n5368) );
  INV_X4 U3629 ( .A(n2843), .ZN(n2345) );
  NOR2_X2 U3630 ( .A1(n5704), .A2(n5415), .ZN(n5416) );
  NOR2_X2 U3631 ( .A1(n5704), .A2(n5463), .ZN(n5464) );
  NOR2_X2 U3632 ( .A1(n5704), .A2(n5511), .ZN(n5512) );
  NOR2_X2 U3633 ( .A1(n5704), .A2(n5559), .ZN(n5560) );
  INV_X4 U3634 ( .A(n2843), .ZN(n2343) );
  NOR2_X2 U3635 ( .A1(n5704), .A2(n5607), .ZN(n5608) );
  INV_X4 U3636 ( .A(n2845), .ZN(n2339) );
  NOR2_X2 U3637 ( .A1(n5704), .A2(n5655), .ZN(n5656) );
  NOR2_X2 U3638 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  AOI211_X2 U3639 ( .C1(n5821), .C2(n5820), .A(n2385), .B(n2518), .ZN(n5831)
         );
  NOR3_X2 U3640 ( .A1(n5816), .A2(n5815), .A3(n5814), .ZN(n5821) );
  NOR3_X2 U3641 ( .A1(n5819), .A2(n5818), .A3(n5817), .ZN(n5820) );
  NOR3_X2 U3642 ( .A1(n5824), .A2(n5823), .A3(n5822), .ZN(n5829) );
  NOR3_X2 U3643 ( .A1(n5827), .A2(n5826), .A3(n5825), .ZN(n5828) );
  AOI211_X2 U3644 ( .C1(n5811), .C2(n5810), .A(n2384), .B(n2517), .ZN(n5812)
         );
  NOR3_X2 U3645 ( .A1(n5806), .A2(n5805), .A3(n5804), .ZN(n5811) );
  AOI211_X2 U3646 ( .C1(n5869), .C2(n5868), .A(n2389), .B(n2521), .ZN(n5870)
         );
  NOR3_X2 U3647 ( .A1(n5864), .A2(n5863), .A3(n5862), .ZN(n5869) );
  AOI211_X2 U3648 ( .C1(n5861), .C2(n5860), .A(n2388), .B(n2520), .ZN(n5871)
         );
  NOR3_X2 U3649 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(n5861) );
  AOI211_X2 U3650 ( .C1(n5851), .C2(n5850), .A(n2387), .B(n2519), .ZN(n5852)
         );
  NOR3_X2 U3651 ( .A1(n5846), .A2(n5845), .A3(n5844), .ZN(n5851) );
  AOI211_X2 U3652 ( .C1(n5891), .C2(n5890), .A(n2391), .B(n2522), .ZN(n5892)
         );
  NOR3_X2 U3653 ( .A1(n5886), .A2(n5885), .A3(n5884), .ZN(n5891) );
  AOI211_X2 U3654 ( .C1(n5883), .C2(n5882), .A(n2390), .B(n2545), .ZN(n5893)
         );
  NOR3_X2 U3655 ( .A1(n5878), .A2(n5877), .A3(n5876), .ZN(n5883) );
  AOI211_X2 U3656 ( .C1(n5901), .C2(n5900), .A(n2392), .B(n2523), .ZN(n5911)
         );
  AOI211_X2 U3657 ( .C1(n5909), .C2(n5908), .A(n2393), .B(n2524), .ZN(n5910)
         );
  AOI211_X2 U3658 ( .C1(n5931), .C2(n5930), .A(n2395), .B(n2525), .ZN(n5932)
         );
  NOR3_X2 U3659 ( .A1(n5929), .A2(n5928), .A3(n5927), .ZN(n5930) );
  NOR3_X2 U3660 ( .A1(n5926), .A2(n5925), .A3(n5924), .ZN(n5931) );
  AOI211_X2 U3661 ( .C1(n5923), .C2(n5922), .A(n2394), .B(n2546), .ZN(n5933)
         );
  NOR3_X2 U3662 ( .A1(n5918), .A2(n5917), .A3(n5916), .ZN(n5923) );
  NOR3_X2 U3663 ( .A1(n5921), .A2(n5920), .A3(n5919), .ZN(n5922) );
  AOI211_X2 U3664 ( .C1(n5949), .C2(n5948), .A(n2397), .B(n2527), .ZN(n5950)
         );
  AOI211_X2 U3665 ( .C1(n5941), .C2(n5940), .A(n2396), .B(n2526), .ZN(n5951)
         );
  NOR3_X2 U3666 ( .A1(n5944), .A2(n5943), .A3(n5942), .ZN(n5949) );
  AOI211_X2 U3667 ( .C1(n5989), .C2(n5988), .A(n2401), .B(n2530), .ZN(n5990)
         );
  NOR3_X2 U3668 ( .A1(n5984), .A2(n5983), .A3(n5982), .ZN(n5989) );
  AOI211_X2 U3669 ( .C1(n5981), .C2(n5980), .A(n2400), .B(n2529), .ZN(n5991)
         );
  NOR3_X2 U3670 ( .A1(n5976), .A2(n5975), .A3(n5974), .ZN(n5981) );
  AOI211_X2 U3671 ( .C1(n5971), .C2(n5970), .A(n2399), .B(n2528), .ZN(n5972)
         );
  AOI211_X2 U3672 ( .C1(n6011), .C2(n6010), .A(n2403), .B(n2531), .ZN(n6012)
         );
  NOR3_X2 U3673 ( .A1(n6009), .A2(n6008), .A3(n6007), .ZN(n6010) );
  AOI211_X2 U3674 ( .C1(n6003), .C2(n6002), .A(n2402), .B(n2548), .ZN(n6013)
         );
  NOR3_X2 U3675 ( .A1(n5998), .A2(n5997), .A3(n5996), .ZN(n6003) );
  NOR3_X2 U3676 ( .A1(n6001), .A2(n6000), .A3(n5999), .ZN(n6002) );
  AOI211_X2 U3677 ( .C1(n6021), .C2(n6020), .A(n2404), .B(n2532), .ZN(n6031)
         );
  AOI211_X2 U3678 ( .C1(n6029), .C2(n6028), .A(n2405), .B(n2533), .ZN(n6030)
         );
  AOI211_X2 U3679 ( .C1(n6069), .C2(n6068), .A(n2409), .B(n2536), .ZN(n6070)
         );
  NOR3_X2 U3680 ( .A1(n6064), .A2(n6063), .A3(n6062), .ZN(n6069) );
  AOI211_X2 U3681 ( .C1(n6061), .C2(n6060), .A(n2408), .B(n2535), .ZN(n6071)
         );
  NOR3_X2 U3682 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n6061) );
  NOR3_X2 U3683 ( .A1(n6059), .A2(n6058), .A3(n6057), .ZN(n6060) );
  AOI211_X2 U3684 ( .C1(n6051), .C2(n6050), .A(n2407), .B(n2534), .ZN(n6052)
         );
  AOI211_X2 U3685 ( .C1(n6043), .C2(n6042), .A(n2406), .B(n2549), .ZN(n6053)
         );
  AOI211_X2 U3686 ( .C1(n6109), .C2(n6108), .A(n2413), .B(n2539), .ZN(n6110)
         );
  NOR3_X2 U3687 ( .A1(n6104), .A2(n6103), .A3(n6102), .ZN(n6109) );
  AOI211_X2 U3688 ( .C1(n6101), .C2(n6100), .A(n2412), .B(n2538), .ZN(n6111)
         );
  NOR3_X2 U3689 ( .A1(n6096), .A2(n6095), .A3(n6094), .ZN(n6101) );
  NOR3_X2 U3690 ( .A1(n6099), .A2(n6098), .A3(n6097), .ZN(n6100) );
  AOI211_X2 U3691 ( .C1(n6091), .C2(n6090), .A(n2411), .B(n2537), .ZN(n6092)
         );
  AOI211_X2 U3692 ( .C1(n6083), .C2(n6082), .A(n2410), .B(n2550), .ZN(n6093)
         );
  AOI211_X2 U3693 ( .C1(n6151), .C2(n6150), .A(n2417), .B(n2542), .ZN(n6152)
         );
  NOR3_X2 U3694 ( .A1(n6144), .A2(n6143), .A3(n6142), .ZN(n6151) );
  AOI211_X2 U3695 ( .C1(n6141), .C2(n6140), .A(n2416), .B(n2541), .ZN(n6153)
         );
  NOR3_X2 U3696 ( .A1(n6136), .A2(n6135), .A3(n6134), .ZN(n6141) );
  AOI211_X2 U3697 ( .C1(n6131), .C2(n6130), .A(n2415), .B(n2540), .ZN(n6132)
         );
  AOI211_X2 U3698 ( .C1(n6123), .C2(n6122), .A(n2414), .B(n2551), .ZN(n6133)
         );
  OAI21_X2 U3699 ( .B1(n2938), .B2(n2982), .A(n745), .ZN(n1182) );
  OAI21_X2 U3700 ( .B1(n2936), .B2(n2984), .A(n734), .ZN(n1183) );
  OAI21_X2 U3701 ( .B1(n2934), .B2(n2983), .A(n723), .ZN(n1184) );
  OAI21_X2 U3702 ( .B1(n2932), .B2(n2982), .A(n720), .ZN(n1185) );
  OAI21_X2 U3703 ( .B1(n2930), .B2(n2982), .A(n719), .ZN(n1186) );
  OAI21_X2 U3704 ( .B1(n2928), .B2(n2982), .A(n718), .ZN(n1187) );
  OAI21_X2 U3705 ( .B1(n2926), .B2(n2982), .A(n717), .ZN(n1188) );
  OAI21_X2 U3706 ( .B1(n2924), .B2(n2982), .A(n716), .ZN(n1189) );
  OAI21_X2 U3707 ( .B1(n2922), .B2(n2982), .A(n715), .ZN(n1190) );
  OAI21_X2 U3708 ( .B1(n2920), .B2(n2982), .A(n714), .ZN(n1191) );
  OAI21_X2 U3709 ( .B1(n2918), .B2(n2982), .A(n744), .ZN(n1192) );
  OAI21_X2 U3710 ( .B1(n2916), .B2(n2982), .A(n743), .ZN(n1193) );
  OAI21_X2 U3711 ( .B1(n2914), .B2(n2982), .A(n742), .ZN(n1194) );
  OAI21_X2 U3712 ( .B1(n2912), .B2(n2983), .A(n741), .ZN(n1195) );
  OAI21_X2 U3713 ( .B1(n2910), .B2(n2983), .A(n740), .ZN(n1196) );
  OAI21_X2 U3714 ( .B1(n2908), .B2(n2983), .A(n739), .ZN(n1197) );
  OAI21_X2 U3715 ( .B1(n2906), .B2(n2984), .A(n738), .ZN(n1198) );
  OAI21_X2 U3716 ( .B1(n2904), .B2(n2984), .A(n737), .ZN(n1199) );
  OAI21_X2 U3717 ( .B1(n2902), .B2(n2984), .A(n736), .ZN(n1200) );
  OAI21_X2 U3718 ( .B1(n2900), .B2(n2984), .A(n735), .ZN(n1201) );
  OAI21_X2 U3719 ( .B1(n2898), .B2(n2984), .A(n733), .ZN(n1202) );
  OAI21_X2 U3720 ( .B1(n2896), .B2(n2983), .A(n732), .ZN(n1203) );
  OAI21_X2 U3721 ( .B1(n2894), .B2(n2984), .A(n731), .ZN(n1204) );
  OAI21_X2 U3722 ( .B1(n2892), .B2(n2984), .A(n730), .ZN(n1205) );
  OAI21_X2 U3723 ( .B1(n2890), .B2(n2983), .A(n729), .ZN(n1206) );
  OAI21_X2 U3724 ( .B1(n2888), .B2(n2983), .A(n728), .ZN(n1207) );
  OAI21_X2 U3725 ( .B1(n2886), .B2(n2983), .A(n727), .ZN(n1208) );
  OAI21_X2 U3726 ( .B1(n2884), .B2(n2983), .A(n726), .ZN(n1209) );
  OAI21_X2 U3727 ( .B1(n2882), .B2(n2983), .A(n725), .ZN(n1210) );
  OAI21_X2 U3728 ( .B1(n2880), .B2(n2983), .A(n724), .ZN(n1211) );
  OAI21_X2 U3729 ( .B1(n2878), .B2(n2983), .A(n722), .ZN(n1212) );
  OAI21_X2 U3730 ( .B1(n2876), .B2(n2982), .A(n721), .ZN(n1213) );
  OAI21_X2 U3731 ( .B1(n2939), .B2(n3025), .A(n376), .ZN(n1214) );
  OAI21_X2 U3732 ( .B1(n2937), .B2(n3027), .A(n365), .ZN(n1215) );
  OAI21_X2 U3733 ( .B1(n2935), .B2(n3026), .A(n354), .ZN(n1216) );
  OAI21_X2 U3734 ( .B1(n2933), .B2(n3025), .A(n351), .ZN(n1217) );
  OAI21_X2 U3735 ( .B1(n2931), .B2(n3025), .A(n350), .ZN(n1218) );
  OAI21_X2 U3736 ( .B1(n2929), .B2(n3025), .A(n349), .ZN(n1219) );
  OAI21_X2 U3737 ( .B1(n2927), .B2(n3025), .A(n348), .ZN(n1220) );
  OAI21_X2 U3738 ( .B1(n2925), .B2(n3025), .A(n347), .ZN(n1221) );
  OAI21_X2 U3739 ( .B1(n2923), .B2(n3025), .A(n346), .ZN(n1222) );
  OAI21_X2 U3740 ( .B1(n2921), .B2(n3025), .A(n345), .ZN(n1223) );
  OAI21_X2 U3741 ( .B1(n2919), .B2(n3025), .A(n375), .ZN(n1224) );
  OAI21_X2 U3742 ( .B1(n2917), .B2(n3025), .A(n374), .ZN(n1225) );
  OAI21_X2 U3743 ( .B1(n2915), .B2(n3025), .A(n373), .ZN(n1226) );
  OAI21_X2 U3744 ( .B1(n2913), .B2(n3026), .A(n372), .ZN(n1227) );
  OAI21_X2 U3745 ( .B1(n2911), .B2(n3026), .A(n371), .ZN(n1228) );
  OAI21_X2 U3746 ( .B1(n2909), .B2(n3026), .A(n370), .ZN(n1229) );
  OAI21_X2 U3747 ( .B1(n2907), .B2(n3027), .A(n369), .ZN(n1230) );
  OAI21_X2 U3748 ( .B1(n2905), .B2(n3027), .A(n368), .ZN(n1231) );
  OAI21_X2 U3749 ( .B1(n2903), .B2(n3027), .A(n367), .ZN(n1232) );
  OAI21_X2 U3750 ( .B1(n2901), .B2(n3027), .A(n366), .ZN(n1233) );
  OAI21_X2 U3751 ( .B1(n2899), .B2(n3027), .A(n364), .ZN(n1234) );
  OAI21_X2 U3752 ( .B1(n2897), .B2(n3026), .A(n363), .ZN(n1235) );
  OAI21_X2 U3753 ( .B1(n2895), .B2(n3027), .A(n362), .ZN(n1236) );
  OAI21_X2 U3754 ( .B1(n2893), .B2(n3027), .A(n361), .ZN(n1237) );
  OAI21_X2 U3755 ( .B1(n2891), .B2(n3026), .A(n360), .ZN(n1238) );
  OAI21_X2 U3756 ( .B1(n2889), .B2(n3026), .A(n359), .ZN(n1239) );
  OAI21_X2 U3757 ( .B1(n2887), .B2(n3026), .A(n358), .ZN(n1240) );
  OAI21_X2 U3758 ( .B1(n2885), .B2(n3026), .A(n357), .ZN(n1241) );
  OAI21_X2 U3759 ( .B1(n2883), .B2(n3026), .A(n356), .ZN(n1242) );
  OAI21_X2 U3760 ( .B1(n2881), .B2(n3026), .A(n355), .ZN(n1243) );
  OAI21_X2 U3761 ( .B1(n2879), .B2(n3026), .A(n353), .ZN(n1244) );
  OAI21_X2 U3762 ( .B1(n2877), .B2(n3025), .A(n352), .ZN(n1245) );
  OAI21_X2 U3763 ( .B1(n2939), .B2(n3036), .A(n275), .ZN(n1246) );
  OAI21_X2 U3764 ( .B1(n2937), .B2(n3038), .A(n264), .ZN(n1247) );
  OAI21_X2 U3765 ( .B1(n2935), .B2(n3037), .A(n253), .ZN(n1248) );
  OAI21_X2 U3766 ( .B1(n2933), .B2(n3036), .A(n250), .ZN(n1249) );
  OAI21_X2 U3767 ( .B1(n2931), .B2(n3036), .A(n249), .ZN(n1250) );
  OAI21_X2 U3768 ( .B1(n2929), .B2(n3036), .A(n248), .ZN(n1251) );
  OAI21_X2 U3769 ( .B1(n2927), .B2(n3036), .A(n247), .ZN(n1252) );
  OAI21_X2 U3770 ( .B1(n2925), .B2(n3036), .A(n246), .ZN(n1253) );
  OAI21_X2 U3771 ( .B1(n2923), .B2(n3036), .A(n245), .ZN(n1254) );
  OAI21_X2 U3772 ( .B1(n2921), .B2(n3036), .A(n244), .ZN(n1255) );
  OAI21_X2 U3773 ( .B1(n2919), .B2(n3036), .A(n274), .ZN(n1256) );
  OAI21_X2 U3774 ( .B1(n2917), .B2(n3036), .A(n273), .ZN(n1257) );
  OAI21_X2 U3775 ( .B1(n2915), .B2(n3036), .A(n272), .ZN(n1258) );
  OAI21_X2 U3776 ( .B1(n2913), .B2(n3037), .A(n271), .ZN(n1259) );
  OAI21_X2 U3777 ( .B1(n2911), .B2(n3037), .A(n270), .ZN(n1260) );
  OAI21_X2 U3778 ( .B1(n2909), .B2(n3037), .A(n269), .ZN(n1261) );
  OAI21_X2 U3779 ( .B1(n2907), .B2(n3038), .A(n268), .ZN(n1262) );
  OAI21_X2 U3780 ( .B1(n2905), .B2(n3038), .A(n267), .ZN(n1263) );
  OAI21_X2 U3781 ( .B1(n2903), .B2(n3038), .A(n266), .ZN(n1264) );
  OAI21_X2 U3782 ( .B1(n2901), .B2(n3038), .A(n265), .ZN(n1265) );
  OAI21_X2 U3783 ( .B1(n2899), .B2(n3038), .A(n263), .ZN(n1266) );
  OAI21_X2 U3784 ( .B1(n2897), .B2(n3037), .A(n262), .ZN(n1267) );
  OAI21_X2 U3785 ( .B1(n2895), .B2(n3038), .A(n261), .ZN(n1268) );
  OAI21_X2 U3786 ( .B1(n2893), .B2(n3038), .A(n260), .ZN(n1269) );
  OAI21_X2 U3787 ( .B1(n2891), .B2(n3037), .A(n259), .ZN(n1270) );
  OAI21_X2 U3788 ( .B1(n2889), .B2(n3037), .A(n258), .ZN(n1271) );
  OAI21_X2 U3789 ( .B1(n2887), .B2(n3037), .A(n257), .ZN(n1272) );
  OAI21_X2 U3790 ( .B1(n2885), .B2(n3037), .A(n256), .ZN(n1273) );
  OAI21_X2 U3791 ( .B1(n2883), .B2(n3037), .A(n255), .ZN(n1274) );
  OAI21_X2 U3792 ( .B1(n2881), .B2(n3037), .A(n254), .ZN(n1275) );
  OAI21_X2 U3793 ( .B1(n2879), .B2(n3037), .A(n252), .ZN(n1276) );
  OAI21_X2 U3794 ( .B1(n2877), .B2(n3036), .A(n251), .ZN(n1277) );
  OAI21_X2 U3795 ( .B1(n2939), .B2(n3039), .A(n240), .ZN(n1278) );
  OAI21_X2 U3796 ( .B1(n2936), .B2(n3041), .A(n229), .ZN(n1279) );
  OAI21_X2 U3797 ( .B1(n2935), .B2(n3040), .A(n218), .ZN(n1280) );
  OAI21_X2 U3798 ( .B1(n2933), .B2(n3039), .A(n215), .ZN(n1281) );
  OAI21_X2 U3799 ( .B1(n2931), .B2(n3039), .A(n214), .ZN(n1282) );
  OAI21_X2 U3800 ( .B1(n2929), .B2(n3039), .A(n213), .ZN(n1283) );
  OAI21_X2 U3801 ( .B1(n2927), .B2(n3039), .A(n212), .ZN(n1284) );
  OAI21_X2 U3802 ( .B1(n2925), .B2(n3039), .A(n211), .ZN(n1285) );
  OAI21_X2 U3803 ( .B1(n2923), .B2(n3039), .A(n210), .ZN(n1286) );
  OAI21_X2 U3804 ( .B1(n2920), .B2(n3039), .A(n209), .ZN(n1287) );
  OAI21_X2 U3805 ( .B1(n2918), .B2(n3039), .A(n239), .ZN(n1288) );
  OAI21_X2 U3806 ( .B1(n2917), .B2(n3039), .A(n238), .ZN(n1289) );
  OAI21_X2 U3807 ( .B1(n2914), .B2(n3039), .A(n237), .ZN(n1290) );
  OAI21_X2 U3808 ( .B1(n2913), .B2(n3040), .A(n236), .ZN(n1291) );
  OAI21_X2 U3809 ( .B1(n2911), .B2(n3040), .A(n235), .ZN(n1292) );
  OAI21_X2 U3810 ( .B1(n2909), .B2(n3040), .A(n234), .ZN(n1293) );
  OAI21_X2 U3811 ( .B1(n2907), .B2(n3041), .A(n233), .ZN(n1294) );
  OAI21_X2 U3812 ( .B1(n2905), .B2(n3041), .A(n232), .ZN(n1295) );
  OAI21_X2 U3813 ( .B1(n2903), .B2(n3041), .A(n231), .ZN(n1296) );
  OAI21_X2 U3814 ( .B1(n2901), .B2(n3041), .A(n230), .ZN(n1297) );
  OAI21_X2 U3815 ( .B1(n2899), .B2(n3041), .A(n228), .ZN(n1298) );
  OAI21_X2 U3816 ( .B1(n2897), .B2(n3040), .A(n227), .ZN(n1299) );
  OAI21_X2 U3817 ( .B1(n2894), .B2(n3041), .A(n226), .ZN(n1300) );
  OAI21_X2 U3818 ( .B1(n2892), .B2(n3041), .A(n225), .ZN(n1301) );
  OAI21_X2 U3819 ( .B1(n2890), .B2(n3040), .A(n224), .ZN(n1302) );
  OAI21_X2 U3820 ( .B1(n2888), .B2(n3040), .A(n223), .ZN(n1303) );
  OAI21_X2 U3821 ( .B1(n2886), .B2(n3040), .A(n222), .ZN(n1304) );
  OAI21_X2 U3822 ( .B1(n2884), .B2(n3040), .A(n221), .ZN(n1305) );
  OAI21_X2 U3823 ( .B1(n2882), .B2(n3040), .A(n220), .ZN(n1306) );
  OAI21_X2 U3824 ( .B1(n2880), .B2(n3040), .A(n219), .ZN(n1307) );
  OAI21_X2 U3825 ( .B1(n2878), .B2(n3040), .A(n217), .ZN(n1308) );
  OAI21_X2 U3826 ( .B1(n2876), .B2(n3039), .A(n216), .ZN(n1309) );
  OAI21_X2 U3827 ( .B1(n2939), .B2(n3042), .A(n207), .ZN(n1310) );
  OAI21_X2 U3828 ( .B1(n2936), .B2(n3044), .A(n196), .ZN(n1311) );
  OAI21_X2 U3829 ( .B1(n2935), .B2(n3043), .A(n185), .ZN(n1312) );
  OAI21_X2 U3830 ( .B1(n2933), .B2(n3042), .A(n182), .ZN(n1313) );
  OAI21_X2 U3831 ( .B1(n2931), .B2(n3042), .A(n181), .ZN(n1314) );
  OAI21_X2 U3832 ( .B1(n2929), .B2(n3042), .A(n180), .ZN(n1315) );
  OAI21_X2 U3833 ( .B1(n2927), .B2(n3042), .A(n179), .ZN(n1316) );
  OAI21_X2 U3834 ( .B1(n2925), .B2(n3042), .A(n178), .ZN(n1317) );
  OAI21_X2 U3835 ( .B1(n2923), .B2(n3042), .A(n177), .ZN(n1318) );
  OAI21_X2 U3836 ( .B1(n2920), .B2(n3042), .A(n176), .ZN(n1319) );
  OAI21_X2 U3837 ( .B1(n2919), .B2(n3042), .A(n206), .ZN(n1320) );
  OAI21_X2 U3838 ( .B1(n2917), .B2(n3042), .A(n205), .ZN(n1321) );
  OAI21_X2 U3839 ( .B1(n2915), .B2(n3042), .A(n204), .ZN(n1322) );
  OAI21_X2 U3840 ( .B1(n2913), .B2(n3043), .A(n203), .ZN(n1323) );
  OAI21_X2 U3841 ( .B1(n2911), .B2(n3043), .A(n202), .ZN(n1324) );
  OAI21_X2 U3842 ( .B1(n2909), .B2(n3043), .A(n201), .ZN(n1325) );
  OAI21_X2 U3843 ( .B1(n2907), .B2(n3044), .A(n200), .ZN(n1326) );
  OAI21_X2 U3844 ( .B1(n2905), .B2(n3044), .A(n199), .ZN(n1327) );
  OAI21_X2 U3845 ( .B1(n2903), .B2(n3044), .A(n198), .ZN(n1328) );
  OAI21_X2 U3846 ( .B1(n2901), .B2(n3044), .A(n197), .ZN(n1329) );
  OAI21_X2 U3847 ( .B1(n2899), .B2(n3044), .A(n195), .ZN(n1330) );
  OAI21_X2 U3848 ( .B1(n2897), .B2(n3043), .A(n194), .ZN(n1331) );
  OAI21_X2 U3849 ( .B1(n2894), .B2(n3044), .A(n193), .ZN(n1332) );
  OAI21_X2 U3850 ( .B1(n2893), .B2(n3044), .A(n192), .ZN(n1333) );
  OAI21_X2 U3851 ( .B1(n2891), .B2(n3043), .A(n191), .ZN(n1334) );
  OAI21_X2 U3852 ( .B1(n2889), .B2(n3043), .A(n190), .ZN(n1335) );
  OAI21_X2 U3853 ( .B1(n2887), .B2(n3043), .A(n189), .ZN(n1336) );
  OAI21_X2 U3854 ( .B1(n2885), .B2(n3043), .A(n188), .ZN(n1337) );
  OAI21_X2 U3855 ( .B1(n2883), .B2(n3043), .A(n187), .ZN(n1338) );
  OAI21_X2 U3856 ( .B1(n2881), .B2(n3043), .A(n186), .ZN(n1339) );
  OAI21_X2 U3857 ( .B1(n2879), .B2(n3043), .A(n184), .ZN(n1340) );
  OAI21_X2 U3858 ( .B1(n2877), .B2(n3042), .A(n183), .ZN(n1341) );
  OAI21_X2 U3859 ( .B1(n2938), .B2(n3045), .A(n173), .ZN(n1342) );
  OAI21_X2 U3860 ( .B1(n2937), .B2(n3047), .A(n162), .ZN(n1343) );
  OAI21_X2 U3861 ( .B1(n2934), .B2(n3046), .A(n151), .ZN(n1344) );
  OAI21_X2 U3862 ( .B1(n2932), .B2(n3045), .A(n148), .ZN(n1345) );
  OAI21_X2 U3863 ( .B1(n2930), .B2(n3045), .A(n147), .ZN(n1346) );
  OAI21_X2 U3864 ( .B1(n2928), .B2(n3045), .A(n146), .ZN(n1347) );
  OAI21_X2 U3865 ( .B1(n2926), .B2(n3045), .A(n145), .ZN(n1348) );
  OAI21_X2 U3866 ( .B1(n2924), .B2(n3045), .A(n144), .ZN(n1349) );
  OAI21_X2 U3867 ( .B1(n2922), .B2(n3045), .A(n143), .ZN(n1350) );
  OAI21_X2 U3868 ( .B1(n2921), .B2(n3045), .A(n142), .ZN(n1351) );
  OAI21_X2 U3869 ( .B1(n2919), .B2(n3045), .A(n172), .ZN(n1352) );
  OAI21_X2 U3870 ( .B1(n2916), .B2(n3045), .A(n171), .ZN(n1353) );
  OAI21_X2 U3871 ( .B1(n2915), .B2(n3045), .A(n170), .ZN(n1354) );
  OAI21_X2 U3872 ( .B1(n2912), .B2(n3046), .A(n169), .ZN(n1355) );
  OAI21_X2 U3873 ( .B1(n2910), .B2(n3046), .A(n168), .ZN(n1356) );
  OAI21_X2 U3874 ( .B1(n2908), .B2(n3046), .A(n167), .ZN(n1357) );
  OAI21_X2 U3875 ( .B1(n2906), .B2(n3047), .A(n166), .ZN(n1358) );
  OAI21_X2 U3876 ( .B1(n2904), .B2(n3047), .A(n165), .ZN(n1359) );
  OAI21_X2 U3877 ( .B1(n2902), .B2(n3047), .A(n164), .ZN(n1360) );
  OAI21_X2 U3878 ( .B1(n2900), .B2(n3047), .A(n163), .ZN(n1361) );
  OAI21_X2 U3879 ( .B1(n2898), .B2(n3047), .A(n161), .ZN(n1362) );
  OAI21_X2 U3880 ( .B1(n2896), .B2(n3046), .A(n160), .ZN(n1363) );
  OAI21_X2 U3881 ( .B1(n2895), .B2(n3047), .A(n159), .ZN(n1364) );
  OAI21_X2 U3882 ( .B1(n2893), .B2(n3047), .A(n158), .ZN(n1365) );
  OAI21_X2 U3883 ( .B1(n2891), .B2(n3046), .A(n157), .ZN(n1366) );
  OAI21_X2 U3884 ( .B1(n2889), .B2(n3046), .A(n156), .ZN(n1367) );
  OAI21_X2 U3885 ( .B1(n2887), .B2(n3046), .A(n155), .ZN(n1368) );
  OAI21_X2 U3886 ( .B1(n2885), .B2(n3046), .A(n154), .ZN(n1369) );
  OAI21_X2 U3887 ( .B1(n2883), .B2(n3046), .A(n153), .ZN(n1370) );
  OAI21_X2 U3888 ( .B1(n2881), .B2(n3046), .A(n152), .ZN(n1371) );
  OAI21_X2 U3889 ( .B1(n2879), .B2(n3046), .A(n150), .ZN(n1372) );
  OAI21_X2 U3890 ( .B1(n2877), .B2(n3045), .A(n149), .ZN(n1373) );
  OAI21_X2 U3891 ( .B1(n2939), .B2(n3048), .A(n138), .ZN(n1374) );
  OAI21_X2 U3892 ( .B1(n2937), .B2(n3050), .A(n127), .ZN(n1375) );
  OAI21_X2 U3893 ( .B1(n2935), .B2(n3049), .A(n116), .ZN(n1376) );
  OAI21_X2 U3894 ( .B1(n2933), .B2(n3048), .A(n113), .ZN(n1377) );
  OAI21_X2 U3895 ( .B1(n2931), .B2(n3048), .A(n112), .ZN(n1378) );
  OAI21_X2 U3896 ( .B1(n2929), .B2(n3048), .A(n111), .ZN(n1379) );
  OAI21_X2 U3897 ( .B1(n2927), .B2(n3048), .A(n110), .ZN(n1380) );
  OAI21_X2 U3898 ( .B1(n2925), .B2(n3048), .A(n109), .ZN(n1381) );
  OAI21_X2 U3899 ( .B1(n2923), .B2(n3048), .A(n108), .ZN(n1382) );
  OAI21_X2 U3900 ( .B1(n2920), .B2(n3048), .A(n107), .ZN(n1383) );
  OAI21_X2 U3901 ( .B1(n2918), .B2(n3048), .A(n137), .ZN(n1384) );
  OAI21_X2 U3902 ( .B1(n2917), .B2(n3048), .A(n136), .ZN(n1385) );
  OAI21_X2 U3903 ( .B1(n2915), .B2(n3048), .A(n135), .ZN(n1386) );
  OAI21_X2 U3904 ( .B1(n2913), .B2(n3049), .A(n134), .ZN(n1387) );
  OAI21_X2 U3905 ( .B1(n2911), .B2(n3049), .A(n133), .ZN(n1388) );
  OAI21_X2 U3906 ( .B1(n2909), .B2(n3049), .A(n132), .ZN(n1389) );
  OAI21_X2 U3907 ( .B1(n2907), .B2(n3050), .A(n131), .ZN(n1390) );
  OAI21_X2 U3908 ( .B1(n2905), .B2(n3050), .A(n130), .ZN(n1391) );
  OAI21_X2 U3909 ( .B1(n2903), .B2(n3050), .A(n129), .ZN(n1392) );
  OAI21_X2 U3910 ( .B1(n2901), .B2(n3050), .A(n128), .ZN(n1393) );
  OAI21_X2 U3911 ( .B1(n2899), .B2(n3050), .A(n126), .ZN(n1394) );
  OAI21_X2 U3912 ( .B1(n2897), .B2(n3049), .A(n125), .ZN(n1395) );
  OAI21_X2 U3913 ( .B1(n2895), .B2(n3050), .A(n124), .ZN(n1396) );
  OAI21_X2 U3914 ( .B1(n2892), .B2(n3050), .A(n123), .ZN(n1397) );
  OAI21_X2 U3915 ( .B1(n2890), .B2(n3049), .A(n122), .ZN(n1398) );
  OAI21_X2 U3916 ( .B1(n2888), .B2(n3049), .A(n121), .ZN(n1399) );
  OAI21_X2 U3917 ( .B1(n2886), .B2(n3049), .A(n120), .ZN(n1400) );
  OAI21_X2 U3918 ( .B1(n2884), .B2(n3049), .A(n119), .ZN(n1401) );
  OAI21_X2 U3919 ( .B1(n2882), .B2(n3049), .A(n118), .ZN(n1402) );
  OAI21_X2 U3920 ( .B1(n2880), .B2(n3049), .A(n117), .ZN(n1403) );
  OAI21_X2 U3921 ( .B1(n2878), .B2(n3049), .A(n115), .ZN(n1404) );
  OAI21_X2 U3922 ( .B1(n2876), .B2(n3048), .A(n114), .ZN(n1405) );
  OAI21_X2 U3923 ( .B1(n2938), .B2(n3052), .A(n104), .ZN(n1406) );
  OAI21_X2 U3924 ( .B1(n2937), .B2(n3054), .A(n93), .ZN(n1407) );
  OAI21_X2 U3925 ( .B1(n2934), .B2(n3053), .A(n82), .ZN(n1408) );
  OAI21_X2 U3926 ( .B1(n2932), .B2(n3052), .A(n79), .ZN(n1409) );
  OAI21_X2 U3927 ( .B1(n2930), .B2(n3052), .A(n78), .ZN(n1410) );
  OAI21_X2 U3928 ( .B1(n2928), .B2(n3052), .A(n77), .ZN(n1411) );
  OAI21_X2 U3929 ( .B1(n2926), .B2(n3052), .A(n76), .ZN(n1412) );
  OAI21_X2 U3930 ( .B1(n2924), .B2(n3052), .A(n75), .ZN(n1413) );
  OAI21_X2 U3931 ( .B1(n2922), .B2(n3052), .A(n74), .ZN(n1414) );
  OAI21_X2 U3932 ( .B1(n2920), .B2(n3052), .A(n73), .ZN(n1415) );
  OAI21_X2 U3933 ( .B1(n2919), .B2(n3052), .A(n103), .ZN(n1416) );
  OAI21_X2 U3934 ( .B1(n2916), .B2(n3052), .A(n102), .ZN(n1417) );
  OAI21_X2 U3935 ( .B1(n2914), .B2(n3052), .A(n101), .ZN(n1418) );
  OAI21_X2 U3936 ( .B1(n2912), .B2(n3053), .A(n100), .ZN(n1419) );
  OAI21_X2 U3937 ( .B1(n2910), .B2(n3053), .A(n99), .ZN(n1420) );
  OAI21_X2 U3938 ( .B1(n2908), .B2(n3053), .A(n98), .ZN(n1421) );
  OAI21_X2 U3939 ( .B1(n2906), .B2(n3054), .A(n97), .ZN(n1422) );
  OAI21_X2 U3940 ( .B1(n2904), .B2(n3054), .A(n96), .ZN(n1423) );
  OAI21_X2 U3941 ( .B1(n2902), .B2(n3054), .A(n95), .ZN(n1424) );
  OAI21_X2 U3942 ( .B1(n2900), .B2(n3054), .A(n94), .ZN(n1425) );
  OAI21_X2 U3943 ( .B1(n2898), .B2(n3054), .A(n92), .ZN(n1426) );
  OAI21_X2 U3944 ( .B1(n2896), .B2(n3053), .A(n91), .ZN(n1427) );
  OAI21_X2 U3945 ( .B1(n2895), .B2(n3054), .A(n90), .ZN(n1428) );
  OAI21_X2 U3946 ( .B1(n2893), .B2(n3054), .A(n89), .ZN(n1429) );
  OAI21_X2 U3947 ( .B1(n2891), .B2(n3053), .A(n88), .ZN(n1430) );
  OAI21_X2 U3948 ( .B1(n2889), .B2(n3053), .A(n87), .ZN(n1431) );
  OAI21_X2 U3949 ( .B1(n2887), .B2(n3053), .A(n86), .ZN(n1432) );
  OAI21_X2 U3950 ( .B1(n2885), .B2(n3053), .A(n85), .ZN(n1433) );
  OAI21_X2 U3951 ( .B1(n2883), .B2(n3053), .A(n84), .ZN(n1434) );
  OAI21_X2 U3952 ( .B1(n2881), .B2(n3053), .A(n83), .ZN(n1435) );
  OAI21_X2 U3953 ( .B1(n2879), .B2(n3053), .A(n81), .ZN(n1436) );
  OAI21_X2 U3954 ( .B1(n2877), .B2(n3052), .A(n80), .ZN(n1437) );
  OAI21_X2 U3955 ( .B1(n3056), .B2(n2938), .A(n69), .ZN(n1438) );
  OAI21_X2 U3956 ( .B1(n3058), .B2(n2936), .A(n47), .ZN(n1439) );
  OAI21_X2 U3957 ( .B1(n3056), .B2(n2934), .A(n25), .ZN(n1440) );
  OAI21_X2 U3958 ( .B1(n3056), .B2(n2932), .A(n19), .ZN(n1441) );
  OAI21_X2 U3959 ( .B1(n3056), .B2(n2930), .A(n17), .ZN(n1442) );
  OAI21_X2 U3960 ( .B1(n3056), .B2(n2928), .A(n15), .ZN(n1443) );
  OAI21_X2 U3961 ( .B1(n3056), .B2(n2926), .A(n13), .ZN(n1444) );
  OAI21_X2 U3962 ( .B1(n3056), .B2(n2924), .A(n11), .ZN(n1445) );
  OAI21_X2 U3963 ( .B1(n3056), .B2(n2922), .A(n9), .ZN(n1446) );
  OAI21_X2 U3964 ( .B1(n2921), .B2(n3058), .A(n7), .ZN(n1447) );
  OAI21_X2 U3965 ( .B1(n3056), .B2(n2918), .A(n67), .ZN(n1448) );
  OAI21_X2 U3966 ( .B1(n3056), .B2(n2916), .A(n65), .ZN(n1449) );
  OAI21_X2 U3967 ( .B1(n3056), .B2(n2914), .A(n63), .ZN(n1450) );
  OAI21_X2 U3968 ( .B1(n3057), .B2(n2912), .A(n61), .ZN(n1451) );
  OAI21_X2 U3969 ( .B1(n3057), .B2(n2910), .A(n59), .ZN(n1452) );
  OAI21_X2 U3970 ( .B1(n3057), .B2(n2908), .A(n57), .ZN(n1453) );
  OAI21_X2 U3971 ( .B1(n3058), .B2(n2906), .A(n55), .ZN(n1454) );
  OAI21_X2 U3972 ( .B1(n3058), .B2(n2904), .A(n53), .ZN(n1455) );
  OAI21_X2 U3973 ( .B1(n3057), .B2(n2902), .A(n51), .ZN(n1456) );
  OAI21_X2 U3974 ( .B1(n3058), .B2(n2900), .A(n49), .ZN(n1457) );
  OAI21_X2 U3975 ( .B1(n3058), .B2(n2898), .A(n45), .ZN(n1458) );
  OAI21_X2 U3976 ( .B1(n3057), .B2(n2896), .A(n43), .ZN(n1459) );
  OAI21_X2 U3977 ( .B1(n3058), .B2(n2894), .A(n41), .ZN(n1460) );
  OAI21_X2 U3978 ( .B1(n3058), .B2(n2892), .A(n39), .ZN(n1461) );
  OAI21_X2 U3979 ( .B1(n3057), .B2(n2890), .A(n37), .ZN(n1462) );
  OAI21_X2 U3980 ( .B1(n3057), .B2(n2888), .A(n35), .ZN(n1463) );
  OAI21_X2 U3981 ( .B1(n3057), .B2(n2886), .A(n33), .ZN(n1464) );
  OAI21_X2 U3982 ( .B1(n3057), .B2(n2884), .A(n31), .ZN(n1465) );
  OAI21_X2 U3983 ( .B1(n3057), .B2(n2882), .A(n29), .ZN(n1466) );
  OAI21_X2 U3984 ( .B1(n3057), .B2(n2880), .A(n27), .ZN(n1467) );
  OAI21_X2 U3985 ( .B1(n3057), .B2(n2878), .A(n23), .ZN(n1468) );
  OAI21_X2 U3986 ( .B1(n3056), .B2(n2876), .A(n21), .ZN(n1469) );
  OAI21_X2 U3987 ( .B1(n2938), .B2(n2943), .A(n1080), .ZN(n1470) );
  OAI21_X2 U3988 ( .B1(n2936), .B2(n2945), .A(n1069), .ZN(n1471) );
  OAI21_X2 U3989 ( .B1(n2934), .B2(n2944), .A(n1058), .ZN(n1472) );
  OAI21_X2 U3990 ( .B1(n2932), .B2(n2943), .A(n1055), .ZN(n1473) );
  OAI21_X2 U3991 ( .B1(n2930), .B2(n2943), .A(n1054), .ZN(n1474) );
  OAI21_X2 U3992 ( .B1(n2928), .B2(n2943), .A(n1053), .ZN(n1475) );
  OAI21_X2 U3993 ( .B1(n2926), .B2(n2943), .A(n1052), .ZN(n1476) );
  OAI21_X2 U3994 ( .B1(n2924), .B2(n2943), .A(n1051), .ZN(n1477) );
  OAI21_X2 U3995 ( .B1(n2922), .B2(n2943), .A(n1050), .ZN(n1478) );
  OAI21_X2 U3996 ( .B1(n2920), .B2(n2943), .A(n1049), .ZN(n1479) );
  OAI21_X2 U3997 ( .B1(n2918), .B2(n2943), .A(n1079), .ZN(n1480) );
  OAI21_X2 U3998 ( .B1(n2916), .B2(n2943), .A(n1078), .ZN(n1481) );
  OAI21_X2 U3999 ( .B1(n2914), .B2(n2943), .A(n1077), .ZN(n1482) );
  OAI21_X2 U4000 ( .B1(n2912), .B2(n2944), .A(n1076), .ZN(n1483) );
  OAI21_X2 U4001 ( .B1(n2910), .B2(n2944), .A(n1075), .ZN(n1484) );
  OAI21_X2 U4002 ( .B1(n2908), .B2(n2944), .A(n1074), .ZN(n1485) );
  OAI21_X2 U4003 ( .B1(n2906), .B2(n2945), .A(n1073), .ZN(n1486) );
  OAI21_X2 U4004 ( .B1(n2904), .B2(n2945), .A(n1072), .ZN(n1487) );
  OAI21_X2 U4005 ( .B1(n2902), .B2(n2945), .A(n1071), .ZN(n1488) );
  OAI21_X2 U4006 ( .B1(n2900), .B2(n2945), .A(n1070), .ZN(n1489) );
  OAI21_X2 U4007 ( .B1(n2898), .B2(n2945), .A(n1068), .ZN(n1490) );
  OAI21_X2 U4008 ( .B1(n2896), .B2(n2944), .A(n1067), .ZN(n1491) );
  OAI21_X2 U4009 ( .B1(n2894), .B2(n2945), .A(n1066), .ZN(n1492) );
  OAI21_X2 U4010 ( .B1(n2892), .B2(n2945), .A(n1065), .ZN(n1493) );
  OAI21_X2 U4011 ( .B1(n2890), .B2(n2944), .A(n1064), .ZN(n1494) );
  OAI21_X2 U4012 ( .B1(n2888), .B2(n2944), .A(n1063), .ZN(n1495) );
  OAI21_X2 U4013 ( .B1(n2886), .B2(n2944), .A(n1062), .ZN(n1496) );
  OAI21_X2 U4014 ( .B1(n2884), .B2(n2944), .A(n1061), .ZN(n1497) );
  OAI21_X2 U4015 ( .B1(n2882), .B2(n2944), .A(n1060), .ZN(n1498) );
  OAI21_X2 U4016 ( .B1(n2880), .B2(n2944), .A(n1059), .ZN(n1499) );
  OAI21_X2 U4017 ( .B1(n2878), .B2(n2944), .A(n1057), .ZN(n1500) );
  OAI21_X2 U4018 ( .B1(n2876), .B2(n2943), .A(n1056), .ZN(n1501) );
  OAI21_X2 U4019 ( .B1(n2938), .B2(n2947), .A(n1047), .ZN(n1502) );
  OAI21_X2 U4020 ( .B1(n2936), .B2(n2949), .A(n1036), .ZN(n1503) );
  OAI21_X2 U4021 ( .B1(n2934), .B2(n2948), .A(n1025), .ZN(n1504) );
  OAI21_X2 U4022 ( .B1(n2932), .B2(n2947), .A(n1022), .ZN(n1505) );
  OAI21_X2 U4023 ( .B1(n2930), .B2(n2947), .A(n1021), .ZN(n1506) );
  OAI21_X2 U4024 ( .B1(n2928), .B2(n2947), .A(n1020), .ZN(n1507) );
  OAI21_X2 U4025 ( .B1(n2926), .B2(n2947), .A(n1019), .ZN(n1508) );
  OAI21_X2 U4026 ( .B1(n2924), .B2(n2947), .A(n1018), .ZN(n1509) );
  OAI21_X2 U4027 ( .B1(n2922), .B2(n2947), .A(n1017), .ZN(n1510) );
  OAI21_X2 U4028 ( .B1(n2920), .B2(n2947), .A(n1016), .ZN(n1511) );
  OAI21_X2 U4029 ( .B1(n2918), .B2(n2947), .A(n1046), .ZN(n1512) );
  OAI21_X2 U4030 ( .B1(n2916), .B2(n2947), .A(n1045), .ZN(n1513) );
  OAI21_X2 U4031 ( .B1(n2914), .B2(n2947), .A(n1044), .ZN(n1514) );
  OAI21_X2 U4032 ( .B1(n2912), .B2(n2948), .A(n1043), .ZN(n1515) );
  OAI21_X2 U4033 ( .B1(n2910), .B2(n2948), .A(n1042), .ZN(n1516) );
  OAI21_X2 U4034 ( .B1(n2908), .B2(n2948), .A(n1041), .ZN(n1517) );
  OAI21_X2 U4035 ( .B1(n2906), .B2(n2949), .A(n1040), .ZN(n1518) );
  OAI21_X2 U4036 ( .B1(n2904), .B2(n2949), .A(n1039), .ZN(n1519) );
  OAI21_X2 U4037 ( .B1(n2902), .B2(n2949), .A(n1038), .ZN(n1520) );
  OAI21_X2 U4038 ( .B1(n2900), .B2(n2949), .A(n1037), .ZN(n1521) );
  OAI21_X2 U4039 ( .B1(n2898), .B2(n2949), .A(n1035), .ZN(n1522) );
  OAI21_X2 U4040 ( .B1(n2896), .B2(n2948), .A(n1034), .ZN(n1523) );
  OAI21_X2 U4041 ( .B1(n2894), .B2(n2949), .A(n1033), .ZN(n1524) );
  OAI21_X2 U4042 ( .B1(n2892), .B2(n2949), .A(n1032), .ZN(n1525) );
  OAI21_X2 U4043 ( .B1(n2890), .B2(n2948), .A(n1031), .ZN(n1526) );
  OAI21_X2 U4044 ( .B1(n2888), .B2(n2948), .A(n1030), .ZN(n1527) );
  OAI21_X2 U4045 ( .B1(n2886), .B2(n2948), .A(n1029), .ZN(n1528) );
  OAI21_X2 U4046 ( .B1(n2884), .B2(n2948), .A(n1028), .ZN(n1529) );
  OAI21_X2 U4047 ( .B1(n2882), .B2(n2948), .A(n1027), .ZN(n1530) );
  OAI21_X2 U4048 ( .B1(n2880), .B2(n2948), .A(n1026), .ZN(n1531) );
  OAI21_X2 U4049 ( .B1(n2878), .B2(n2948), .A(n1024), .ZN(n1532) );
  OAI21_X2 U4050 ( .B1(n2876), .B2(n2947), .A(n1023), .ZN(n1533) );
  OAI21_X2 U4051 ( .B1(n2938), .B2(n2951), .A(n1013), .ZN(n1534) );
  OAI21_X2 U4052 ( .B1(n2936), .B2(n2953), .A(n1002), .ZN(n1535) );
  OAI21_X2 U4053 ( .B1(n2934), .B2(n2952), .A(n991), .ZN(n1536) );
  OAI21_X2 U4054 ( .B1(n2932), .B2(n2951), .A(n988), .ZN(n1537) );
  OAI21_X2 U4055 ( .B1(n2930), .B2(n2951), .A(n987), .ZN(n1538) );
  OAI21_X2 U4056 ( .B1(n2928), .B2(n2951), .A(n986), .ZN(n1539) );
  OAI21_X2 U4057 ( .B1(n2926), .B2(n2951), .A(n985), .ZN(n1540) );
  OAI21_X2 U4058 ( .B1(n2924), .B2(n2951), .A(n984), .ZN(n1541) );
  OAI21_X2 U4059 ( .B1(n2922), .B2(n2951), .A(n983), .ZN(n1542) );
  OAI21_X2 U4060 ( .B1(n2920), .B2(n2951), .A(n982), .ZN(n1543) );
  OAI21_X2 U4061 ( .B1(n2918), .B2(n2951), .A(n1012), .ZN(n1544) );
  OAI21_X2 U4062 ( .B1(n2916), .B2(n2951), .A(n1011), .ZN(n1545) );
  OAI21_X2 U4063 ( .B1(n2914), .B2(n2951), .A(n1010), .ZN(n1546) );
  OAI21_X2 U4064 ( .B1(n2912), .B2(n2952), .A(n1009), .ZN(n1547) );
  OAI21_X2 U4065 ( .B1(n2910), .B2(n2952), .A(n1008), .ZN(n1548) );
  OAI21_X2 U4066 ( .B1(n2908), .B2(n2952), .A(n1007), .ZN(n1549) );
  OAI21_X2 U4067 ( .B1(n2906), .B2(n2953), .A(n1006), .ZN(n1550) );
  OAI21_X2 U4068 ( .B1(n2904), .B2(n2953), .A(n1005), .ZN(n1551) );
  OAI21_X2 U4069 ( .B1(n2902), .B2(n2953), .A(n1004), .ZN(n1552) );
  OAI21_X2 U4070 ( .B1(n2900), .B2(n2953), .A(n1003), .ZN(n1553) );
  OAI21_X2 U4071 ( .B1(n2898), .B2(n2953), .A(n1001), .ZN(n1554) );
  OAI21_X2 U4072 ( .B1(n2896), .B2(n2952), .A(n1000), .ZN(n1555) );
  OAI21_X2 U4073 ( .B1(n2894), .B2(n2953), .A(n999), .ZN(n1556) );
  OAI21_X2 U4074 ( .B1(n2892), .B2(n2953), .A(n998), .ZN(n1557) );
  OAI21_X2 U4075 ( .B1(n2890), .B2(n2952), .A(n997), .ZN(n1558) );
  OAI21_X2 U4076 ( .B1(n2888), .B2(n2952), .A(n996), .ZN(n1559) );
  OAI21_X2 U4077 ( .B1(n2886), .B2(n2952), .A(n995), .ZN(n1560) );
  OAI21_X2 U4078 ( .B1(n2884), .B2(n2952), .A(n994), .ZN(n1561) );
  OAI21_X2 U4079 ( .B1(n2882), .B2(n2952), .A(n993), .ZN(n1562) );
  OAI21_X2 U4080 ( .B1(n2880), .B2(n2952), .A(n992), .ZN(n1563) );
  OAI21_X2 U4081 ( .B1(n2878), .B2(n2952), .A(n990), .ZN(n1564) );
  OAI21_X2 U4082 ( .B1(n2876), .B2(n2951), .A(n989), .ZN(n1565) );
  OAI21_X2 U4083 ( .B1(n2938), .B2(n2954), .A(n979), .ZN(n1566) );
  OAI21_X2 U4084 ( .B1(n2936), .B2(n2956), .A(n968), .ZN(n1567) );
  OAI21_X2 U4085 ( .B1(n2934), .B2(n2955), .A(n957), .ZN(n1568) );
  OAI21_X2 U4086 ( .B1(n2932), .B2(n2954), .A(n954), .ZN(n1569) );
  OAI21_X2 U4087 ( .B1(n2930), .B2(n2954), .A(n953), .ZN(n1570) );
  OAI21_X2 U4088 ( .B1(n2928), .B2(n2954), .A(n952), .ZN(n1571) );
  OAI21_X2 U4089 ( .B1(n2926), .B2(n2954), .A(n951), .ZN(n1572) );
  OAI21_X2 U4090 ( .B1(n2924), .B2(n2954), .A(n950), .ZN(n1573) );
  OAI21_X2 U4091 ( .B1(n2922), .B2(n2954), .A(n949), .ZN(n1574) );
  OAI21_X2 U4092 ( .B1(n2920), .B2(n2954), .A(n948), .ZN(n1575) );
  OAI21_X2 U4093 ( .B1(n2918), .B2(n2954), .A(n978), .ZN(n1576) );
  OAI21_X2 U4094 ( .B1(n2916), .B2(n2954), .A(n977), .ZN(n1577) );
  OAI21_X2 U4095 ( .B1(n2914), .B2(n2954), .A(n976), .ZN(n1578) );
  OAI21_X2 U4096 ( .B1(n2912), .B2(n2955), .A(n975), .ZN(n1579) );
  OAI21_X2 U4097 ( .B1(n2910), .B2(n2955), .A(n974), .ZN(n1580) );
  OAI21_X2 U4098 ( .B1(n2908), .B2(n2955), .A(n973), .ZN(n1581) );
  OAI21_X2 U4099 ( .B1(n2906), .B2(n2956), .A(n972), .ZN(n1582) );
  OAI21_X2 U4100 ( .B1(n2904), .B2(n2956), .A(n971), .ZN(n1583) );
  OAI21_X2 U4101 ( .B1(n2902), .B2(n2956), .A(n970), .ZN(n1584) );
  OAI21_X2 U4102 ( .B1(n2900), .B2(n2956), .A(n969), .ZN(n1585) );
  OAI21_X2 U4103 ( .B1(n2898), .B2(n2956), .A(n967), .ZN(n1586) );
  OAI21_X2 U4104 ( .B1(n2896), .B2(n2955), .A(n966), .ZN(n1587) );
  OAI21_X2 U4105 ( .B1(n2894), .B2(n2956), .A(n965), .ZN(n1588) );
  OAI21_X2 U4106 ( .B1(n2892), .B2(n2956), .A(n964), .ZN(n1589) );
  OAI21_X2 U4107 ( .B1(n2890), .B2(n2955), .A(n963), .ZN(n1590) );
  OAI21_X2 U4108 ( .B1(n2888), .B2(n2955), .A(n962), .ZN(n1591) );
  OAI21_X2 U4109 ( .B1(n2886), .B2(n2955), .A(n961), .ZN(n1592) );
  OAI21_X2 U4110 ( .B1(n2884), .B2(n2955), .A(n960), .ZN(n1593) );
  OAI21_X2 U4111 ( .B1(n2882), .B2(n2955), .A(n959), .ZN(n1594) );
  OAI21_X2 U4112 ( .B1(n2880), .B2(n2955), .A(n958), .ZN(n1595) );
  OAI21_X2 U4113 ( .B1(n2878), .B2(n2955), .A(n956), .ZN(n1596) );
  OAI21_X2 U4114 ( .B1(n2876), .B2(n2954), .A(n955), .ZN(n1597) );
  OAI21_X2 U4115 ( .B1(n2938), .B2(n2959), .A(n946), .ZN(n1598) );
  OAI21_X2 U4116 ( .B1(n2936), .B2(n2961), .A(n935), .ZN(n1599) );
  OAI21_X2 U4117 ( .B1(n2934), .B2(n2960), .A(n924), .ZN(n1600) );
  OAI21_X2 U4118 ( .B1(n2932), .B2(n2959), .A(n921), .ZN(n1601) );
  OAI21_X2 U4119 ( .B1(n2930), .B2(n2959), .A(n920), .ZN(n1602) );
  OAI21_X2 U4120 ( .B1(n2928), .B2(n2959), .A(n919), .ZN(n1603) );
  OAI21_X2 U4121 ( .B1(n2926), .B2(n2959), .A(n918), .ZN(n1604) );
  OAI21_X2 U4122 ( .B1(n2924), .B2(n2959), .A(n917), .ZN(n1605) );
  OAI21_X2 U4123 ( .B1(n2922), .B2(n2959), .A(n916), .ZN(n1606) );
  OAI21_X2 U4124 ( .B1(n2920), .B2(n2959), .A(n915), .ZN(n1607) );
  OAI21_X2 U4125 ( .B1(n2918), .B2(n2959), .A(n945), .ZN(n1608) );
  OAI21_X2 U4126 ( .B1(n2916), .B2(n2959), .A(n944), .ZN(n1609) );
  OAI21_X2 U4127 ( .B1(n2914), .B2(n2959), .A(n943), .ZN(n1610) );
  OAI21_X2 U4128 ( .B1(n2912), .B2(n2960), .A(n942), .ZN(n1611) );
  OAI21_X2 U4129 ( .B1(n2910), .B2(n2960), .A(n941), .ZN(n1612) );
  OAI21_X2 U4130 ( .B1(n2908), .B2(n2960), .A(n940), .ZN(n1613) );
  OAI21_X2 U4131 ( .B1(n2906), .B2(n2961), .A(n939), .ZN(n1614) );
  OAI21_X2 U4132 ( .B1(n2904), .B2(n2961), .A(n938), .ZN(n1615) );
  OAI21_X2 U4133 ( .B1(n2902), .B2(n2961), .A(n937), .ZN(n1616) );
  OAI21_X2 U4134 ( .B1(n2900), .B2(n2961), .A(n936), .ZN(n1617) );
  OAI21_X2 U4135 ( .B1(n2898), .B2(n2961), .A(n934), .ZN(n1618) );
  OAI21_X2 U4136 ( .B1(n2896), .B2(n2960), .A(n933), .ZN(n1619) );
  OAI21_X2 U4137 ( .B1(n2894), .B2(n2961), .A(n932), .ZN(n1620) );
  OAI21_X2 U4138 ( .B1(n2892), .B2(n2961), .A(n931), .ZN(n1621) );
  OAI21_X2 U4139 ( .B1(n2890), .B2(n2960), .A(n930), .ZN(n1622) );
  OAI21_X2 U4140 ( .B1(n2888), .B2(n2960), .A(n929), .ZN(n1623) );
  OAI21_X2 U4141 ( .B1(n2886), .B2(n2960), .A(n928), .ZN(n1624) );
  OAI21_X2 U4142 ( .B1(n2884), .B2(n2960), .A(n927), .ZN(n1625) );
  OAI21_X2 U4143 ( .B1(n2882), .B2(n2960), .A(n926), .ZN(n1626) );
  OAI21_X2 U4144 ( .B1(n2880), .B2(n2960), .A(n925), .ZN(n1627) );
  OAI21_X2 U4145 ( .B1(n2878), .B2(n2960), .A(n923), .ZN(n1628) );
  OAI21_X2 U4146 ( .B1(n2876), .B2(n2959), .A(n922), .ZN(n1629) );
  OAI21_X2 U4147 ( .B1(n2938), .B2(n2963), .A(n912), .ZN(n1630) );
  OAI21_X2 U4148 ( .B1(n2936), .B2(n2965), .A(n901), .ZN(n1631) );
  OAI21_X2 U4149 ( .B1(n2934), .B2(n2964), .A(n890), .ZN(n1632) );
  OAI21_X2 U4150 ( .B1(n2932), .B2(n2963), .A(n887), .ZN(n1633) );
  OAI21_X2 U4151 ( .B1(n2930), .B2(n2963), .A(n886), .ZN(n1634) );
  OAI21_X2 U4152 ( .B1(n2928), .B2(n2963), .A(n885), .ZN(n1635) );
  OAI21_X2 U4153 ( .B1(n2926), .B2(n2963), .A(n884), .ZN(n1636) );
  OAI21_X2 U4154 ( .B1(n2924), .B2(n2963), .A(n883), .ZN(n1637) );
  OAI21_X2 U4155 ( .B1(n2922), .B2(n2963), .A(n882), .ZN(n1638) );
  OAI21_X2 U4156 ( .B1(n2920), .B2(n2963), .A(n881), .ZN(n1639) );
  OAI21_X2 U4157 ( .B1(n2918), .B2(n2963), .A(n911), .ZN(n1640) );
  OAI21_X2 U4158 ( .B1(n2916), .B2(n2963), .A(n910), .ZN(n1641) );
  OAI21_X2 U4159 ( .B1(n2914), .B2(n2963), .A(n909), .ZN(n1642) );
  OAI21_X2 U4160 ( .B1(n2912), .B2(n2964), .A(n908), .ZN(n1643) );
  OAI21_X2 U4161 ( .B1(n2910), .B2(n2964), .A(n907), .ZN(n1644) );
  OAI21_X2 U4162 ( .B1(n2908), .B2(n2964), .A(n906), .ZN(n1645) );
  OAI21_X2 U4163 ( .B1(n2906), .B2(n2965), .A(n905), .ZN(n1646) );
  OAI21_X2 U4164 ( .B1(n2904), .B2(n2965), .A(n904), .ZN(n1647) );
  OAI21_X2 U4165 ( .B1(n2902), .B2(n2965), .A(n903), .ZN(n1648) );
  OAI21_X2 U4166 ( .B1(n2900), .B2(n2965), .A(n902), .ZN(n1649) );
  OAI21_X2 U4167 ( .B1(n2898), .B2(n2965), .A(n900), .ZN(n1650) );
  OAI21_X2 U4168 ( .B1(n2896), .B2(n2964), .A(n899), .ZN(n1651) );
  OAI21_X2 U4169 ( .B1(n2894), .B2(n2965), .A(n898), .ZN(n1652) );
  OAI21_X2 U4170 ( .B1(n2892), .B2(n2965), .A(n897), .ZN(n1653) );
  OAI21_X2 U4171 ( .B1(n2890), .B2(n2964), .A(n896), .ZN(n1654) );
  OAI21_X2 U4172 ( .B1(n2886), .B2(n2964), .A(n894), .ZN(n1656) );
  OAI21_X2 U4173 ( .B1(n2884), .B2(n2964), .A(n893), .ZN(n1657) );
  OAI21_X2 U4174 ( .B1(n2880), .B2(n2964), .A(n891), .ZN(n1659) );
  OAI21_X2 U4175 ( .B1(n2878), .B2(n2964), .A(n889), .ZN(n1660) );
  OAI21_X2 U4176 ( .B1(n2876), .B2(n2963), .A(n888), .ZN(n1661) );
  OAI21_X2 U4177 ( .B1(n2938), .B2(n2966), .A(n879), .ZN(n1662) );
  OAI21_X2 U4178 ( .B1(n2936), .B2(n2968), .A(n868), .ZN(n1663) );
  OAI21_X2 U4179 ( .B1(n2934), .B2(n2967), .A(n857), .ZN(n1664) );
  OAI21_X2 U4180 ( .B1(n2932), .B2(n2966), .A(n854), .ZN(n1665) );
  OAI21_X2 U4181 ( .B1(n2930), .B2(n2966), .A(n853), .ZN(n1666) );
  OAI21_X2 U4182 ( .B1(n2928), .B2(n2966), .A(n852), .ZN(n1667) );
  OAI21_X2 U4183 ( .B1(n2926), .B2(n2966), .A(n851), .ZN(n1668) );
  OAI21_X2 U4184 ( .B1(n2924), .B2(n2966), .A(n850), .ZN(n1669) );
  OAI21_X2 U4185 ( .B1(n2922), .B2(n2966), .A(n849), .ZN(n1670) );
  OAI21_X2 U4186 ( .B1(n2920), .B2(n2966), .A(n848), .ZN(n1671) );
  OAI21_X2 U4187 ( .B1(n2918), .B2(n2966), .A(n878), .ZN(n1672) );
  OAI21_X2 U4188 ( .B1(n2916), .B2(n2966), .A(n877), .ZN(n1673) );
  OAI21_X2 U4189 ( .B1(n2914), .B2(n2966), .A(n876), .ZN(n1674) );
  OAI21_X2 U4190 ( .B1(n2912), .B2(n2967), .A(n875), .ZN(n1675) );
  OAI21_X2 U4191 ( .B1(n2910), .B2(n2967), .A(n874), .ZN(n1676) );
  OAI21_X2 U4192 ( .B1(n2908), .B2(n2967), .A(n873), .ZN(n1677) );
  OAI21_X2 U4193 ( .B1(n2906), .B2(n2968), .A(n872), .ZN(n1678) );
  OAI21_X2 U4194 ( .B1(n2904), .B2(n2968), .A(n871), .ZN(n1679) );
  OAI21_X2 U4195 ( .B1(n2902), .B2(n2968), .A(n870), .ZN(n1680) );
  OAI21_X2 U4196 ( .B1(n2900), .B2(n2968), .A(n869), .ZN(n1681) );
  OAI21_X2 U4197 ( .B1(n2898), .B2(n2968), .A(n867), .ZN(n1682) );
  OAI21_X2 U4198 ( .B1(n2896), .B2(n2967), .A(n866), .ZN(n1683) );
  OAI21_X2 U4199 ( .B1(n2894), .B2(n2968), .A(n865), .ZN(n1684) );
  OAI21_X2 U4200 ( .B1(n2892), .B2(n2968), .A(n864), .ZN(n1685) );
  OAI21_X2 U4201 ( .B1(n2890), .B2(n2967), .A(n863), .ZN(n1686) );
  OAI21_X2 U4202 ( .B1(n2888), .B2(n2967), .A(n862), .ZN(n1687) );
  OAI21_X2 U4203 ( .B1(n2886), .B2(n2967), .A(n861), .ZN(n1688) );
  OAI21_X2 U4204 ( .B1(n2884), .B2(n2967), .A(n860), .ZN(n1689) );
  OAI21_X2 U4205 ( .B1(n2882), .B2(n2967), .A(n859), .ZN(n1690) );
  OAI21_X2 U4206 ( .B1(n2880), .B2(n2967), .A(n858), .ZN(n1691) );
  OAI21_X2 U4207 ( .B1(n2878), .B2(n2967), .A(n856), .ZN(n1692) );
  OAI21_X2 U4208 ( .B1(n2876), .B2(n2966), .A(n855), .ZN(n1693) );
  OAI21_X2 U4209 ( .B1(n2938), .B2(n2970), .A(n846), .ZN(n1694) );
  OAI21_X2 U4210 ( .B1(n2936), .B2(n2972), .A(n835), .ZN(n1695) );
  OAI21_X2 U4211 ( .B1(n2934), .B2(n2971), .A(n824), .ZN(n1696) );
  OAI21_X2 U4212 ( .B1(n2932), .B2(n2970), .A(n821), .ZN(n1697) );
  OAI21_X2 U4213 ( .B1(n2930), .B2(n2970), .A(n820), .ZN(n1698) );
  OAI21_X2 U4214 ( .B1(n2928), .B2(n2970), .A(n819), .ZN(n1699) );
  OAI21_X2 U4215 ( .B1(n2926), .B2(n2970), .A(n818), .ZN(n1700) );
  OAI21_X2 U4216 ( .B1(n2924), .B2(n2970), .A(n817), .ZN(n1701) );
  OAI21_X2 U4217 ( .B1(n2922), .B2(n2970), .A(n816), .ZN(n1702) );
  OAI21_X2 U4218 ( .B1(n2920), .B2(n2970), .A(n815), .ZN(n1703) );
  OAI21_X2 U4219 ( .B1(n2918), .B2(n2970), .A(n845), .ZN(n1704) );
  OAI21_X2 U4220 ( .B1(n2916), .B2(n2970), .A(n844), .ZN(n1705) );
  OAI21_X2 U4221 ( .B1(n2914), .B2(n2970), .A(n843), .ZN(n1706) );
  OAI21_X2 U4222 ( .B1(n2912), .B2(n2971), .A(n842), .ZN(n1707) );
  OAI21_X2 U4223 ( .B1(n2910), .B2(n2971), .A(n841), .ZN(n1708) );
  OAI21_X2 U4224 ( .B1(n2908), .B2(n2971), .A(n840), .ZN(n1709) );
  OAI21_X2 U4225 ( .B1(n2906), .B2(n2972), .A(n839), .ZN(n1710) );
  OAI21_X2 U4226 ( .B1(n2904), .B2(n2972), .A(n838), .ZN(n1711) );
  OAI21_X2 U4227 ( .B1(n2902), .B2(n2972), .A(n837), .ZN(n1712) );
  OAI21_X2 U4228 ( .B1(n2900), .B2(n2972), .A(n836), .ZN(n1713) );
  OAI21_X2 U4229 ( .B1(n2898), .B2(n2972), .A(n834), .ZN(n1714) );
  OAI21_X2 U4230 ( .B1(n2896), .B2(n2971), .A(n833), .ZN(n1715) );
  OAI21_X2 U4231 ( .B1(n2894), .B2(n2972), .A(n832), .ZN(n1716) );
  OAI21_X2 U4232 ( .B1(n2892), .B2(n2972), .A(n831), .ZN(n1717) );
  OAI21_X2 U4233 ( .B1(n2890), .B2(n2971), .A(n830), .ZN(n1718) );
  OAI21_X2 U4234 ( .B1(n2888), .B2(n2971), .A(n829), .ZN(n1719) );
  OAI21_X2 U4235 ( .B1(n2886), .B2(n2971), .A(n828), .ZN(n1720) );
  OAI21_X2 U4236 ( .B1(n2884), .B2(n2971), .A(n827), .ZN(n1721) );
  OAI21_X2 U4237 ( .B1(n2882), .B2(n2971), .A(n826), .ZN(n1722) );
  OAI21_X2 U4238 ( .B1(n2880), .B2(n2971), .A(n825), .ZN(n1723) );
  OAI21_X2 U4239 ( .B1(n2878), .B2(n2971), .A(n823), .ZN(n1724) );
  OAI21_X2 U4240 ( .B1(n2876), .B2(n2970), .A(n822), .ZN(n1725) );
  OAI21_X2 U4241 ( .B1(n2938), .B2(n2975), .A(n813), .ZN(n1726) );
  OAI21_X2 U4242 ( .B1(n2936), .B2(n2977), .A(n802), .ZN(n1727) );
  OAI21_X2 U4243 ( .B1(n2934), .B2(n2976), .A(n791), .ZN(n1728) );
  OAI21_X2 U4244 ( .B1(n2932), .B2(n2975), .A(n788), .ZN(n1729) );
  OAI21_X2 U4245 ( .B1(n2930), .B2(n2975), .A(n787), .ZN(n1730) );
  OAI21_X2 U4246 ( .B1(n2928), .B2(n2975), .A(n786), .ZN(n1731) );
  OAI21_X2 U4247 ( .B1(n2926), .B2(n2975), .A(n785), .ZN(n1732) );
  OAI21_X2 U4248 ( .B1(n2924), .B2(n2975), .A(n784), .ZN(n1733) );
  OAI21_X2 U4249 ( .B1(n2922), .B2(n2975), .A(n783), .ZN(n1734) );
  OAI21_X2 U4250 ( .B1(n2920), .B2(n2975), .A(n782), .ZN(n1735) );
  OAI21_X2 U4251 ( .B1(n2918), .B2(n2975), .A(n812), .ZN(n1736) );
  OAI21_X2 U4252 ( .B1(n2916), .B2(n2975), .A(n811), .ZN(n1737) );
  OAI21_X2 U4253 ( .B1(n2914), .B2(n2975), .A(n810), .ZN(n1738) );
  OAI21_X2 U4254 ( .B1(n2912), .B2(n2976), .A(n809), .ZN(n1739) );
  OAI21_X2 U4255 ( .B1(n2910), .B2(n2976), .A(n808), .ZN(n1740) );
  OAI21_X2 U4256 ( .B1(n2908), .B2(n2976), .A(n807), .ZN(n1741) );
  OAI21_X2 U4257 ( .B1(n2906), .B2(n2977), .A(n806), .ZN(n1742) );
  OAI21_X2 U4258 ( .B1(n2904), .B2(n2977), .A(n805), .ZN(n1743) );
  OAI21_X2 U4259 ( .B1(n2902), .B2(n2977), .A(n804), .ZN(n1744) );
  OAI21_X2 U4260 ( .B1(n2900), .B2(n2977), .A(n803), .ZN(n1745) );
  OAI21_X2 U4261 ( .B1(n2898), .B2(n2977), .A(n801), .ZN(n1746) );
  OAI21_X2 U4262 ( .B1(n2896), .B2(n2976), .A(n800), .ZN(n1747) );
  OAI21_X2 U4263 ( .B1(n2894), .B2(n2977), .A(n799), .ZN(n1748) );
  OAI21_X2 U4264 ( .B1(n2892), .B2(n2977), .A(n798), .ZN(n1749) );
  OAI21_X2 U4265 ( .B1(n2890), .B2(n2976), .A(n797), .ZN(n1750) );
  OAI21_X2 U4266 ( .B1(n2888), .B2(n2976), .A(n796), .ZN(n1751) );
  OAI21_X2 U4267 ( .B1(n2886), .B2(n2976), .A(n795), .ZN(n1752) );
  OAI21_X2 U4268 ( .B1(n2884), .B2(n2976), .A(n794), .ZN(n1753) );
  OAI21_X2 U4269 ( .B1(n2882), .B2(n2976), .A(n793), .ZN(n1754) );
  OAI21_X2 U4270 ( .B1(n2880), .B2(n2976), .A(n792), .ZN(n1755) );
  OAI21_X2 U4271 ( .B1(n2878), .B2(n2976), .A(n790), .ZN(n1756) );
  OAI21_X2 U4272 ( .B1(n2876), .B2(n2975), .A(n789), .ZN(n1757) );
  OAI21_X2 U4273 ( .B1(n2938), .B2(n2979), .A(n779), .ZN(n1758) );
  OAI21_X2 U4274 ( .B1(n2936), .B2(n2981), .A(n768), .ZN(n1759) );
  OAI21_X2 U4275 ( .B1(n2934), .B2(n2980), .A(n757), .ZN(n1760) );
  OAI21_X2 U4276 ( .B1(n2932), .B2(n2979), .A(n754), .ZN(n1761) );
  OAI21_X2 U4277 ( .B1(n2930), .B2(n2979), .A(n753), .ZN(n1762) );
  OAI21_X2 U4278 ( .B1(n2928), .B2(n2979), .A(n752), .ZN(n1763) );
  OAI21_X2 U4279 ( .B1(n2926), .B2(n2979), .A(n751), .ZN(n1764) );
  OAI21_X2 U4280 ( .B1(n2924), .B2(n2979), .A(n750), .ZN(n1765) );
  OAI21_X2 U4281 ( .B1(n2922), .B2(n2979), .A(n749), .ZN(n1766) );
  OAI21_X2 U4282 ( .B1(n2920), .B2(n2979), .A(n748), .ZN(n1767) );
  OAI21_X2 U4283 ( .B1(n2918), .B2(n2979), .A(n778), .ZN(n1768) );
  OAI21_X2 U4284 ( .B1(n2916), .B2(n2979), .A(n777), .ZN(n1769) );
  OAI21_X2 U4285 ( .B1(n2914), .B2(n2979), .A(n776), .ZN(n1770) );
  OAI21_X2 U4286 ( .B1(n2912), .B2(n2980), .A(n775), .ZN(n1771) );
  OAI21_X2 U4287 ( .B1(n2910), .B2(n2980), .A(n774), .ZN(n1772) );
  OAI21_X2 U4288 ( .B1(n2908), .B2(n2980), .A(n773), .ZN(n1773) );
  OAI21_X2 U4289 ( .B1(n2906), .B2(n2981), .A(n772), .ZN(n1774) );
  OAI21_X2 U4290 ( .B1(n2904), .B2(n2981), .A(n771), .ZN(n1775) );
  OAI21_X2 U4291 ( .B1(n2902), .B2(n2981), .A(n770), .ZN(n1776) );
  OAI21_X2 U4292 ( .B1(n2900), .B2(n2981), .A(n769), .ZN(n1777) );
  OAI21_X2 U4293 ( .B1(n2898), .B2(n2981), .A(n767), .ZN(n1778) );
  OAI21_X2 U4294 ( .B1(n2896), .B2(n2980), .A(n766), .ZN(n1779) );
  OAI21_X2 U4295 ( .B1(n2894), .B2(n2981), .A(n765), .ZN(n1780) );
  OAI21_X2 U4296 ( .B1(n2892), .B2(n2981), .A(n764), .ZN(n1781) );
  OAI21_X2 U4297 ( .B1(n2890), .B2(n2980), .A(n763), .ZN(n1782) );
  OAI21_X2 U4298 ( .B1(n2888), .B2(n2980), .A(n762), .ZN(n1783) );
  OAI21_X2 U4299 ( .B1(n2886), .B2(n2980), .A(n761), .ZN(n1784) );
  OAI21_X2 U4300 ( .B1(n2884), .B2(n2980), .A(n760), .ZN(n1785) );
  OAI21_X2 U4301 ( .B1(n2882), .B2(n2980), .A(n759), .ZN(n1786) );
  OAI21_X2 U4302 ( .B1(n2880), .B2(n2980), .A(n758), .ZN(n1787) );
  OAI21_X2 U4303 ( .B1(n2878), .B2(n2980), .A(n756), .ZN(n1788) );
  OAI21_X2 U4304 ( .B1(n2876), .B2(n2979), .A(n755), .ZN(n1789) );
  OAI21_X2 U4305 ( .B1(n2938), .B2(n2985), .A(n711), .ZN(n1790) );
  OAI21_X2 U4306 ( .B1(n2936), .B2(n2987), .A(n700), .ZN(n1791) );
  OAI21_X2 U4307 ( .B1(n2934), .B2(n2986), .A(n689), .ZN(n1792) );
  OAI21_X2 U4308 ( .B1(n2932), .B2(n2985), .A(n686), .ZN(n1793) );
  OAI21_X2 U4309 ( .B1(n2930), .B2(n2985), .A(n685), .ZN(n1794) );
  OAI21_X2 U4310 ( .B1(n2928), .B2(n2985), .A(n684), .ZN(n1795) );
  OAI21_X2 U4311 ( .B1(n2926), .B2(n2985), .A(n683), .ZN(n1796) );
  OAI21_X2 U4312 ( .B1(n2924), .B2(n2985), .A(n682), .ZN(n1797) );
  OAI21_X2 U4313 ( .B1(n2922), .B2(n2985), .A(n681), .ZN(n1798) );
  OAI21_X2 U4314 ( .B1(n2920), .B2(n2985), .A(n680), .ZN(n1799) );
  OAI21_X2 U4315 ( .B1(n2918), .B2(n2985), .A(n710), .ZN(n1800) );
  OAI21_X2 U4316 ( .B1(n2916), .B2(n2985), .A(n709), .ZN(n1801) );
  OAI21_X2 U4317 ( .B1(n2914), .B2(n2985), .A(n708), .ZN(n1802) );
  OAI21_X2 U4318 ( .B1(n2912), .B2(n2986), .A(n707), .ZN(n1803) );
  OAI21_X2 U4319 ( .B1(n2910), .B2(n2986), .A(n706), .ZN(n1804) );
  OAI21_X2 U4320 ( .B1(n2908), .B2(n2986), .A(n705), .ZN(n1805) );
  OAI21_X2 U4321 ( .B1(n2906), .B2(n2987), .A(n704), .ZN(n1806) );
  OAI21_X2 U4322 ( .B1(n2904), .B2(n2987), .A(n703), .ZN(n1807) );
  OAI21_X2 U4323 ( .B1(n2902), .B2(n2987), .A(n702), .ZN(n1808) );
  OAI21_X2 U4324 ( .B1(n2900), .B2(n2987), .A(n701), .ZN(n1809) );
  OAI21_X2 U4325 ( .B1(n2898), .B2(n2987), .A(n699), .ZN(n1810) );
  OAI21_X2 U4326 ( .B1(n2896), .B2(n2986), .A(n698), .ZN(n1811) );
  OAI21_X2 U4327 ( .B1(n2894), .B2(n2987), .A(n697), .ZN(n1812) );
  OAI21_X2 U4328 ( .B1(n2892), .B2(n2987), .A(n696), .ZN(n1813) );
  OAI21_X2 U4329 ( .B1(n2890), .B2(n2986), .A(n695), .ZN(n1814) );
  OAI21_X2 U4330 ( .B1(n2888), .B2(n2986), .A(n694), .ZN(n1815) );
  OAI21_X2 U4331 ( .B1(n2886), .B2(n2986), .A(n693), .ZN(n1816) );
  OAI21_X2 U4332 ( .B1(n2884), .B2(n2986), .A(n692), .ZN(n1817) );
  OAI21_X2 U4333 ( .B1(n2882), .B2(n2986), .A(n691), .ZN(n1818) );
  OAI21_X2 U4334 ( .B1(n2880), .B2(n2986), .A(n690), .ZN(n1819) );
  OAI21_X2 U4335 ( .B1(n2878), .B2(n2986), .A(n688), .ZN(n1820) );
  OAI21_X2 U4336 ( .B1(n2876), .B2(n2985), .A(n687), .ZN(n1821) );
  OAI21_X2 U4337 ( .B1(n2939), .B2(n2989), .A(n678), .ZN(n1822) );
  OAI21_X2 U4338 ( .B1(n2937), .B2(n2991), .A(n667), .ZN(n1823) );
  OAI21_X2 U4339 ( .B1(n2935), .B2(n2990), .A(n656), .ZN(n1824) );
  OAI21_X2 U4340 ( .B1(n2933), .B2(n2989), .A(n653), .ZN(n1825) );
  OAI21_X2 U4341 ( .B1(n2931), .B2(n2989), .A(n652), .ZN(n1826) );
  OAI21_X2 U4342 ( .B1(n2929), .B2(n2989), .A(n651), .ZN(n1827) );
  OAI21_X2 U4343 ( .B1(n2927), .B2(n2989), .A(n650), .ZN(n1828) );
  OAI21_X2 U4344 ( .B1(n2925), .B2(n2989), .A(n649), .ZN(n1829) );
  OAI21_X2 U4345 ( .B1(n2923), .B2(n2989), .A(n648), .ZN(n1830) );
  OAI21_X2 U4346 ( .B1(n2921), .B2(n2989), .A(n647), .ZN(n1831) );
  OAI21_X2 U4347 ( .B1(n2919), .B2(n2989), .A(n677), .ZN(n1832) );
  OAI21_X2 U4348 ( .B1(n2917), .B2(n2989), .A(n676), .ZN(n1833) );
  OAI21_X2 U4349 ( .B1(n2915), .B2(n2989), .A(n675), .ZN(n1834) );
  OAI21_X2 U4350 ( .B1(n2913), .B2(n2990), .A(n674), .ZN(n1835) );
  OAI21_X2 U4351 ( .B1(n2911), .B2(n2990), .A(n673), .ZN(n1836) );
  OAI21_X2 U4352 ( .B1(n2909), .B2(n2990), .A(n672), .ZN(n1837) );
  OAI21_X2 U4353 ( .B1(n2907), .B2(n2991), .A(n671), .ZN(n1838) );
  OAI21_X2 U4354 ( .B1(n2905), .B2(n2991), .A(n670), .ZN(n1839) );
  OAI21_X2 U4355 ( .B1(n2903), .B2(n2991), .A(n669), .ZN(n1840) );
  OAI21_X2 U4356 ( .B1(n2901), .B2(n2991), .A(n668), .ZN(n1841) );
  OAI21_X2 U4357 ( .B1(n2899), .B2(n2991), .A(n666), .ZN(n1842) );
  OAI21_X2 U4358 ( .B1(n2897), .B2(n2990), .A(n665), .ZN(n1843) );
  OAI21_X2 U4359 ( .B1(n2895), .B2(n2991), .A(n664), .ZN(n1844) );
  OAI21_X2 U4360 ( .B1(n2893), .B2(n2991), .A(n663), .ZN(n1845) );
  OAI21_X2 U4361 ( .B1(n2891), .B2(n2990), .A(n662), .ZN(n1846) );
  OAI21_X2 U4362 ( .B1(n2889), .B2(n2990), .A(n661), .ZN(n1847) );
  OAI21_X2 U4363 ( .B1(n2887), .B2(n2990), .A(n660), .ZN(n1848) );
  OAI21_X2 U4364 ( .B1(n2885), .B2(n2990), .A(n659), .ZN(n1849) );
  OAI21_X2 U4365 ( .B1(n2883), .B2(n2990), .A(n658), .ZN(n1850) );
  OAI21_X2 U4366 ( .B1(n2881), .B2(n2990), .A(n657), .ZN(n1851) );
  OAI21_X2 U4367 ( .B1(n2879), .B2(n2990), .A(n655), .ZN(n1852) );
  OAI21_X2 U4368 ( .B1(n2877), .B2(n2989), .A(n654), .ZN(n1853) );
  OAI21_X2 U4369 ( .B1(n2939), .B2(n2994), .A(n645), .ZN(n1854) );
  OAI21_X2 U4370 ( .B1(n2937), .B2(n2996), .A(n634), .ZN(n1855) );
  OAI21_X2 U4371 ( .B1(n2935), .B2(n2995), .A(n623), .ZN(n1856) );
  OAI21_X2 U4372 ( .B1(n2933), .B2(n2994), .A(n620), .ZN(n1857) );
  OAI21_X2 U4373 ( .B1(n2931), .B2(n2994), .A(n619), .ZN(n1858) );
  OAI21_X2 U4374 ( .B1(n2929), .B2(n2994), .A(n618), .ZN(n1859) );
  OAI21_X2 U4375 ( .B1(n2927), .B2(n2994), .A(n617), .ZN(n1860) );
  OAI21_X2 U4376 ( .B1(n2925), .B2(n2994), .A(n616), .ZN(n1861) );
  OAI21_X2 U4377 ( .B1(n2923), .B2(n2994), .A(n615), .ZN(n1862) );
  OAI21_X2 U4378 ( .B1(n2921), .B2(n2994), .A(n614), .ZN(n1863) );
  OAI21_X2 U4379 ( .B1(n2919), .B2(n2994), .A(n644), .ZN(n1864) );
  OAI21_X2 U4380 ( .B1(n2917), .B2(n2994), .A(n643), .ZN(n1865) );
  OAI21_X2 U4381 ( .B1(n2915), .B2(n2994), .A(n642), .ZN(n1866) );
  OAI21_X2 U4382 ( .B1(n2913), .B2(n2995), .A(n641), .ZN(n1867) );
  OAI21_X2 U4383 ( .B1(n2911), .B2(n2995), .A(n640), .ZN(n1868) );
  OAI21_X2 U4384 ( .B1(n2909), .B2(n2995), .A(n639), .ZN(n1869) );
  OAI21_X2 U4385 ( .B1(n2907), .B2(n2996), .A(n638), .ZN(n1870) );
  OAI21_X2 U4386 ( .B1(n2905), .B2(n2996), .A(n637), .ZN(n1871) );
  OAI21_X2 U4387 ( .B1(n2903), .B2(n2996), .A(n636), .ZN(n1872) );
  OAI21_X2 U4388 ( .B1(n2901), .B2(n2996), .A(n635), .ZN(n1873) );
  OAI21_X2 U4389 ( .B1(n2899), .B2(n2996), .A(n633), .ZN(n1874) );
  OAI21_X2 U4390 ( .B1(n2897), .B2(n2995), .A(n632), .ZN(n1875) );
  OAI21_X2 U4391 ( .B1(n2895), .B2(n2996), .A(n631), .ZN(n1876) );
  OAI21_X2 U4392 ( .B1(n2893), .B2(n2996), .A(n630), .ZN(n1877) );
  OAI21_X2 U4393 ( .B1(n2891), .B2(n2995), .A(n629), .ZN(n1878) );
  OAI21_X2 U4394 ( .B1(n2889), .B2(n2995), .A(n628), .ZN(n1879) );
  OAI21_X2 U4395 ( .B1(n2887), .B2(n2995), .A(n627), .ZN(n1880) );
  OAI21_X2 U4396 ( .B1(n2885), .B2(n2995), .A(n626), .ZN(n1881) );
  OAI21_X2 U4397 ( .B1(n2883), .B2(n2995), .A(n625), .ZN(n1882) );
  OAI21_X2 U4398 ( .B1(n2881), .B2(n2995), .A(n624), .ZN(n1883) );
  OAI21_X2 U4399 ( .B1(n2879), .B2(n2995), .A(n622), .ZN(n1884) );
  OAI21_X2 U4400 ( .B1(n2877), .B2(n2994), .A(n621), .ZN(n1885) );
  OAI21_X2 U4401 ( .B1(n2939), .B2(n2998), .A(n611), .ZN(n1886) );
  OAI21_X2 U4402 ( .B1(n2937), .B2(n3000), .A(n600), .ZN(n1887) );
  OAI21_X2 U4403 ( .B1(n2935), .B2(n2999), .A(n589), .ZN(n1888) );
  OAI21_X2 U4404 ( .B1(n2933), .B2(n2998), .A(n586), .ZN(n1889) );
  OAI21_X2 U4405 ( .B1(n2931), .B2(n2998), .A(n585), .ZN(n1890) );
  OAI21_X2 U4406 ( .B1(n2929), .B2(n2998), .A(n584), .ZN(n1891) );
  OAI21_X2 U4407 ( .B1(n2927), .B2(n2998), .A(n583), .ZN(n1892) );
  OAI21_X2 U4408 ( .B1(n2925), .B2(n2998), .A(n582), .ZN(n1893) );
  OAI21_X2 U4409 ( .B1(n2923), .B2(n2998), .A(n581), .ZN(n1894) );
  OAI21_X2 U4410 ( .B1(n2921), .B2(n2998), .A(n580), .ZN(n1895) );
  OAI21_X2 U4411 ( .B1(n2919), .B2(n2998), .A(n610), .ZN(n1896) );
  OAI21_X2 U4412 ( .B1(n2917), .B2(n2998), .A(n609), .ZN(n1897) );
  OAI21_X2 U4413 ( .B1(n2915), .B2(n2998), .A(n608), .ZN(n1898) );
  OAI21_X2 U4414 ( .B1(n2913), .B2(n2999), .A(n607), .ZN(n1899) );
  OAI21_X2 U4415 ( .B1(n2911), .B2(n2999), .A(n606), .ZN(n1900) );
  OAI21_X2 U4416 ( .B1(n2909), .B2(n2999), .A(n605), .ZN(n1901) );
  OAI21_X2 U4417 ( .B1(n2907), .B2(n3000), .A(n604), .ZN(n1902) );
  OAI21_X2 U4418 ( .B1(n2905), .B2(n3000), .A(n603), .ZN(n1903) );
  OAI21_X2 U4419 ( .B1(n2903), .B2(n3000), .A(n602), .ZN(n1904) );
  OAI21_X2 U4420 ( .B1(n2901), .B2(n3000), .A(n601), .ZN(n1905) );
  OAI21_X2 U4421 ( .B1(n2899), .B2(n3000), .A(n599), .ZN(n1906) );
  OAI21_X2 U4422 ( .B1(n2897), .B2(n2999), .A(n598), .ZN(n1907) );
  OAI21_X2 U4423 ( .B1(n2895), .B2(n3000), .A(n597), .ZN(n1908) );
  OAI21_X2 U4424 ( .B1(n2893), .B2(n3000), .A(n596), .ZN(n1909) );
  OAI21_X2 U4425 ( .B1(n2891), .B2(n2999), .A(n595), .ZN(n1910) );
  OAI21_X2 U4426 ( .B1(n2889), .B2(n2999), .A(n594), .ZN(n1911) );
  OAI21_X2 U4427 ( .B1(n2887), .B2(n2999), .A(n593), .ZN(n1912) );
  OAI21_X2 U4428 ( .B1(n2885), .B2(n2999), .A(n592), .ZN(n1913) );
  OAI21_X2 U4429 ( .B1(n2883), .B2(n2999), .A(n591), .ZN(n1914) );
  OAI21_X2 U4430 ( .B1(n2881), .B2(n2999), .A(n590), .ZN(n1915) );
  OAI21_X2 U4431 ( .B1(n2879), .B2(n2999), .A(n588), .ZN(n1916) );
  OAI21_X2 U4432 ( .B1(n2877), .B2(n2998), .A(n587), .ZN(n1917) );
  OAI21_X2 U4433 ( .B1(n2939), .B2(n3001), .A(n577), .ZN(n1918) );
  OAI21_X2 U4434 ( .B1(n2937), .B2(n3003), .A(n566), .ZN(n1919) );
  OAI21_X2 U4435 ( .B1(n2935), .B2(n3002), .A(n555), .ZN(n1920) );
  OAI21_X2 U4436 ( .B1(n2933), .B2(n3001), .A(n552), .ZN(n1921) );
  OAI21_X2 U4437 ( .B1(n2931), .B2(n3001), .A(n551), .ZN(n1922) );
  OAI21_X2 U4438 ( .B1(n2929), .B2(n3001), .A(n550), .ZN(n1923) );
  OAI21_X2 U4439 ( .B1(n2927), .B2(n3001), .A(n549), .ZN(n1924) );
  OAI21_X2 U4440 ( .B1(n2925), .B2(n3001), .A(n548), .ZN(n1925) );
  OAI21_X2 U4441 ( .B1(n2923), .B2(n3001), .A(n547), .ZN(n1926) );
  OAI21_X2 U4442 ( .B1(n2921), .B2(n3001), .A(n546), .ZN(n1927) );
  OAI21_X2 U4443 ( .B1(n2919), .B2(n3001), .A(n576), .ZN(n1928) );
  OAI21_X2 U4444 ( .B1(n2917), .B2(n3001), .A(n575), .ZN(n1929) );
  OAI21_X2 U4445 ( .B1(n2915), .B2(n3001), .A(n574), .ZN(n1930) );
  OAI21_X2 U4446 ( .B1(n2913), .B2(n3002), .A(n573), .ZN(n1931) );
  OAI21_X2 U4447 ( .B1(n2911), .B2(n3002), .A(n572), .ZN(n1932) );
  OAI21_X2 U4448 ( .B1(n2909), .B2(n3002), .A(n571), .ZN(n1933) );
  OAI21_X2 U4449 ( .B1(n2907), .B2(n3003), .A(n570), .ZN(n1934) );
  OAI21_X2 U4450 ( .B1(n2905), .B2(n3003), .A(n569), .ZN(n1935) );
  OAI21_X2 U4451 ( .B1(n2903), .B2(n3003), .A(n568), .ZN(n1936) );
  OAI21_X2 U4452 ( .B1(n2901), .B2(n3003), .A(n567), .ZN(n1937) );
  OAI21_X2 U4453 ( .B1(n2899), .B2(n3003), .A(n565), .ZN(n1938) );
  OAI21_X2 U4454 ( .B1(n2897), .B2(n3002), .A(n564), .ZN(n1939) );
  OAI21_X2 U4455 ( .B1(n2895), .B2(n3003), .A(n563), .ZN(n1940) );
  OAI21_X2 U4456 ( .B1(n2893), .B2(n3003), .A(n562), .ZN(n1941) );
  OAI21_X2 U4457 ( .B1(n2891), .B2(n3002), .A(n561), .ZN(n1942) );
  OAI21_X2 U4458 ( .B1(n2889), .B2(n3002), .A(n560), .ZN(n1943) );
  OAI21_X2 U4459 ( .B1(n2887), .B2(n3002), .A(n559), .ZN(n1944) );
  OAI21_X2 U4460 ( .B1(n2885), .B2(n3002), .A(n558), .ZN(n1945) );
  OAI21_X2 U4461 ( .B1(n2883), .B2(n3002), .A(n557), .ZN(n1946) );
  OAI21_X2 U4462 ( .B1(n2881), .B2(n3002), .A(n556), .ZN(n1947) );
  OAI21_X2 U4463 ( .B1(n2879), .B2(n3002), .A(n554), .ZN(n1948) );
  OAI21_X2 U4464 ( .B1(n2877), .B2(n3001), .A(n553), .ZN(n1949) );
  OAI21_X2 U4465 ( .B1(n2939), .B2(n3005), .A(n544), .ZN(n1950) );
  OAI21_X2 U4466 ( .B1(n2937), .B2(n3007), .A(n533), .ZN(n1951) );
  OAI21_X2 U4467 ( .B1(n2935), .B2(n3006), .A(n522), .ZN(n1952) );
  OAI21_X2 U4468 ( .B1(n2933), .B2(n3005), .A(n519), .ZN(n1953) );
  OAI21_X2 U4469 ( .B1(n2931), .B2(n3005), .A(n518), .ZN(n1954) );
  OAI21_X2 U4470 ( .B1(n2929), .B2(n3005), .A(n517), .ZN(n1955) );
  OAI21_X2 U4471 ( .B1(n2927), .B2(n3005), .A(n516), .ZN(n1956) );
  OAI21_X2 U4472 ( .B1(n2925), .B2(n3005), .A(n515), .ZN(n1957) );
  OAI21_X2 U4473 ( .B1(n2923), .B2(n3005), .A(n514), .ZN(n1958) );
  OAI21_X2 U4474 ( .B1(n2921), .B2(n3005), .A(n513), .ZN(n1959) );
  OAI21_X2 U4475 ( .B1(n2919), .B2(n3005), .A(n543), .ZN(n1960) );
  OAI21_X2 U4476 ( .B1(n2917), .B2(n3005), .A(n542), .ZN(n1961) );
  OAI21_X2 U4477 ( .B1(n2915), .B2(n3005), .A(n541), .ZN(n1962) );
  OAI21_X2 U4478 ( .B1(n2913), .B2(n3006), .A(n540), .ZN(n1963) );
  OAI21_X2 U4479 ( .B1(n2911), .B2(n3006), .A(n539), .ZN(n1964) );
  OAI21_X2 U4480 ( .B1(n2909), .B2(n3006), .A(n538), .ZN(n1965) );
  OAI21_X2 U4481 ( .B1(n2907), .B2(n3007), .A(n537), .ZN(n1966) );
  OAI21_X2 U4482 ( .B1(n2905), .B2(n3007), .A(n536), .ZN(n1967) );
  OAI21_X2 U4483 ( .B1(n2903), .B2(n3007), .A(n535), .ZN(n1968) );
  OAI21_X2 U4484 ( .B1(n2901), .B2(n3007), .A(n534), .ZN(n1969) );
  OAI21_X2 U4485 ( .B1(n2899), .B2(n3007), .A(n532), .ZN(n1970) );
  OAI21_X2 U4486 ( .B1(n2897), .B2(n3006), .A(n531), .ZN(n1971) );
  OAI21_X2 U4487 ( .B1(n2895), .B2(n3007), .A(n530), .ZN(n1972) );
  OAI21_X2 U4488 ( .B1(n2893), .B2(n3007), .A(n529), .ZN(n1973) );
  OAI21_X2 U4489 ( .B1(n2891), .B2(n3006), .A(n528), .ZN(n1974) );
  OAI21_X2 U4490 ( .B1(n2889), .B2(n3006), .A(n527), .ZN(n1975) );
  OAI21_X2 U4491 ( .B1(n2887), .B2(n3006), .A(n526), .ZN(n1976) );
  OAI21_X2 U4492 ( .B1(n2885), .B2(n3006), .A(n525), .ZN(n1977) );
  OAI21_X2 U4493 ( .B1(n2883), .B2(n3006), .A(n524), .ZN(n1978) );
  OAI21_X2 U4494 ( .B1(n2881), .B2(n3006), .A(n523), .ZN(n1979) );
  OAI21_X2 U4495 ( .B1(n2879), .B2(n3006), .A(n521), .ZN(n1980) );
  OAI21_X2 U4496 ( .B1(n2877), .B2(n3005), .A(n520), .ZN(n1981) );
  OAI21_X2 U4497 ( .B1(n2939), .B2(n3010), .A(n511), .ZN(n1982) );
  OAI21_X2 U4498 ( .B1(n2937), .B2(n3012), .A(n500), .ZN(n1983) );
  OAI21_X2 U4499 ( .B1(n2935), .B2(n3011), .A(n489), .ZN(n1984) );
  OAI21_X2 U4500 ( .B1(n2933), .B2(n3010), .A(n486), .ZN(n1985) );
  OAI21_X2 U4501 ( .B1(n2931), .B2(n3010), .A(n485), .ZN(n1986) );
  OAI21_X2 U4502 ( .B1(n2929), .B2(n3010), .A(n484), .ZN(n1987) );
  OAI21_X2 U4503 ( .B1(n2927), .B2(n3010), .A(n483), .ZN(n1988) );
  OAI21_X2 U4504 ( .B1(n2925), .B2(n3010), .A(n482), .ZN(n1989) );
  OAI21_X2 U4505 ( .B1(n2923), .B2(n3010), .A(n481), .ZN(n1990) );
  OAI21_X2 U4506 ( .B1(n2921), .B2(n3010), .A(n480), .ZN(n1991) );
  OAI21_X2 U4507 ( .B1(n2919), .B2(n3010), .A(n510), .ZN(n1992) );
  OAI21_X2 U4508 ( .B1(n2917), .B2(n3010), .A(n509), .ZN(n1993) );
  OAI21_X2 U4509 ( .B1(n2915), .B2(n3010), .A(n508), .ZN(n1994) );
  OAI21_X2 U4510 ( .B1(n2913), .B2(n3011), .A(n507), .ZN(n1995) );
  OAI21_X2 U4511 ( .B1(n2911), .B2(n3011), .A(n506), .ZN(n1996) );
  OAI21_X2 U4512 ( .B1(n2909), .B2(n3011), .A(n505), .ZN(n1997) );
  OAI21_X2 U4513 ( .B1(n2907), .B2(n3012), .A(n504), .ZN(n1998) );
  OAI21_X2 U4514 ( .B1(n2905), .B2(n3012), .A(n503), .ZN(n1999) );
  OAI21_X2 U4515 ( .B1(n2903), .B2(n3012), .A(n502), .ZN(n2000) );
  OAI21_X2 U4516 ( .B1(n2901), .B2(n3012), .A(n501), .ZN(n2001) );
  OAI21_X2 U4517 ( .B1(n2899), .B2(n3012), .A(n499), .ZN(n2002) );
  OAI21_X2 U4518 ( .B1(n2897), .B2(n3011), .A(n498), .ZN(n2003) );
  OAI21_X2 U4519 ( .B1(n2895), .B2(n3012), .A(n497), .ZN(n2004) );
  OAI21_X2 U4520 ( .B1(n2893), .B2(n3012), .A(n496), .ZN(n2005) );
  OAI21_X2 U4521 ( .B1(n2891), .B2(n3011), .A(n495), .ZN(n2006) );
  OAI21_X2 U4522 ( .B1(n2889), .B2(n3011), .A(n494), .ZN(n2007) );
  OAI21_X2 U4523 ( .B1(n2887), .B2(n3011), .A(n493), .ZN(n2008) );
  OAI21_X2 U4524 ( .B1(n2885), .B2(n3011), .A(n492), .ZN(n2009) );
  OAI21_X2 U4525 ( .B1(n2883), .B2(n3011), .A(n491), .ZN(n2010) );
  OAI21_X2 U4526 ( .B1(n2881), .B2(n3011), .A(n490), .ZN(n2011) );
  OAI21_X2 U4527 ( .B1(n2879), .B2(n3011), .A(n488), .ZN(n2012) );
  OAI21_X2 U4528 ( .B1(n2877), .B2(n3010), .A(n487), .ZN(n2013) );
  OAI21_X2 U4529 ( .B1(n2939), .B2(n3014), .A(n477), .ZN(n2014) );
  OAI21_X2 U4530 ( .B1(n2937), .B2(n3014), .A(n466), .ZN(n2015) );
  OAI21_X2 U4531 ( .B1(n2935), .B2(n3015), .A(n455), .ZN(n2016) );
  OAI21_X2 U4532 ( .B1(n2933), .B2(n3014), .A(n452), .ZN(n2017) );
  OAI21_X2 U4533 ( .B1(n2931), .B2(n3014), .A(n451), .ZN(n2018) );
  OAI21_X2 U4534 ( .B1(n2929), .B2(n3014), .A(n450), .ZN(n2019) );
  OAI21_X2 U4535 ( .B1(n2927), .B2(n3014), .A(n449), .ZN(n2020) );
  OAI21_X2 U4536 ( .B1(n2925), .B2(n3014), .A(n448), .ZN(n2021) );
  OAI21_X2 U4537 ( .B1(n2923), .B2(n3014), .A(n447), .ZN(n2022) );
  OAI21_X2 U4538 ( .B1(n2921), .B2(n3014), .A(n446), .ZN(n2023) );
  OAI21_X2 U4539 ( .B1(n2919), .B2(n3014), .A(n476), .ZN(n2024) );
  OAI21_X2 U4540 ( .B1(n2917), .B2(n3014), .A(n475), .ZN(n2025) );
  OAI21_X2 U4541 ( .B1(n2915), .B2(n3014), .A(n474), .ZN(n2026) );
  OAI21_X2 U4542 ( .B1(n2913), .B2(n3015), .A(n473), .ZN(n2027) );
  OAI21_X2 U4543 ( .B1(n2911), .B2(n3015), .A(n472), .ZN(n2028) );
  OAI21_X2 U4544 ( .B1(n2909), .B2(n3015), .A(n471), .ZN(n2029) );
  OAI21_X2 U4545 ( .B1(n2907), .B2(n445), .A(n470), .ZN(n2030) );
  OAI21_X2 U4546 ( .B1(n2905), .B2(n3015), .A(n469), .ZN(n2031) );
  OAI21_X2 U4547 ( .B1(n2903), .B2(n445), .A(n468), .ZN(n2032) );
  OAI21_X2 U4548 ( .B1(n2901), .B2(n445), .A(n467), .ZN(n2033) );
  OAI21_X2 U4549 ( .B1(n2899), .B2(n3016), .A(n465), .ZN(n2034) );
  OAI21_X2 U4550 ( .B1(n2897), .B2(n3015), .A(n464), .ZN(n2035) );
  OAI21_X2 U4551 ( .B1(n2895), .B2(n445), .A(n463), .ZN(n2036) );
  OAI21_X2 U4552 ( .B1(n2893), .B2(n445), .A(n462), .ZN(n2037) );
  OAI21_X2 U4553 ( .B1(n2891), .B2(n3015), .A(n461), .ZN(n2038) );
  OAI21_X2 U4554 ( .B1(n2889), .B2(n3015), .A(n460), .ZN(n2039) );
  OAI21_X2 U4555 ( .B1(n2887), .B2(n3015), .A(n459), .ZN(n2040) );
  OAI21_X2 U4556 ( .B1(n2885), .B2(n3015), .A(n458), .ZN(n2041) );
  OAI21_X2 U4557 ( .B1(n2883), .B2(n3015), .A(n457), .ZN(n2042) );
  OAI21_X2 U4558 ( .B1(n2881), .B2(n3015), .A(n456), .ZN(n2043) );
  OAI21_X2 U4559 ( .B1(n2879), .B2(n3015), .A(n454), .ZN(n2044) );
  OAI21_X2 U4560 ( .B1(n2877), .B2(n3014), .A(n453), .ZN(n2045) );
  OAI21_X2 U4561 ( .B1(n2939), .B2(n3018), .A(n442), .ZN(n2046) );
  OAI21_X2 U4562 ( .B1(n2937), .B2(n3020), .A(n431), .ZN(n2047) );
  OAI21_X2 U4563 ( .B1(n2935), .B2(n3019), .A(n420), .ZN(n2048) );
  OAI21_X2 U4564 ( .B1(n2933), .B2(n3018), .A(n417), .ZN(n2049) );
  OAI21_X2 U4565 ( .B1(n2931), .B2(n3018), .A(n416), .ZN(n2050) );
  OAI21_X2 U4566 ( .B1(n2929), .B2(n3018), .A(n415), .ZN(n2051) );
  OAI21_X2 U4567 ( .B1(n2927), .B2(n3018), .A(n414), .ZN(n2052) );
  OAI21_X2 U4568 ( .B1(n2925), .B2(n3018), .A(n413), .ZN(n2053) );
  OAI21_X2 U4569 ( .B1(n2923), .B2(n3018), .A(n412), .ZN(n2054) );
  OAI21_X2 U4570 ( .B1(n2921), .B2(n3018), .A(n411), .ZN(n2055) );
  OAI21_X2 U4571 ( .B1(n2919), .B2(n3018), .A(n441), .ZN(n2056) );
  OAI21_X2 U4572 ( .B1(n2917), .B2(n3018), .A(n440), .ZN(n2057) );
  OAI21_X2 U4573 ( .B1(n2915), .B2(n3018), .A(n439), .ZN(n2058) );
  OAI21_X2 U4574 ( .B1(n2913), .B2(n3019), .A(n438), .ZN(n2059) );
  OAI21_X2 U4575 ( .B1(n2911), .B2(n3019), .A(n437), .ZN(n2060) );
  OAI21_X2 U4576 ( .B1(n2909), .B2(n3019), .A(n436), .ZN(n2061) );
  OAI21_X2 U4577 ( .B1(n2907), .B2(n3020), .A(n435), .ZN(n2062) );
  OAI21_X2 U4578 ( .B1(n2905), .B2(n3020), .A(n434), .ZN(n2063) );
  OAI21_X2 U4579 ( .B1(n2903), .B2(n3020), .A(n433), .ZN(n2064) );
  OAI21_X2 U4580 ( .B1(n2901), .B2(n3020), .A(n432), .ZN(n2065) );
  OAI21_X2 U4581 ( .B1(n2899), .B2(n3020), .A(n430), .ZN(n2066) );
  OAI21_X2 U4582 ( .B1(n2897), .B2(n3019), .A(n429), .ZN(n2067) );
  OAI21_X2 U4583 ( .B1(n2895), .B2(n3020), .A(n428), .ZN(n2068) );
  OAI21_X2 U4584 ( .B1(n2893), .B2(n3020), .A(n427), .ZN(n2069) );
  OAI21_X2 U4585 ( .B1(n2891), .B2(n3019), .A(n426), .ZN(n2070) );
  OAI21_X2 U4586 ( .B1(n2889), .B2(n3019), .A(n425), .ZN(n2071) );
  OAI21_X2 U4587 ( .B1(n2887), .B2(n3019), .A(n424), .ZN(n2072) );
  OAI21_X2 U4588 ( .B1(n2885), .B2(n3019), .A(n423), .ZN(n2073) );
  OAI21_X2 U4589 ( .B1(n2883), .B2(n3019), .A(n422), .ZN(n2074) );
  OAI21_X2 U4590 ( .B1(n2881), .B2(n3019), .A(n421), .ZN(n2075) );
  OAI21_X2 U4591 ( .B1(n2879), .B2(n3019), .A(n419), .ZN(n2076) );
  OAI21_X2 U4592 ( .B1(n2877), .B2(n3018), .A(n418), .ZN(n2077) );
  OAI21_X2 U4593 ( .B1(n2939), .B2(n3021), .A(n409), .ZN(n2078) );
  OAI21_X2 U4594 ( .B1(n2937), .B2(n3023), .A(n398), .ZN(n2079) );
  OAI21_X2 U4595 ( .B1(n2935), .B2(n3022), .A(n387), .ZN(n2080) );
  OAI21_X2 U4596 ( .B1(n2933), .B2(n3021), .A(n384), .ZN(n2081) );
  OAI21_X2 U4597 ( .B1(n2931), .B2(n3021), .A(n383), .ZN(n2082) );
  OAI21_X2 U4598 ( .B1(n2929), .B2(n3021), .A(n382), .ZN(n2083) );
  OAI21_X2 U4599 ( .B1(n2927), .B2(n3021), .A(n381), .ZN(n2084) );
  OAI21_X2 U4600 ( .B1(n2925), .B2(n3021), .A(n380), .ZN(n2085) );
  OAI21_X2 U4601 ( .B1(n2923), .B2(n3021), .A(n379), .ZN(n2086) );
  OAI21_X2 U4602 ( .B1(n2921), .B2(n3021), .A(n378), .ZN(n2087) );
  OAI21_X2 U4603 ( .B1(n2919), .B2(n3021), .A(n408), .ZN(n2088) );
  OAI21_X2 U4604 ( .B1(n2917), .B2(n3021), .A(n407), .ZN(n2089) );
  OAI21_X2 U4605 ( .B1(n2915), .B2(n3021), .A(n406), .ZN(n2090) );
  OAI21_X2 U4606 ( .B1(n2913), .B2(n3022), .A(n405), .ZN(n2091) );
  OAI21_X2 U4607 ( .B1(n2911), .B2(n3022), .A(n404), .ZN(n2092) );
  OAI21_X2 U4608 ( .B1(n2909), .B2(n3022), .A(n403), .ZN(n2093) );
  OAI21_X2 U4609 ( .B1(n2907), .B2(n3023), .A(n402), .ZN(n2094) );
  OAI21_X2 U4610 ( .B1(n2905), .B2(n3023), .A(n401), .ZN(n2095) );
  OAI21_X2 U4611 ( .B1(n2903), .B2(n3023), .A(n400), .ZN(n2096) );
  OAI21_X2 U4612 ( .B1(n2901), .B2(n3023), .A(n399), .ZN(n2097) );
  OAI21_X2 U4613 ( .B1(n2899), .B2(n3023), .A(n397), .ZN(n2098) );
  OAI21_X2 U4614 ( .B1(n2897), .B2(n3022), .A(n396), .ZN(n2099) );
  OAI21_X2 U4615 ( .B1(n2895), .B2(n3023), .A(n395), .ZN(n2100) );
  OAI21_X2 U4616 ( .B1(n2893), .B2(n3023), .A(n394), .ZN(n2101) );
  OAI21_X2 U4617 ( .B1(n2891), .B2(n3022), .A(n393), .ZN(n2102) );
  OAI21_X2 U4618 ( .B1(n2889), .B2(n3022), .A(n392), .ZN(n2103) );
  OAI21_X2 U4619 ( .B1(n2887), .B2(n3022), .A(n391), .ZN(n2104) );
  OAI21_X2 U4620 ( .B1(n2885), .B2(n3022), .A(n390), .ZN(n2105) );
  OAI21_X2 U4621 ( .B1(n2883), .B2(n3022), .A(n389), .ZN(n2106) );
  OAI21_X2 U4622 ( .B1(n2881), .B2(n3022), .A(n388), .ZN(n2107) );
  OAI21_X2 U4623 ( .B1(n2879), .B2(n3022), .A(n386), .ZN(n2108) );
  OAI21_X2 U4624 ( .B1(n2877), .B2(n3021), .A(n385), .ZN(n2109) );
  OAI21_X2 U4625 ( .B1(n2939), .B2(n3029), .A(n343), .ZN(n2110) );
  OAI21_X2 U4626 ( .B1(n2937), .B2(n3031), .A(n332), .ZN(n2111) );
  OAI21_X2 U4627 ( .B1(n2935), .B2(n3030), .A(n321), .ZN(n2112) );
  OAI21_X2 U4628 ( .B1(n2933), .B2(n3029), .A(n318), .ZN(n2113) );
  OAI21_X2 U4629 ( .B1(n2931), .B2(n3029), .A(n317), .ZN(n2114) );
  OAI21_X2 U4630 ( .B1(n2929), .B2(n3029), .A(n316), .ZN(n2115) );
  OAI21_X2 U4631 ( .B1(n2927), .B2(n3029), .A(n315), .ZN(n2116) );
  OAI21_X2 U4632 ( .B1(n2925), .B2(n3029), .A(n314), .ZN(n2117) );
  OAI21_X2 U4633 ( .B1(n2923), .B2(n3029), .A(n313), .ZN(n2118) );
  OAI21_X2 U4634 ( .B1(n2921), .B2(n3029), .A(n312), .ZN(n2119) );
  OAI21_X2 U4635 ( .B1(n2919), .B2(n3029), .A(n342), .ZN(n2120) );
  OAI21_X2 U4636 ( .B1(n2917), .B2(n3029), .A(n341), .ZN(n2121) );
  OAI21_X2 U4637 ( .B1(n2915), .B2(n3029), .A(n340), .ZN(n2122) );
  OAI21_X2 U4638 ( .B1(n2913), .B2(n3030), .A(n339), .ZN(n2123) );
  OAI21_X2 U4639 ( .B1(n2911), .B2(n3030), .A(n338), .ZN(n2124) );
  OAI21_X2 U4640 ( .B1(n2909), .B2(n3030), .A(n337), .ZN(n2125) );
  OAI21_X2 U4641 ( .B1(n2907), .B2(n3031), .A(n336), .ZN(n2126) );
  OAI21_X2 U4642 ( .B1(n2905), .B2(n3031), .A(n335), .ZN(n2127) );
  OAI21_X2 U4643 ( .B1(n2903), .B2(n3031), .A(n334), .ZN(n2128) );
  OAI21_X2 U4644 ( .B1(n2901), .B2(n3031), .A(n333), .ZN(n2129) );
  OAI21_X2 U4645 ( .B1(n2899), .B2(n3031), .A(n331), .ZN(n2130) );
  OAI21_X2 U4646 ( .B1(n2897), .B2(n3030), .A(n330), .ZN(n2131) );
  OAI21_X2 U4647 ( .B1(n2895), .B2(n3031), .A(n329), .ZN(n2132) );
  OAI21_X2 U4648 ( .B1(n2893), .B2(n3031), .A(n328), .ZN(n2133) );
  OAI21_X2 U4649 ( .B1(n2891), .B2(n3030), .A(n327), .ZN(n2134) );
  OAI21_X2 U4650 ( .B1(n2889), .B2(n3030), .A(n326), .ZN(n2135) );
  OAI21_X2 U4651 ( .B1(n2887), .B2(n3030), .A(n325), .ZN(n2136) );
  OAI21_X2 U4652 ( .B1(n2885), .B2(n3030), .A(n324), .ZN(n2137) );
  OAI21_X2 U4653 ( .B1(n2883), .B2(n3030), .A(n323), .ZN(n2138) );
  OAI21_X2 U4654 ( .B1(n2881), .B2(n3030), .A(n322), .ZN(n2139) );
  OAI21_X2 U4655 ( .B1(n2879), .B2(n3030), .A(n320), .ZN(n2140) );
  OAI21_X2 U4656 ( .B1(n2877), .B2(n3029), .A(n319), .ZN(n2141) );
  OAI21_X2 U4657 ( .B1(n2939), .B2(n3033), .A(n309), .ZN(n2142) );
  OAI21_X2 U4658 ( .B1(n2937), .B2(n3035), .A(n298), .ZN(n2143) );
  OAI21_X2 U4659 ( .B1(n2935), .B2(n3034), .A(n287), .ZN(n2144) );
  OAI21_X2 U4660 ( .B1(n2933), .B2(n3033), .A(n284), .ZN(n2145) );
  OAI21_X2 U4661 ( .B1(n2931), .B2(n3033), .A(n283), .ZN(n2146) );
  OAI21_X2 U4662 ( .B1(n2929), .B2(n3033), .A(n282), .ZN(n2147) );
  OAI21_X2 U4663 ( .B1(n2927), .B2(n3033), .A(n281), .ZN(n2148) );
  OAI21_X2 U4664 ( .B1(n2925), .B2(n3033), .A(n280), .ZN(n2149) );
  OAI21_X2 U4665 ( .B1(n2923), .B2(n3033), .A(n279), .ZN(n2150) );
  OAI21_X2 U4666 ( .B1(n2921), .B2(n3033), .A(n278), .ZN(n2151) );
  OAI21_X2 U4667 ( .B1(n2919), .B2(n3033), .A(n308), .ZN(n2152) );
  OAI21_X2 U4668 ( .B1(n2917), .B2(n3033), .A(n307), .ZN(n2153) );
  OAI21_X2 U4669 ( .B1(n2915), .B2(n3033), .A(n306), .ZN(n2154) );
  OAI21_X2 U4670 ( .B1(n2913), .B2(n3034), .A(n305), .ZN(n2155) );
  OAI21_X2 U4671 ( .B1(n2911), .B2(n3034), .A(n304), .ZN(n2156) );
  OAI21_X2 U4672 ( .B1(n2909), .B2(n3034), .A(n303), .ZN(n2157) );
  OAI21_X2 U4673 ( .B1(n2907), .B2(n3035), .A(n302), .ZN(n2158) );
  OAI21_X2 U4674 ( .B1(n2905), .B2(n3035), .A(n301), .ZN(n2159) );
  OAI21_X2 U4675 ( .B1(n2903), .B2(n3035), .A(n300), .ZN(n2160) );
  OAI21_X2 U4676 ( .B1(n2901), .B2(n3035), .A(n299), .ZN(n2161) );
  OAI21_X2 U4677 ( .B1(n2899), .B2(n3035), .A(n297), .ZN(n2162) );
  OAI21_X2 U4678 ( .B1(n2897), .B2(n3034), .A(n296), .ZN(n2163) );
  OAI21_X2 U4679 ( .B1(n2895), .B2(n3035), .A(n295), .ZN(n2164) );
  OAI21_X2 U4680 ( .B1(n2893), .B2(n3035), .A(n294), .ZN(n2165) );
  OAI21_X2 U4681 ( .B1(n2891), .B2(n3034), .A(n293), .ZN(n2166) );
  OAI21_X2 U4682 ( .B1(n2889), .B2(n3034), .A(n292), .ZN(n2167) );
  OAI21_X2 U4683 ( .B1(n2887), .B2(n3034), .A(n291), .ZN(n2168) );
  OAI21_X2 U4684 ( .B1(n2885), .B2(n3034), .A(n290), .ZN(n2169) );
  OAI21_X2 U4685 ( .B1(n2883), .B2(n3034), .A(n289), .ZN(n2170) );
  OAI21_X2 U4686 ( .B1(n2881), .B2(n3034), .A(n288), .ZN(n2171) );
  OAI21_X2 U4687 ( .B1(n2879), .B2(n3034), .A(n286), .ZN(n2172) );
  OAI21_X2 U4688 ( .B1(n2877), .B2(n3033), .A(n285), .ZN(n2173) );
  OAI21_X2 U4689 ( .B1(n3259), .B2(n3258), .A(n3257), .ZN(N194) );
  AOI211_X2 U4690 ( .C1(n3216), .C2(n3215), .A(n2556), .B(n2435), .ZN(n3229)
         );
  OAI21_X2 U4691 ( .B1(n3700), .B2(n3699), .A(n3698), .ZN(N205) );
  OAI21_X2 U4692 ( .B1(n4107), .B2(n4106), .A(n4105), .ZN(N215) );
  OAI21_X2 U4693 ( .B1(n5211), .B2(n5210), .A(n5209), .ZN(n5212) );
  OAI21_X2 U4694 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5794) );
  OAI21_X2 U4695 ( .B1(n2888), .B2(n2964), .A(n895), .ZN(n1655) );
  INV_X4 U4696 ( .A(n2324), .ZN(n2325) );
  NOR2_X2 U4697 ( .A1(n2325), .A2(n2803), .ZN(n4439) );
  OAI21_X2 U4698 ( .B1(n2882), .B2(n2964), .A(n892), .ZN(n1658) );
  NAND2_X4 U4699 ( .A1(n4383), .A2(n4382), .ZN(n4386) );
  NAND2_X4 U4700 ( .A1(n4444), .A2(n3161), .ZN(n4445) );
  NOR2_X2 U4701 ( .A1(n2762), .A2(n4250), .ZN(n4251) );
  NAND2_X4 U4702 ( .A1(n4126), .A2(n4125), .ZN(n4135) );
  NAND2_X4 U4703 ( .A1(n4504), .A2(n4503), .ZN(n4513) );
  NAND2_X4 U4704 ( .A1(n4446), .A2(n4445), .ZN(n4449) );
  NAND2_X4 U4705 ( .A1(n4257), .A2(n4256), .ZN(n4260) );
  NAND2_X4 U4706 ( .A1(n4320), .A2(n4319), .ZN(n4323) );
  INV_X4 U4707 ( .A(n2847), .ZN(n2327) );
  INV_X4 U4708 ( .A(n2847), .ZN(n2328) );
  INV_X4 U4709 ( .A(n2847), .ZN(n2329) );
  INV_X4 U4710 ( .A(n2847), .ZN(n2330) );
  INV_X4 U4711 ( .A(n2842), .ZN(n2331) );
  INV_X4 U4712 ( .A(n2842), .ZN(n2332) );
  INV_X4 U4713 ( .A(n2842), .ZN(n2333) );
  INV_X4 U4714 ( .A(n2842), .ZN(n2334) );
  INV_X4 U4715 ( .A(n2844), .ZN(n2335) );
  INV_X4 U4716 ( .A(n2844), .ZN(n2336) );
  INV_X4 U4717 ( .A(n2844), .ZN(n2337) );
  INV_X4 U4718 ( .A(n2844), .ZN(n2338) );
  INV_X2 U4719 ( .A(n2845), .ZN(n2340) );
  INV_X4 U4720 ( .A(n2845), .ZN(n2341) );
  INV_X4 U4721 ( .A(n2845), .ZN(n2342) );
  INV_X2 U4722 ( .A(n5737), .ZN(n2347) );
  NAND2_X4 U4723 ( .A1(n4684), .A2(n2365), .ZN(n5737) );
  INV_X4 U4724 ( .A(n2844), .ZN(n2841) );
  INV_X4 U4725 ( .A(n2846), .ZN(n2845) );
  NOR3_X1 U4726 ( .A1(n3214), .A2(n2761), .A3(n3213), .ZN(n3215) );
  NOR3_X1 U4727 ( .A1(n3225), .A2(n2761), .A3(n3224), .ZN(n3226) );
  NOR2_X2 U4728 ( .A1(n2761), .A2(n4362), .ZN(n4363) );
  NOR2_X2 U4729 ( .A1(n2761), .A2(n4299), .ZN(n4300) );
  NOR2_X2 U4730 ( .A1(n2761), .A2(n4425), .ZN(n4426) );
  NOR2_X2 U4731 ( .A1(n2761), .A2(n4614), .ZN(n4615) );
  NOR2_X2 U4732 ( .A1(n2761), .A2(n4551), .ZN(n4552) );
  NOR2_X2 U4733 ( .A1(n2761), .A2(n4392), .ZN(n4393) );
  NOR2_X2 U4734 ( .A1(n2761), .A2(n4518), .ZN(n4519) );
  NOR2_X2 U4735 ( .A1(n2761), .A2(n4644), .ZN(n4645) );
  NOR2_X2 U4736 ( .A1(n2761), .A2(n4581), .ZN(n4582) );
  NOR2_X2 U4737 ( .A1(n2761), .A2(n4376), .ZN(n4377) );
  NOR2_X2 U4738 ( .A1(n2761), .A2(n4628), .ZN(n4629) );
  NOR2_X2 U4739 ( .A1(n2761), .A2(n4439), .ZN(n4440) );
  NOR2_X2 U4740 ( .A1(n2761), .A2(n4313), .ZN(n4314) );
  NOR2_X2 U4741 ( .A1(n2761), .A2(n4565), .ZN(n4566) );
  NOR2_X2 U4742 ( .A1(n2761), .A2(n4343), .ZN(n4344) );
  NOR2_X2 U4743 ( .A1(n2761), .A2(n4329), .ZN(n4330) );
  NOR2_X2 U4744 ( .A1(n2761), .A2(n4661), .ZN(n4662) );
  NOR2_X2 U4745 ( .A1(n2761), .A2(n4532), .ZN(n4533) );
  NOR2_X2 U4746 ( .A1(n2761), .A2(n4595), .ZN(n4596) );
  NOR3_X1 U4747 ( .A1(n3087), .A2(n3065), .A3(mem_2__29_), .ZN(n6038) );
  NOR3_X2 U4748 ( .A1(n3088), .A2(n3065), .A3(mem_2__23_), .ZN(n5797) );
  NOR3_X2 U4749 ( .A1(n3087), .A2(n3065), .A3(mem_2__25_), .ZN(n5878) );
  NOR3_X2 U4750 ( .A1(n3087), .A2(n3065), .A3(mem_2__27_), .ZN(n5958) );
  NOR3_X2 U4751 ( .A1(n3087), .A2(n3065), .A3(mem_2__26_), .ZN(n5918) );
  NOR3_X2 U4752 ( .A1(n3087), .A2(n3065), .A3(mem_18__26_), .ZN(n5936) );
  NOR3_X2 U4753 ( .A1(n3087), .A2(n3065), .A3(mem_18__25_), .ZN(n5896) );
  NOR3_X2 U4754 ( .A1(n3088), .A2(n3065), .A3(mem_26__25_), .ZN(n5904) );
  NOR3_X2 U4755 ( .A1(n3087), .A2(n3065), .A3(mem_26__26_), .ZN(n5944) );
  NAND3_X1 U4756 ( .A1(n2267), .A2(mem_0__30_), .A3(n3147), .ZN(n4560) );
  NAND3_X2 U4757 ( .A1(n2249), .A2(mem_0__31_), .A3(n3147), .ZN(n4623) );
  NAND3_X2 U4758 ( .A1(n2772), .A2(mem_1__30_), .A3(n3147), .ZN(n4559) );
  NAND3_X2 U4759 ( .A1(n2772), .A2(mem_1__31_), .A3(n3147), .ZN(n4622) );
  NAND3_X2 U4760 ( .A1(n2256), .A2(mem_16__30_), .A3(n3147), .ZN(n4590) );
  NAND3_X2 U4761 ( .A1(n2772), .A2(mem_17__30_), .A3(n3147), .ZN(n4589) );
  NAND3_X2 U4762 ( .A1(n2254), .A2(mem_8__30_), .A3(n3147), .ZN(n4574) );
  NAND3_X2 U4763 ( .A1(n2772), .A2(mem_9__30_), .A3(n3147), .ZN(n4573) );
  NAND3_X2 U4764 ( .A1(n2292), .A2(mem_24__29_), .A3(n3147), .ZN(n4541) );
  NAND3_X2 U4765 ( .A1(n2291), .A2(mem_24__30_), .A3(n3147), .ZN(n4604) );
  NAND3_X2 U4766 ( .A1(n2771), .A2(mem_25__29_), .A3(n3147), .ZN(n4540) );
  NAND3_X2 U4767 ( .A1(n2771), .A2(mem_25__30_), .A3(n3147), .ZN(n4603) );
  INV_X16 U4768 ( .A(n3122), .ZN(n3144) );
  INV_X4 U4769 ( .A(n4097), .ZN(n2348) );
  INV_X4 U4770 ( .A(n4097), .ZN(n2349) );
  INV_X4 U4771 ( .A(n4097), .ZN(n2350) );
  INV_X2 U4772 ( .A(n4097), .ZN(n2351) );
  INV_X4 U4773 ( .A(n2348), .ZN(n2352) );
  INV_X4 U4774 ( .A(n2348), .ZN(n2353) );
  INV_X4 U4775 ( .A(n2348), .ZN(n2354) );
  INV_X4 U4776 ( .A(n2348), .ZN(n2355) );
  INV_X2 U4777 ( .A(n2348), .ZN(n2356) );
  INV_X8 U4778 ( .A(n2786), .ZN(n2785) );
  INV_X16 U4779 ( .A(n2872), .ZN(n2870) );
  AND2_X4 U4780 ( .A1(n139), .A2(n140), .ZN(n2357) );
  AND2_X4 U4781 ( .A1(n174), .A2(n140), .ZN(n2358) );
  AND2_X4 U4782 ( .A1(n276), .A2(n174), .ZN(n2359) );
  AND2_X4 U4783 ( .A1(n276), .A2(n139), .ZN(n2360) );
  AND2_X4 U4784 ( .A1(n140), .A2(n105), .ZN(n2361) );
  AND2_X4 U4785 ( .A1(n140), .A2(n70), .ZN(n2362) );
  AND2_X4 U4786 ( .A1(n276), .A2(n70), .ZN(n2363) );
  INV_X4 U4787 ( .A(n4664), .ZN(n2829) );
  INV_X4 U4788 ( .A(n2841), .ZN(n2843) );
  INV_X4 U4789 ( .A(n3122), .ZN(n3143) );
  INV_X4 U4790 ( .A(n3136), .ZN(n3121) );
  INV_X4 U4791 ( .A(n3121), .ZN(n3147) );
  INV_X4 U4792 ( .A(n4665), .ZN(n2831) );
  INV_X16 U4793 ( .A(n2839), .ZN(n2836) );
  INV_X16 U4794 ( .A(n2839), .ZN(n2837) );
  INV_X16 U4795 ( .A(n2839), .ZN(n2838) );
  INV_X8 U4796 ( .A(n3161), .ZN(n3157) );
  AND2_X4 U4797 ( .A1(n3064), .A2(n3072), .ZN(n2364) );
  INV_X4 U4798 ( .A(n2363), .ZN(n2984) );
  INV_X4 U4799 ( .A(n2361), .ZN(n3041) );
  INV_X4 U4800 ( .A(n2362), .ZN(n3044) );
  INV_X4 U4801 ( .A(n2358), .ZN(n3047) );
  INV_X4 U4802 ( .A(n2357), .ZN(n3050) );
  INV_X4 U4803 ( .A(n2359), .ZN(n3027) );
  INV_X4 U4804 ( .A(n2360), .ZN(n3038) );
  INV_X4 U4805 ( .A(n2788), .ZN(n2787) );
  AND2_X4 U4806 ( .A1(n2505), .A2(n2381), .ZN(n2365) );
  INV_X4 U4807 ( .A(n2765), .ZN(n2764) );
  INV_X4 U4808 ( .A(n4050), .ZN(n2765) );
  INV_X8 U4809 ( .A(n2763), .ZN(n2761) );
  INV_X4 U4810 ( .A(n3122), .ZN(n3145) );
  INV_X1 U4811 ( .A(n3136), .ZN(n3120) );
  INV_X4 U4812 ( .A(n3120), .ZN(n3148) );
  INV_X4 U4813 ( .A(n3120), .ZN(n3149) );
  INV_X4 U4814 ( .A(n3109), .ZN(n3098) );
  INV_X8 U4815 ( .A(n3110), .ZN(n3101) );
  INV_X16 U4816 ( .A(n2840), .ZN(n2834) );
  INV_X4 U4817 ( .A(n3084), .ZN(n3077) );
  INV_X4 U4818 ( .A(n3084), .ZN(n3079) );
  INV_X4 U4819 ( .A(n3084), .ZN(n3080) );
  INV_X8 U4820 ( .A(n3162), .ZN(n3156) );
  INV_X16 U4821 ( .A(n2872), .ZN(n2871) );
  INV_X16 U4822 ( .A(n2872), .ZN(n2869) );
  INV_X4 U4823 ( .A(n2371), .ZN(n2855) );
  INV_X4 U4824 ( .A(n2846), .ZN(n2844) );
  INV_X4 U4825 ( .A(n2785), .ZN(n2773) );
  INV_X8 U4826 ( .A(n2786), .ZN(n2784) );
  INV_X8 U4827 ( .A(rs2[2]), .ZN(n3137) );
  AND2_X4 U4828 ( .A1(n3067), .A2(n3064), .ZN(n2366) );
  AND2_X4 U4829 ( .A1(n3071), .A2(n3062), .ZN(n2367) );
  AND2_X4 U4830 ( .A1(n2364), .A2(n3062), .ZN(n2368) );
  AND2_X4 U4831 ( .A1(n2366), .A2(n3062), .ZN(n2369) );
  INV_X4 U4832 ( .A(n3064), .ZN(n3063) );
  INV_X8 U4833 ( .A(rs1[0]), .ZN(n3107) );
  INV_X4 U4834 ( .A(n3109), .ZN(n3099) );
  INV_X4 U4835 ( .A(n3110), .ZN(n3102) );
  INV_X8 U4836 ( .A(n3163), .ZN(n3159) );
  INV_X8 U4837 ( .A(n2801), .ZN(n2811) );
  INV_X16 U4838 ( .A(n2811), .ZN(n2806) );
  AND2_X4 U4839 ( .A1(n3150), .A2(n3118), .ZN(n2370) );
  NAND2_X2 U4840 ( .A1(n3109), .A2(n3083), .ZN(n2371) );
  INV_X4 U4841 ( .A(rs1[1]), .ZN(n3083) );
  INV_X4 U4842 ( .A(n3084), .ZN(n3078) );
  AND3_X4 U4843 ( .A1(mem_1__2_), .A2(n2768), .A3(n3148), .ZN(n2372) );
  AND2_X4 U4844 ( .A1(n2352), .A2(n3118), .ZN(n2373) );
  INV_X16 U4845 ( .A(n2830), .ZN(n2840) );
  INV_X8 U4846 ( .A(n2773), .ZN(n2769) );
  INV_X4 U4847 ( .A(n2774), .ZN(n2766) );
  INV_X4 U4848 ( .A(n3066), .ZN(n3070) );
  INV_X4 U4849 ( .A(n3065), .ZN(n3071) );
  INV_X4 U4850 ( .A(n3137), .ZN(n3119) );
  INV_X4 U4851 ( .A(n3124), .ZN(n3150) );
  INV_X4 U4852 ( .A(n3119), .ZN(n3153) );
  AND2_X2 U4853 ( .A1(n3063), .A2(n3067), .ZN(n2374) );
  INV_X4 U4854 ( .A(n3112), .ZN(n3111) );
  AND2_X4 U4855 ( .A1(n3104), .A2(n3069), .ZN(n2375) );
  AND2_X2 U4856 ( .A1(n3134), .A2(n3118), .ZN(n2376) );
  AND3_X4 U4857 ( .A1(n6162), .A2(n6161), .A3(n6160), .ZN(n2377) );
  AND2_X4 U4858 ( .A1(n3085), .A2(n3069), .ZN(n2378) );
  AND4_X4 U4859 ( .A1(n746), .A2(n105), .A3(regWr), .A4(n7227), .ZN(n2379) );
  INV_X4 U4860 ( .A(n3066), .ZN(n3073) );
  INV_X4 U4861 ( .A(rs1[2]), .ZN(n3072) );
  NAND3_X2 U4862 ( .A1(n3206), .A2(n2377), .A3(n3205), .ZN(n4097) );
  AND2_X2 U4863 ( .A1(n3134), .A2(n3112), .ZN(n2380) );
  XNOR2_X2 U4864 ( .A(rs1[4]), .B(rd[4]), .ZN(n2381) );
  AND2_X2 U4865 ( .A1(n3075), .A2(n3064), .ZN(n2382) );
  AND3_X4 U4866 ( .A1(mem_1__23_), .A2(n2866), .A3(n3073), .ZN(n2383) );
  AND3_X4 U4867 ( .A1(mem_9__23_), .A2(n2866), .A3(n3073), .ZN(n2384) );
  AND3_X4 U4868 ( .A1(mem_17__23_), .A2(n2866), .A3(n3073), .ZN(n2385) );
  AND3_X4 U4869 ( .A1(mem_1__24_), .A2(n2866), .A3(n3073), .ZN(n2386) );
  AND3_X4 U4870 ( .A1(mem_9__24_), .A2(n2866), .A3(n3073), .ZN(n2387) );
  AND3_X4 U4871 ( .A1(mem_17__24_), .A2(n2866), .A3(n3072), .ZN(n2388) );
  AND3_X4 U4872 ( .A1(mem_25__24_), .A2(n2866), .A3(n3072), .ZN(n2389) );
  AND3_X4 U4873 ( .A1(mem_1__25_), .A2(n2866), .A3(n3072), .ZN(n2390) );
  AND3_X4 U4874 ( .A1(mem_9__25_), .A2(n2866), .A3(n3072), .ZN(n2391) );
  AND3_X4 U4875 ( .A1(mem_17__25_), .A2(n2866), .A3(n3072), .ZN(n2392) );
  AND3_X4 U4876 ( .A1(mem_25__25_), .A2(n2867), .A3(n3072), .ZN(n2393) );
  AND3_X4 U4877 ( .A1(mem_1__26_), .A2(n2867), .A3(n3072), .ZN(n2394) );
  AND3_X4 U4878 ( .A1(mem_9__26_), .A2(n2867), .A3(n3073), .ZN(n2395) );
  AND3_X4 U4879 ( .A1(mem_17__26_), .A2(n2867), .A3(n3072), .ZN(n2396) );
  AND3_X4 U4880 ( .A1(mem_25__26_), .A2(n2867), .A3(n3073), .ZN(n2397) );
  AND3_X4 U4881 ( .A1(mem_1__27_), .A2(n2867), .A3(n3073), .ZN(n2398) );
  AND3_X4 U4882 ( .A1(mem_9__27_), .A2(n2867), .A3(n3072), .ZN(n2399) );
  AND3_X4 U4883 ( .A1(mem_17__27_), .A2(n2867), .A3(n3071), .ZN(n2400) );
  AND3_X4 U4884 ( .A1(mem_25__27_), .A2(n2867), .A3(n3071), .ZN(n2401) );
  AND3_X4 U4885 ( .A1(mem_1__28_), .A2(n2867), .A3(n3071), .ZN(n2402) );
  AND3_X4 U4886 ( .A1(mem_9__28_), .A2(n2867), .A3(n3071), .ZN(n2403) );
  AND3_X4 U4887 ( .A1(mem_17__28_), .A2(n2867), .A3(n3071), .ZN(n2404) );
  AND3_X4 U4888 ( .A1(mem_25__28_), .A2(n2868), .A3(n3071), .ZN(n2405) );
  AND3_X4 U4889 ( .A1(mem_1__29_), .A2(n2868), .A3(n3070), .ZN(n2406) );
  AND3_X4 U4890 ( .A1(mem_9__29_), .A2(n2868), .A3(n3070), .ZN(n2407) );
  AND3_X4 U4891 ( .A1(mem_17__29_), .A2(n2868), .A3(n3070), .ZN(n2408) );
  AND3_X4 U4892 ( .A1(mem_25__29_), .A2(n2868), .A3(n3070), .ZN(n2409) );
  AND3_X4 U4893 ( .A1(mem_1__30_), .A2(n2868), .A3(n3070), .ZN(n2410) );
  AND3_X4 U4894 ( .A1(mem_9__30_), .A2(n2868), .A3(n3070), .ZN(n2411) );
  AND3_X4 U4895 ( .A1(mem_17__30_), .A2(n2868), .A3(n3070), .ZN(n2412) );
  AND3_X4 U4896 ( .A1(mem_25__30_), .A2(n2868), .A3(n3070), .ZN(n2413) );
  AND3_X4 U4897 ( .A1(mem_1__31_), .A2(n2868), .A3(n3070), .ZN(n2414) );
  AND3_X4 U4898 ( .A1(mem_9__31_), .A2(n2868), .A3(n3071), .ZN(n2415) );
  AND3_X4 U4899 ( .A1(mem_17__31_), .A2(n2868), .A3(n3071), .ZN(n2416) );
  AND3_X4 U4900 ( .A1(mem_25__31_), .A2(n2867), .A3(n3071), .ZN(n2417) );
  AND2_X2 U4901 ( .A1(n2621), .A2(n3134), .ZN(n2418) );
  AND3_X4 U4902 ( .A1(mem_17__15_), .A2(n2769), .A3(n3138), .ZN(n2419) );
  AND3_X4 U4903 ( .A1(mem_25__15_), .A2(n2769), .A3(n3138), .ZN(n2420) );
  AND3_X4 U4904 ( .A1(mem_1__16_), .A2(n2768), .A3(n3138), .ZN(n2421) );
  AND3_X4 U4905 ( .A1(mem_9__16_), .A2(n2784), .A3(n3138), .ZN(n2422) );
  AND3_X4 U4906 ( .A1(mem_17__16_), .A2(n2784), .A3(n3138), .ZN(n2423) );
  AND3_X4 U4907 ( .A1(mem_25__16_), .A2(n2784), .A3(n3138), .ZN(n2424) );
  AND3_X4 U4908 ( .A1(mem_1__17_), .A2(n2784), .A3(n3139), .ZN(n2425) );
  AND3_X4 U4909 ( .A1(mem_9__17_), .A2(n2784), .A3(n3139), .ZN(n2426) );
  AND3_X4 U4910 ( .A1(mem_17__17_), .A2(n2784), .A3(n3139), .ZN(n2427) );
  AND3_X4 U4911 ( .A1(mem_25__17_), .A2(n2769), .A3(n3139), .ZN(n2428) );
  AND3_X4 U4912 ( .A1(mem_1__18_), .A2(n2784), .A3(n3139), .ZN(n2429) );
  AND3_X4 U4913 ( .A1(mem_9__18_), .A2(n2769), .A3(n3139), .ZN(n2430) );
  AND2_X4 U4914 ( .A1(n3103), .A2(n3085), .ZN(n2431) );
  AND3_X4 U4915 ( .A1(mem_8__0_), .A2(n2288), .A3(n3146), .ZN(n2432) );
  AND3_X4 U4916 ( .A1(mem_16__0_), .A2(n2296), .A3(n3146), .ZN(n2433) );
  AND3_X4 U4917 ( .A1(mem_24__0_), .A2(n2264), .A3(n3147), .ZN(n2434) );
  AND3_X4 U4918 ( .A1(mem_16__1_), .A2(n2302), .A3(n3148), .ZN(n2435) );
  AND3_X4 U4919 ( .A1(mem_24__1_), .A2(n2301), .A3(n3148), .ZN(n2436) );
  AND3_X4 U4920 ( .A1(mem_8__2_), .A2(n2295), .A3(n3148), .ZN(n2437) );
  AND3_X4 U4921 ( .A1(mem_16__2_), .A2(n2261), .A3(n3148), .ZN(n2438) );
  AND3_X4 U4922 ( .A1(mem_24__2_), .A2(n2241), .A3(n3148), .ZN(n2439) );
  AND3_X4 U4923 ( .A1(mem_8__3_), .A2(n2273), .A3(n3149), .ZN(n2440) );
  AND3_X4 U4924 ( .A1(mem_16__3_), .A2(n2260), .A3(n3149), .ZN(n2441) );
  AND3_X4 U4925 ( .A1(mem_24__3_), .A2(n2270), .A3(n3149), .ZN(n2442) );
  AND3_X4 U4926 ( .A1(mem_8__4_), .A2(n2283), .A3(n3149), .ZN(n2443) );
  AND3_X4 U4927 ( .A1(mem_16__4_), .A2(n2277), .A3(n3147), .ZN(n2444) );
  AND3_X4 U4928 ( .A1(mem_8__5_), .A2(n2279), .A3(n3146), .ZN(n2445) );
  AND3_X4 U4929 ( .A1(mem_16__5_), .A2(n2278), .A3(n3146), .ZN(n2446) );
  AND3_X4 U4930 ( .A1(mem_8__6_), .A2(n2270), .A3(n3150), .ZN(n2447) );
  AND3_X4 U4931 ( .A1(mem_16__6_), .A2(n2256), .A3(n3150), .ZN(n2448) );
  AND3_X4 U4932 ( .A1(mem_24__6_), .A2(n2264), .A3(n3150), .ZN(n2449) );
  AND3_X4 U4933 ( .A1(mem_8__7_), .A2(n2271), .A3(n3150), .ZN(n2450) );
  AND3_X4 U4934 ( .A1(mem_16__7_), .A2(n2259), .A3(n3151), .ZN(n2451) );
  AND3_X4 U4935 ( .A1(mem_24__7_), .A2(n2268), .A3(n3151), .ZN(n2452) );
  AND3_X4 U4936 ( .A1(mem_8__8_), .A2(n2272), .A3(n3151), .ZN(n2453) );
  AND3_X4 U4937 ( .A1(mem_16__8_), .A2(n2258), .A3(n3151), .ZN(n2454) );
  AND3_X4 U4938 ( .A1(mem_24__8_), .A2(n2253), .A3(n3141), .ZN(n2455) );
  AND3_X4 U4939 ( .A1(mem_8__9_), .A2(n2268), .A3(n3147), .ZN(n2456) );
  AND3_X4 U4940 ( .A1(mem_16__9_), .A2(n2273), .A3(n3140), .ZN(n2457) );
  AND3_X4 U4941 ( .A1(mem_24__9_), .A2(n2262), .A3(n3140), .ZN(n2458) );
  AND3_X4 U4942 ( .A1(mem_8__10_), .A2(n2295), .A3(n3152), .ZN(n2459) );
  AND3_X4 U4943 ( .A1(mem_16__10_), .A2(n2297), .A3(n3152), .ZN(n2460) );
  AND3_X4 U4944 ( .A1(mem_24__10_), .A2(n2265), .A3(n3152), .ZN(n2461) );
  AND3_X4 U4945 ( .A1(mem_8__11_), .A2(n2294), .A3(n3152), .ZN(n2462) );
  AND3_X4 U4946 ( .A1(mem_16__11_), .A2(n2298), .A3(n3152), .ZN(n2463) );
  AND3_X4 U4947 ( .A1(mem_24__11_), .A2(n2262), .A3(n3140), .ZN(n2464) );
  AND3_X4 U4948 ( .A1(mem_8__13_), .A2(n2291), .A3(n3141), .ZN(n2465) );
  AND3_X4 U4949 ( .A1(mem_16__13_), .A2(n2276), .A3(n3150), .ZN(n2466) );
  AND3_X4 U4950 ( .A1(mem_24__13_), .A2(n2267), .A3(n3150), .ZN(n2467) );
  AND3_X4 U4951 ( .A1(mem_8__14_), .A2(n2292), .A3(n3153), .ZN(n2468) );
  AND3_X4 U4952 ( .A1(mem_16__14_), .A2(n2274), .A3(n3153), .ZN(n2469) );
  AND3_X4 U4953 ( .A1(mem_24__14_), .A2(n2254), .A3(n3153), .ZN(n2470) );
  AND3_X4 U4954 ( .A1(mem_8__15_), .A2(n2290), .A3(n3143), .ZN(n2471) );
  AND3_X4 U4955 ( .A1(mem_16__18_), .A2(n2284), .A3(n3140), .ZN(n2472) );
  AND3_X4 U4956 ( .A1(mem_24__18_), .A2(n2243), .A3(n3140), .ZN(n2473) );
  AND3_X4 U4957 ( .A1(mem_8__19_), .A2(n2297), .A3(n3140), .ZN(n2474) );
  AND3_X4 U4958 ( .A1(mem_16__19_), .A2(n2300), .A3(n3140), .ZN(n2475) );
  AND3_X4 U4959 ( .A1(mem_24__19_), .A2(n2266), .A3(n3141), .ZN(n2476) );
  AND3_X4 U4960 ( .A1(mem_8__20_), .A2(n2286), .A3(n3141), .ZN(n2477) );
  AND3_X4 U4961 ( .A1(mem_16__20_), .A2(n2271), .A3(n3141), .ZN(n2478) );
  AND3_X4 U4962 ( .A1(mem_24__20_), .A2(n2265), .A3(n3141), .ZN(n2479) );
  AND3_X4 U4963 ( .A1(mem_8__21_), .A2(n2289), .A3(n3142), .ZN(n2480) );
  AND3_X4 U4964 ( .A1(mem_16__21_), .A2(n2272), .A3(n3142), .ZN(n2481) );
  AND3_X4 U4965 ( .A1(mem_24__21_), .A2(n2252), .A3(n3142), .ZN(n2482) );
  AND3_X4 U4966 ( .A1(mem_1__0_), .A2(n2766), .A3(n3144), .ZN(n2483) );
  AND3_X4 U4967 ( .A1(mem_1__3_), .A2(n2767), .A3(n3149), .ZN(n2484) );
  AND3_X4 U4968 ( .A1(mem_1__4_), .A2(n2767), .A3(n3149), .ZN(n2485) );
  AND3_X4 U4969 ( .A1(mem_1__5_), .A2(n2767), .A3(n3146), .ZN(n2486) );
  AND3_X4 U4970 ( .A1(mem_1__6_), .A2(n2768), .A3(n3150), .ZN(n2487) );
  AND3_X4 U4971 ( .A1(mem_1__7_), .A2(n2768), .A3(n3150), .ZN(n2488) );
  AND3_X4 U4972 ( .A1(mem_1__8_), .A2(n2768), .A3(n3151), .ZN(n2489) );
  AND3_X4 U4973 ( .A1(mem_1__9_), .A2(n2769), .A3(n3147), .ZN(n2490) );
  AND3_X4 U4974 ( .A1(mem_1__11_), .A2(n2769), .A3(n3152), .ZN(n2491) );
  AND3_X4 U4975 ( .A1(mem_1__13_), .A2(n2784), .A3(n3153), .ZN(n2492) );
  AND3_X4 U4976 ( .A1(mem_1__14_), .A2(n2769), .A3(n3141), .ZN(n2493) );
  AND3_X4 U4977 ( .A1(mem_1__15_), .A2(n2769), .A3(n3153), .ZN(n2494) );
  AND3_X4 U4978 ( .A1(mem_1__19_), .A2(n2766), .A3(n3140), .ZN(n2495) );
  AND3_X4 U4979 ( .A1(mem_1__20_), .A2(n2766), .A3(n3141), .ZN(n2496) );
  AND3_X4 U4980 ( .A1(mem_1__21_), .A2(n2766), .A3(n3141), .ZN(n2497) );
  AND3_X4 U4981 ( .A1(n2784), .A2(mem_1__10_), .A3(n3140), .ZN(n2498) );
  AND3_X4 U4982 ( .A1(mem_5__1_), .A2(n3156), .A3(n3154), .ZN(n2499) );
  INV_X4 U4983 ( .A(rs1[1]), .ZN(n3084) );
  AND3_X4 U4984 ( .A1(mem_25__23_), .A2(n2866), .A3(n3073), .ZN(n2500) );
  INV_X4 U4985 ( .A(n3118), .ZN(n3113) );
  INV_X4 U4986 ( .A(n3117), .ZN(n3116) );
  INV_X8 U4987 ( .A(n2774), .ZN(n2767) );
  INV_X4 U4988 ( .A(n5737), .ZN(n2847) );
  INV_X16 U4989 ( .A(n2790), .ZN(n2789) );
  AND3_X4 U4990 ( .A1(mem_24__5_), .A2(n2250), .A3(n3149), .ZN(n2501) );
  AND3_X4 U4991 ( .A1(mem_24__4_), .A2(n2260), .A3(n3148), .ZN(n2502) );
  INV_X4 U4992 ( .A(n3135), .ZN(n3124) );
  INV_X4 U4993 ( .A(n3119), .ZN(n3152) );
  INV_X4 U4994 ( .A(n3124), .ZN(n3151) );
  INV_X4 U4995 ( .A(n1048), .ZN(n2942) );
  INV_X4 U4996 ( .A(n1015), .ZN(n2946) );
  INV_X4 U4997 ( .A(n72), .ZN(n3051) );
  INV_X4 U4998 ( .A(n6), .ZN(n3055) );
  INV_X4 U4999 ( .A(n914), .ZN(n2958) );
  INV_X4 U5000 ( .A(n880), .ZN(n2962) );
  INV_X4 U5001 ( .A(n781), .ZN(n2974) );
  INV_X4 U5002 ( .A(n747), .ZN(n2978) );
  INV_X4 U5003 ( .A(n613), .ZN(n2993) );
  INV_X4 U5004 ( .A(n579), .ZN(n2997) );
  INV_X4 U5005 ( .A(n479), .ZN(n3009) );
  INV_X4 U5006 ( .A(n445), .ZN(n3013) );
  INV_X4 U5007 ( .A(n311), .ZN(n3028) );
  INV_X4 U5008 ( .A(n277), .ZN(n3032) );
  INV_X4 U5009 ( .A(n981), .ZN(n2950) );
  INV_X4 U5010 ( .A(n410), .ZN(n3017) );
  AND2_X4 U5011 ( .A1(n3063), .A2(n3073), .ZN(n2503) );
  AND2_X4 U5012 ( .A1(n3067), .A2(n3062), .ZN(n2504) );
  INV_X8 U5013 ( .A(n2864), .ZN(n2862) );
  INV_X8 U5014 ( .A(n2864), .ZN(n2863) );
  INV_X16 U5015 ( .A(n2785), .ZN(n2774) );
  INV_X4 U5016 ( .A(rs1[0]), .ZN(n3108) );
  INV_X4 U5017 ( .A(rs1[0]), .ZN(n3106) );
  INV_X4 U5018 ( .A(rs1[0]), .ZN(n3105) );
  INV_X4 U5019 ( .A(rs2[0]), .ZN(n3162) );
  INV_X4 U5020 ( .A(rs2[0]), .ZN(n3161) );
  INV_X16 U5021 ( .A(n2840), .ZN(n2832) );
  INV_X16 U5022 ( .A(n2840), .ZN(n2833) );
  INV_X8 U5023 ( .A(n2811), .ZN(n2809) );
  INV_X8 U5024 ( .A(n2811), .ZN(n2807) );
  INV_X4 U5025 ( .A(rs2[1]), .ZN(n3154) );
  INV_X4 U5026 ( .A(rs1[1]), .ZN(n3085) );
  INV_X4 U5027 ( .A(n3085), .ZN(n3074) );
  INV_X4 U5028 ( .A(n3085), .ZN(n3075) );
  INV_X4 U5029 ( .A(n3084), .ZN(n3076) );
  XNOR2_X2 U5030 ( .A(rs1[3]), .B(rd[3]), .ZN(n2505) );
  AND3_X4 U5031 ( .A1(mem_16__15_), .A2(n2282), .A3(n3138), .ZN(n2506) );
  AND3_X4 U5032 ( .A1(mem_24__15_), .A2(n2242), .A3(n3138), .ZN(n2507) );
  AND3_X4 U5033 ( .A1(mem_0__16_), .A2(n2314), .A3(n3138), .ZN(n2508) );
  AND3_X4 U5034 ( .A1(mem_8__16_), .A2(n2280), .A3(n3138), .ZN(n2509) );
  AND3_X4 U5035 ( .A1(mem_16__16_), .A2(n2285), .A3(n3138), .ZN(n2510) );
  AND3_X4 U5036 ( .A1(mem_24__16_), .A2(n2300), .A3(n3139), .ZN(n2511) );
  AND3_X4 U5037 ( .A1(mem_0__17_), .A2(n2306), .A3(n3139), .ZN(n2512) );
  AND3_X4 U5038 ( .A1(mem_8__17_), .A2(n2282), .A3(n3139), .ZN(n2513) );
  AND3_X4 U5039 ( .A1(mem_16__17_), .A2(n2274), .A3(n3139), .ZN(n2514) );
  AND3_X4 U5040 ( .A1(mem_24__17_), .A2(n2240), .A3(n3139), .ZN(n2515) );
  AND3_X4 U5041 ( .A1(mem_0__18_), .A2(n2307), .A3(n3139), .ZN(n2516) );
  INV_X4 U5042 ( .A(n6146), .ZN(n2875) );
  INV_X16 U5043 ( .A(n2875), .ZN(n2873) );
  AND3_X4 U5044 ( .A1(mem_8__23_), .A2(n2848), .A3(n3073), .ZN(n2517) );
  AND3_X4 U5045 ( .A1(mem_16__23_), .A2(n2848), .A3(n3073), .ZN(n2518) );
  AND3_X4 U5046 ( .A1(mem_8__24_), .A2(n2848), .A3(n3073), .ZN(n2519) );
  AND3_X4 U5047 ( .A1(mem_16__24_), .A2(n2848), .A3(n3072), .ZN(n2520) );
  AND3_X4 U5048 ( .A1(mem_24__24_), .A2(n2848), .A3(n3072), .ZN(n2521) );
  AND3_X4 U5049 ( .A1(mem_8__25_), .A2(n2848), .A3(n3072), .ZN(n2522) );
  AND3_X4 U5050 ( .A1(mem_16__25_), .A2(n2848), .A3(n3072), .ZN(n2523) );
  AND3_X4 U5051 ( .A1(mem_24__25_), .A2(n2849), .A3(n3072), .ZN(n2524) );
  AND3_X4 U5052 ( .A1(mem_8__26_), .A2(n2849), .A3(n3073), .ZN(n2525) );
  AND3_X4 U5053 ( .A1(mem_16__26_), .A2(n2849), .A3(n3073), .ZN(n2526) );
  AND3_X4 U5054 ( .A1(mem_24__26_), .A2(n2849), .A3(n3073), .ZN(n2527) );
  AND3_X4 U5055 ( .A1(mem_8__27_), .A2(n2849), .A3(n3071), .ZN(n2528) );
  AND3_X4 U5056 ( .A1(mem_16__27_), .A2(n2849), .A3(n3071), .ZN(n2529) );
  AND3_X4 U5057 ( .A1(mem_24__27_), .A2(n2849), .A3(n3071), .ZN(n2530) );
  AND3_X4 U5058 ( .A1(mem_8__28_), .A2(n2849), .A3(n3071), .ZN(n2531) );
  AND3_X4 U5059 ( .A1(mem_16__28_), .A2(n2849), .A3(n3071), .ZN(n2532) );
  AND3_X4 U5060 ( .A1(mem_24__28_), .A2(n2850), .A3(n3070), .ZN(n2533) );
  AND3_X4 U5061 ( .A1(mem_8__29_), .A2(n2850), .A3(n3070), .ZN(n2534) );
  AND3_X4 U5062 ( .A1(mem_16__29_), .A2(n2850), .A3(n3070), .ZN(n2535) );
  AND3_X4 U5063 ( .A1(mem_24__29_), .A2(n2850), .A3(n3070), .ZN(n2536) );
  AND3_X4 U5064 ( .A1(mem_8__30_), .A2(n2850), .A3(n3070), .ZN(n2537) );
  AND3_X4 U5065 ( .A1(mem_16__30_), .A2(n2850), .A3(n3070), .ZN(n2538) );
  AND3_X4 U5066 ( .A1(mem_24__30_), .A2(n2850), .A3(n3070), .ZN(n2539) );
  AND3_X4 U5067 ( .A1(mem_8__31_), .A2(n2850), .A3(n3071), .ZN(n2540) );
  AND3_X4 U5068 ( .A1(mem_16__31_), .A2(n2850), .A3(n3071), .ZN(n2541) );
  AND3_X4 U5069 ( .A1(mem_24__31_), .A2(n2851), .A3(n3072), .ZN(n2542) );
  AND3_X4 U5070 ( .A1(mem_0__23_), .A2(n2848), .A3(n3073), .ZN(n2543) );
  AND3_X4 U5071 ( .A1(mem_0__24_), .A2(n2848), .A3(n3073), .ZN(n2544) );
  AND3_X4 U5072 ( .A1(mem_0__25_), .A2(n2848), .A3(n3072), .ZN(n2545) );
  AND3_X4 U5073 ( .A1(mem_0__26_), .A2(n2849), .A3(n3072), .ZN(n2546) );
  AND3_X4 U5074 ( .A1(mem_0__27_), .A2(n2849), .A3(n3073), .ZN(n2547) );
  AND3_X4 U5075 ( .A1(mem_0__28_), .A2(n2849), .A3(n3071), .ZN(n2548) );
  AND3_X4 U5076 ( .A1(mem_0__29_), .A2(n2850), .A3(n3070), .ZN(n2549) );
  AND3_X4 U5077 ( .A1(mem_0__30_), .A2(n2850), .A3(n3070), .ZN(n2550) );
  AND3_X4 U5078 ( .A1(mem_0__31_), .A2(n2850), .A3(n3071), .ZN(n2551) );
  AND3_X4 U5079 ( .A1(mem_8__18_), .A2(n2296), .A3(n3140), .ZN(n2552) );
  AND3_X4 U5080 ( .A1(mem_9__0_), .A2(n2768), .A3(n3144), .ZN(n2553) );
  AND3_X4 U5081 ( .A1(mem_17__0_), .A2(n2768), .A3(n3146), .ZN(n2554) );
  AND3_X4 U5082 ( .A1(mem_25__0_), .A2(n2767), .A3(n3143), .ZN(n2555) );
  AND3_X4 U5083 ( .A1(mem_17__1_), .A2(n2767), .A3(n3148), .ZN(n2556) );
  AND3_X4 U5084 ( .A1(mem_25__1_), .A2(n2767), .A3(n3148), .ZN(n2557) );
  AND3_X4 U5085 ( .A1(mem_9__2_), .A2(n2767), .A3(n3148), .ZN(n2558) );
  AND3_X4 U5086 ( .A1(mem_17__2_), .A2(n2767), .A3(n3148), .ZN(n2559) );
  AND3_X4 U5087 ( .A1(mem_25__2_), .A2(n2767), .A3(n3148), .ZN(n2560) );
  AND3_X4 U5088 ( .A1(mem_9__3_), .A2(n2767), .A3(n3149), .ZN(n2561) );
  AND3_X4 U5089 ( .A1(mem_17__3_), .A2(n2767), .A3(n3149), .ZN(n2562) );
  AND3_X4 U5090 ( .A1(mem_25__3_), .A2(n2767), .A3(n3149), .ZN(n2563) );
  AND3_X4 U5091 ( .A1(mem_9__4_), .A2(n2767), .A3(n3149), .ZN(n2564) );
  AND3_X4 U5092 ( .A1(mem_17__4_), .A2(n2767), .A3(n3143), .ZN(n2565) );
  AND3_X4 U5093 ( .A1(mem_9__5_), .A2(n2767), .A3(n3144), .ZN(n2566) );
  AND3_X4 U5094 ( .A1(mem_17__5_), .A2(n2768), .A3(n3145), .ZN(n2567) );
  AND3_X4 U5095 ( .A1(mem_9__6_), .A2(n2768), .A3(n3150), .ZN(n2568) );
  AND3_X4 U5096 ( .A1(mem_17__6_), .A2(n2768), .A3(n3150), .ZN(n2569) );
  AND3_X4 U5097 ( .A1(mem_25__6_), .A2(n2768), .A3(n3150), .ZN(n2570) );
  AND3_X4 U5098 ( .A1(mem_9__7_), .A2(n2768), .A3(n3150), .ZN(n2571) );
  AND3_X4 U5099 ( .A1(mem_17__7_), .A2(n2768), .A3(n3151), .ZN(n2572) );
  AND3_X4 U5100 ( .A1(mem_25__7_), .A2(n2768), .A3(n3151), .ZN(n2573) );
  AND3_X4 U5101 ( .A1(mem_9__8_), .A2(n2767), .A3(n3151), .ZN(n2574) );
  AND3_X4 U5102 ( .A1(mem_17__8_), .A2(n2767), .A3(n3151), .ZN(n2575) );
  AND3_X4 U5103 ( .A1(mem_25__8_), .A2(n2767), .A3(n3151), .ZN(n2576) );
  AND3_X4 U5104 ( .A1(mem_9__9_), .A2(n2769), .A3(n3140), .ZN(n2577) );
  AND3_X4 U5105 ( .A1(mem_17__9_), .A2(n2769), .A3(n3147), .ZN(n2578) );
  AND3_X4 U5106 ( .A1(mem_25__9_), .A2(n2769), .A3(n3141), .ZN(n2579) );
  AND3_X4 U5107 ( .A1(mem_9__10_), .A2(n2769), .A3(n3141), .ZN(n2580) );
  AND3_X4 U5108 ( .A1(mem_17__10_), .A2(n2769), .A3(n3152), .ZN(n2581) );
  AND3_X4 U5109 ( .A1(mem_25__10_), .A2(n2769), .A3(n3152), .ZN(n2582) );
  AND3_X4 U5110 ( .A1(mem_9__11_), .A2(n2769), .A3(n3152), .ZN(n2583) );
  AND3_X4 U5111 ( .A1(mem_17__11_), .A2(n2768), .A3(n3152), .ZN(n2584) );
  AND3_X4 U5112 ( .A1(mem_25__11_), .A2(n2768), .A3(n3152), .ZN(n2585) );
  AND3_X4 U5113 ( .A1(mem_9__13_), .A2(n2769), .A3(n3150), .ZN(n2586) );
  AND3_X4 U5114 ( .A1(mem_17__13_), .A2(n2769), .A3(n3153), .ZN(n2587) );
  AND3_X4 U5115 ( .A1(mem_25__13_), .A2(n2769), .A3(n3140), .ZN(n2588) );
  AND3_X4 U5116 ( .A1(mem_9__14_), .A2(n2769), .A3(n3153), .ZN(n2589) );
  AND3_X4 U5117 ( .A1(mem_17__14_), .A2(n2769), .A3(n3153), .ZN(n2590) );
  AND3_X4 U5118 ( .A1(mem_25__14_), .A2(n2769), .A3(n3153), .ZN(n2591) );
  AND3_X4 U5119 ( .A1(mem_9__15_), .A2(n2769), .A3(n3153), .ZN(n2592) );
  AND3_X4 U5120 ( .A1(mem_17__18_), .A2(n2784), .A3(n3140), .ZN(n2593) );
  AND3_X4 U5121 ( .A1(mem_25__18_), .A2(n2769), .A3(n3140), .ZN(n2594) );
  AND3_X4 U5122 ( .A1(mem_9__19_), .A2(n2766), .A3(n3140), .ZN(n2595) );
  AND3_X4 U5123 ( .A1(mem_17__19_), .A2(n2766), .A3(n3140), .ZN(n2596) );
  AND3_X4 U5124 ( .A1(mem_25__19_), .A2(n2766), .A3(n3140), .ZN(n2597) );
  AND3_X4 U5125 ( .A1(mem_9__20_), .A2(n2766), .A3(n3141), .ZN(n2598) );
  AND3_X4 U5126 ( .A1(mem_17__20_), .A2(n2766), .A3(n3141), .ZN(n2599) );
  AND3_X4 U5127 ( .A1(mem_25__20_), .A2(n2766), .A3(n3141), .ZN(n2600) );
  AND3_X4 U5128 ( .A1(mem_9__21_), .A2(n2766), .A3(n3141), .ZN(n2601) );
  AND3_X4 U5129 ( .A1(mem_17__21_), .A2(n2766), .A3(n3142), .ZN(n2602) );
  AND3_X4 U5130 ( .A1(mem_25__21_), .A2(n2766), .A3(n3142), .ZN(n2603) );
  AND3_X4 U5131 ( .A1(mem_0__0_), .A2(n2240), .A3(n3146), .ZN(n2604) );
  AND3_X4 U5132 ( .A1(mem_0__2_), .A2(n2303), .A3(n3148), .ZN(n2605) );
  AND3_X4 U5133 ( .A1(mem_0__3_), .A2(n2248), .A3(n3149), .ZN(n2606) );
  AND3_X4 U5134 ( .A1(mem_0__4_), .A2(n2247), .A3(n3149), .ZN(n2607) );
  AND3_X4 U5135 ( .A1(mem_0__5_), .A2(n2313), .A3(n3147), .ZN(n2608) );
  AND3_X4 U5136 ( .A1(mem_0__6_), .A2(n2310), .A3(n3150), .ZN(n2609) );
  AND3_X4 U5137 ( .A1(mem_0__7_), .A2(n2312), .A3(n3150), .ZN(n2610) );
  AND3_X4 U5138 ( .A1(mem_0__8_), .A2(n2315), .A3(n3151), .ZN(n2611) );
  AND3_X4 U5139 ( .A1(mem_0__9_), .A2(n2242), .A3(n3141), .ZN(n2612) );
  AND3_X4 U5140 ( .A1(mem_0__11_), .A2(n2243), .A3(n3152), .ZN(n2613) );
  AND3_X4 U5141 ( .A1(mem_0__13_), .A2(n2308), .A3(n3150), .ZN(n2614) );
  AND3_X4 U5142 ( .A1(mem_0__14_), .A2(n2241), .A3(n3153), .ZN(n2615) );
  AND3_X4 U5143 ( .A1(mem_0__15_), .A2(n2309), .A3(n3153), .ZN(n2616) );
  AND3_X4 U5144 ( .A1(mem_0__19_), .A2(n2316), .A3(n3140), .ZN(n2617) );
  AND3_X4 U5145 ( .A1(mem_0__20_), .A2(n2244), .A3(n3141), .ZN(n2618) );
  AND3_X4 U5146 ( .A1(mem_0__21_), .A2(n2246), .A3(n3141), .ZN(n2619) );
  AND3_X4 U5147 ( .A1(n2266), .A2(mem_0__10_), .A3(n3149), .ZN(n2620) );
  INV_X4 U5148 ( .A(rs1[2]), .ZN(n3069) );
  INV_X4 U5149 ( .A(n3068), .ZN(n3066) );
  INV_X4 U5150 ( .A(n3068), .ZN(n3065) );
  AND2_X4 U5151 ( .A1(n3111), .A2(n3116), .ZN(n2621) );
  AND3_X4 U5152 ( .A1(mem_4__1_), .A2(n3162), .A3(n3155), .ZN(n2622) );
  AND3_X4 U5153 ( .A1(mem_1__1_), .A2(n3156), .A3(n3155), .ZN(n2623) );
  AND2_X4 U5154 ( .A1(n2621), .A2(n3151), .ZN(n2624) );
  INV_X4 U5155 ( .A(n2379), .ZN(n2940) );
  INV_X4 U5156 ( .A(n2379), .ZN(n2941) );
  AND3_X4 U5157 ( .A1(mem_24__23_), .A2(n2848), .A3(n3073), .ZN(n2625) );
  AND3_X4 U5158 ( .A1(mem_25__5_), .A2(n2767), .A3(n3149), .ZN(n2626) );
  AND3_X4 U5159 ( .A1(mem_25__4_), .A2(n2767), .A3(n3148), .ZN(n2627) );
  OR2_X4 U5160 ( .A1(mem_20__1_), .A2(n2320), .ZN(n2628) );
  OR2_X4 U5161 ( .A1(mem_28__1_), .A2(n2319), .ZN(n2629) );
  INV_X4 U5162 ( .A(rs1[4]), .ZN(n3062) );
  INV_X4 U5163 ( .A(n3062), .ZN(n3060) );
  INV_X4 U5164 ( .A(n3062), .ZN(n3061) );
  INV_X4 U5165 ( .A(n3062), .ZN(n3059) );
  INV_X4 U5166 ( .A(n947), .ZN(n2957) );
  INV_X4 U5167 ( .A(n2957), .ZN(n2954) );
  INV_X4 U5168 ( .A(n2957), .ZN(n2955) );
  INV_X4 U5169 ( .A(n2957), .ZN(n2956) );
  INV_X4 U5170 ( .A(n847), .ZN(n2969) );
  INV_X4 U5171 ( .A(n2969), .ZN(n2966) );
  INV_X4 U5172 ( .A(n2969), .ZN(n2967) );
  INV_X4 U5173 ( .A(n2969), .ZN(n2968) );
  INV_X4 U5174 ( .A(n814), .ZN(n2973) );
  INV_X4 U5175 ( .A(n2973), .ZN(n2970) );
  INV_X4 U5176 ( .A(n2973), .ZN(n2971) );
  INV_X4 U5177 ( .A(n2973), .ZN(n2972) );
  INV_X4 U5178 ( .A(n2363), .ZN(n2982) );
  INV_X4 U5179 ( .A(n2363), .ZN(n2983) );
  INV_X4 U5180 ( .A(n679), .ZN(n2988) );
  INV_X4 U5181 ( .A(n2988), .ZN(n2985) );
  INV_X4 U5182 ( .A(n2988), .ZN(n2986) );
  INV_X4 U5183 ( .A(n2988), .ZN(n2987) );
  INV_X4 U5184 ( .A(n646), .ZN(n2992) );
  INV_X4 U5185 ( .A(n2992), .ZN(n2989) );
  INV_X4 U5186 ( .A(n2992), .ZN(n2990) );
  INV_X4 U5187 ( .A(n2992), .ZN(n2991) );
  INV_X4 U5188 ( .A(n2993), .ZN(n2995) );
  INV_X4 U5189 ( .A(n2993), .ZN(n2994) );
  INV_X4 U5190 ( .A(n2993), .ZN(n2996) );
  INV_X4 U5191 ( .A(n545), .ZN(n3004) );
  INV_X4 U5192 ( .A(n3004), .ZN(n3001) );
  INV_X4 U5193 ( .A(n3004), .ZN(n3002) );
  INV_X4 U5194 ( .A(n3004), .ZN(n3003) );
  INV_X4 U5195 ( .A(n512), .ZN(n3008) );
  INV_X4 U5196 ( .A(n3008), .ZN(n3005) );
  INV_X4 U5197 ( .A(n3008), .ZN(n3006) );
  INV_X4 U5198 ( .A(n3008), .ZN(n3007) );
  INV_X4 U5199 ( .A(n3013), .ZN(n3014) );
  INV_X4 U5200 ( .A(n3013), .ZN(n3015) );
  INV_X4 U5201 ( .A(n3013), .ZN(n3016) );
  INV_X4 U5202 ( .A(n3017), .ZN(n3019) );
  INV_X4 U5203 ( .A(n3017), .ZN(n3018) );
  INV_X4 U5204 ( .A(n3017), .ZN(n3020) );
  INV_X4 U5205 ( .A(n377), .ZN(n3024) );
  INV_X4 U5206 ( .A(n3024), .ZN(n3021) );
  INV_X4 U5207 ( .A(n3024), .ZN(n3022) );
  INV_X4 U5208 ( .A(n3024), .ZN(n3023) );
  INV_X4 U5209 ( .A(n2359), .ZN(n3025) );
  INV_X4 U5210 ( .A(n2359), .ZN(n3026) );
  INV_X4 U5211 ( .A(n3028), .ZN(n3030) );
  INV_X4 U5212 ( .A(n3028), .ZN(n3029) );
  INV_X4 U5213 ( .A(n3028), .ZN(n3031) );
  INV_X4 U5214 ( .A(n3032), .ZN(n3034) );
  INV_X4 U5215 ( .A(n3032), .ZN(n3033) );
  INV_X4 U5216 ( .A(n3032), .ZN(n3035) );
  INV_X4 U5217 ( .A(n2360), .ZN(n3036) );
  INV_X4 U5218 ( .A(n2360), .ZN(n3037) );
  INV_X4 U5219 ( .A(n2361), .ZN(n3039) );
  INV_X4 U5220 ( .A(n2361), .ZN(n3040) );
  INV_X4 U5221 ( .A(n2362), .ZN(n3042) );
  INV_X4 U5222 ( .A(n2362), .ZN(n3043) );
  INV_X4 U5223 ( .A(n2358), .ZN(n3045) );
  INV_X4 U5224 ( .A(n2358), .ZN(n3046) );
  INV_X4 U5225 ( .A(n2357), .ZN(n3048) );
  INV_X4 U5226 ( .A(n2357), .ZN(n3049) );
  INV_X4 U5227 ( .A(n3051), .ZN(n3052) );
  INV_X4 U5228 ( .A(n3051), .ZN(n3053) );
  INV_X4 U5229 ( .A(n3051), .ZN(n3054) );
  INV_X4 U5230 ( .A(n3055), .ZN(n3056) );
  INV_X4 U5231 ( .A(n3055), .ZN(n3057) );
  INV_X4 U5232 ( .A(n3055), .ZN(n3058) );
  INV_X4 U5233 ( .A(n2942), .ZN(n2945) );
  INV_X4 U5234 ( .A(n2942), .ZN(n2944) );
  INV_X4 U5235 ( .A(n2942), .ZN(n2943) );
  INV_X4 U5236 ( .A(n2946), .ZN(n2949) );
  INV_X4 U5237 ( .A(n2946), .ZN(n2948) );
  INV_X4 U5238 ( .A(n2946), .ZN(n2947) );
  INV_X4 U5239 ( .A(n2950), .ZN(n2953) );
  INV_X4 U5240 ( .A(n2950), .ZN(n2952) );
  INV_X4 U5241 ( .A(n2950), .ZN(n2951) );
  INV_X4 U5242 ( .A(n2958), .ZN(n2961) );
  INV_X4 U5243 ( .A(n2958), .ZN(n2960) );
  INV_X4 U5244 ( .A(n2958), .ZN(n2959) );
  INV_X4 U5245 ( .A(n2962), .ZN(n2965) );
  INV_X4 U5246 ( .A(n2962), .ZN(n2964) );
  INV_X4 U5247 ( .A(n2962), .ZN(n2963) );
  INV_X4 U5248 ( .A(n2974), .ZN(n2977) );
  INV_X4 U5249 ( .A(n2974), .ZN(n2976) );
  INV_X4 U5250 ( .A(n2974), .ZN(n2975) );
  INV_X4 U5251 ( .A(n2978), .ZN(n2981) );
  INV_X4 U5252 ( .A(n2978), .ZN(n2980) );
  INV_X4 U5253 ( .A(n2978), .ZN(n2979) );
  INV_X4 U5254 ( .A(n2997), .ZN(n3000) );
  INV_X4 U5255 ( .A(n2997), .ZN(n2999) );
  INV_X4 U5256 ( .A(n2997), .ZN(n2998) );
  INV_X4 U5257 ( .A(n3009), .ZN(n3012) );
  INV_X4 U5258 ( .A(n3009), .ZN(n3011) );
  INV_X4 U5259 ( .A(n3009), .ZN(n3010) );
  INV_X4 U5260 ( .A(n5737), .ZN(n2842) );
  INV_X4 U5261 ( .A(rs2[3]), .ZN(n3117) );
  INV_X4 U5262 ( .A(n3117), .ZN(n3115) );
  INV_X16 U5263 ( .A(n2870), .ZN(n2867) );
  INV_X8 U5264 ( .A(n2763), .ZN(n2762) );
  INV_X4 U5265 ( .A(rs2[4]), .ZN(n3112) );
  INV_X4 U5266 ( .A(rs1[3]), .ZN(n3064) );
  INV_X4 U5267 ( .A(wData[9]), .ZN(n2920) );
  INV_X4 U5268 ( .A(wData[9]), .ZN(n2921) );
  INV_X4 U5269 ( .A(wData[0]), .ZN(n2938) );
  INV_X4 U5270 ( .A(wData[0]), .ZN(n2939) );
  INV_X4 U5271 ( .A(wData[10]), .ZN(n2918) );
  INV_X4 U5272 ( .A(wData[10]), .ZN(n2919) );
  INV_X4 U5273 ( .A(wData[11]), .ZN(n2916) );
  INV_X4 U5274 ( .A(wData[11]), .ZN(n2917) );
  INV_X4 U5275 ( .A(wData[12]), .ZN(n2914) );
  INV_X4 U5276 ( .A(wData[12]), .ZN(n2915) );
  INV_X4 U5277 ( .A(wData[13]), .ZN(n2912) );
  INV_X4 U5278 ( .A(wData[13]), .ZN(n2913) );
  INV_X4 U5279 ( .A(wData[14]), .ZN(n2910) );
  INV_X4 U5280 ( .A(wData[14]), .ZN(n2911) );
  INV_X4 U5281 ( .A(wData[15]), .ZN(n2908) );
  INV_X4 U5282 ( .A(wData[15]), .ZN(n2909) );
  INV_X4 U5283 ( .A(wData[16]), .ZN(n2906) );
  INV_X4 U5284 ( .A(wData[16]), .ZN(n2907) );
  INV_X4 U5285 ( .A(wData[17]), .ZN(n2904) );
  INV_X4 U5286 ( .A(wData[17]), .ZN(n2905) );
  INV_X4 U5287 ( .A(wData[18]), .ZN(n2902) );
  INV_X4 U5288 ( .A(wData[18]), .ZN(n2903) );
  INV_X4 U5289 ( .A(wData[19]), .ZN(n2900) );
  INV_X4 U5290 ( .A(wData[19]), .ZN(n2901) );
  INV_X4 U5291 ( .A(wData[1]), .ZN(n2936) );
  INV_X4 U5292 ( .A(wData[1]), .ZN(n2937) );
  INV_X4 U5293 ( .A(wData[20]), .ZN(n2898) );
  INV_X4 U5294 ( .A(wData[20]), .ZN(n2899) );
  INV_X4 U5295 ( .A(wData[21]), .ZN(n2896) );
  INV_X4 U5296 ( .A(wData[21]), .ZN(n2897) );
  INV_X4 U5297 ( .A(wData[22]), .ZN(n2894) );
  INV_X4 U5298 ( .A(wData[22]), .ZN(n2895) );
  INV_X4 U5299 ( .A(wData[23]), .ZN(n2892) );
  INV_X4 U5300 ( .A(wData[23]), .ZN(n2893) );
  INV_X4 U5301 ( .A(wData[24]), .ZN(n2890) );
  INV_X4 U5302 ( .A(wData[24]), .ZN(n2891) );
  INV_X4 U5303 ( .A(wData[25]), .ZN(n2888) );
  INV_X4 U5304 ( .A(wData[25]), .ZN(n2889) );
  INV_X4 U5305 ( .A(wData[26]), .ZN(n2886) );
  INV_X4 U5306 ( .A(wData[26]), .ZN(n2887) );
  INV_X4 U5307 ( .A(wData[27]), .ZN(n2884) );
  INV_X4 U5308 ( .A(wData[27]), .ZN(n2885) );
  INV_X4 U5309 ( .A(wData[28]), .ZN(n2882) );
  INV_X4 U5310 ( .A(wData[28]), .ZN(n2883) );
  INV_X4 U5311 ( .A(wData[29]), .ZN(n2880) );
  INV_X4 U5312 ( .A(wData[29]), .ZN(n2881) );
  INV_X4 U5313 ( .A(wData[2]), .ZN(n2934) );
  INV_X4 U5314 ( .A(wData[2]), .ZN(n2935) );
  INV_X4 U5315 ( .A(wData[30]), .ZN(n2878) );
  INV_X4 U5316 ( .A(wData[30]), .ZN(n2879) );
  INV_X4 U5317 ( .A(wData[31]), .ZN(n2876) );
  INV_X4 U5318 ( .A(wData[31]), .ZN(n2877) );
  INV_X4 U5319 ( .A(wData[3]), .ZN(n2932) );
  INV_X4 U5320 ( .A(wData[3]), .ZN(n2933) );
  INV_X4 U5321 ( .A(wData[4]), .ZN(n2930) );
  INV_X4 U5322 ( .A(wData[4]), .ZN(n2931) );
  INV_X4 U5323 ( .A(wData[5]), .ZN(n2928) );
  INV_X4 U5324 ( .A(wData[5]), .ZN(n2929) );
  INV_X4 U5325 ( .A(wData[6]), .ZN(n2926) );
  INV_X4 U5326 ( .A(wData[6]), .ZN(n2927) );
  INV_X4 U5327 ( .A(wData[7]), .ZN(n2924) );
  INV_X4 U5328 ( .A(wData[7]), .ZN(n2925) );
  INV_X4 U5329 ( .A(wData[8]), .ZN(n2922) );
  INV_X4 U5330 ( .A(wData[8]), .ZN(n2923) );
  NAND2_X1 U5331 ( .A1(mem_19__27_), .A2(n2981), .ZN(n760) );
  NOR2_X2 U5332 ( .A1(mem_19__27_), .A2(n2857), .ZN(n5974) );
  NAND2_X1 U5333 ( .A1(mem_19__24_), .A2(n2979), .ZN(n763) );
  NOR2_X2 U5334 ( .A1(mem_19__24_), .A2(n2856), .ZN(n5854) );
  NAND2_X1 U5335 ( .A1(mem_12__27_), .A2(n2953), .ZN(n994) );
  NOR2_X2 U5336 ( .A1(mem_12__27_), .A2(n2853), .ZN(n5965) );
  NAND2_X1 U5337 ( .A1(mem_12__24_), .A2(n2951), .ZN(n997) );
  NOR2_X2 U5338 ( .A1(mem_12__24_), .A2(n2853), .ZN(n5845) );
  NAND2_X1 U5339 ( .A1(mem_19__29_), .A2(n2980), .ZN(n758) );
  NOR2_X2 U5340 ( .A1(mem_19__29_), .A2(n2856), .ZN(n6054) );
  NAND2_X1 U5341 ( .A1(mem_19__28_), .A2(n2981), .ZN(n759) );
  NOR2_X2 U5342 ( .A1(mem_19__28_), .A2(n2857), .ZN(n6014) );
  NAND2_X1 U5343 ( .A1(mem_19__25_), .A2(n747), .ZN(n762) );
  NOR2_X2 U5344 ( .A1(mem_19__25_), .A2(n2856), .ZN(n5894) );
  NAND2_X1 U5345 ( .A1(mem_19__23_), .A2(n747), .ZN(n764) );
  NOR2_X2 U5346 ( .A1(mem_19__23_), .A2(n2856), .ZN(n5814) );
  NAND2_X1 U5347 ( .A1(mem_19__31_), .A2(n2981), .ZN(n755) );
  NOR2_X2 U5348 ( .A1(mem_19__31_), .A2(n2857), .ZN(n6134) );
  NAND2_X1 U5349 ( .A1(mem_19__30_), .A2(n747), .ZN(n756) );
  NOR2_X2 U5350 ( .A1(mem_19__30_), .A2(n2856), .ZN(n6094) );
  MUX2_X2 U5351 ( .A(n4419), .B(n4418), .S(n3113), .Z(n4420) );
  MUX2_X2 U5352 ( .A(n4230), .B(n4229), .S(n3114), .Z(n4231) );
  NAND2_X1 U5353 ( .A1(mem_14__27_), .A2(n2961), .ZN(n927) );
  NOR2_X2 U5354 ( .A1(mem_14__27_), .A2(n2873), .ZN(n5967) );
  NAND2_X1 U5355 ( .A1(mem_14__24_), .A2(n2959), .ZN(n930) );
  NOR2_X2 U5356 ( .A1(mem_14__24_), .A2(n2873), .ZN(n5847) );
  NAND2_X1 U5357 ( .A1(mem_12__28_), .A2(n2952), .ZN(n993) );
  NOR2_X2 U5358 ( .A1(mem_12__28_), .A2(n2854), .ZN(n6005) );
  NAND2_X1 U5359 ( .A1(mem_12__25_), .A2(n2953), .ZN(n996) );
  NOR2_X2 U5360 ( .A1(mem_12__25_), .A2(n2852), .ZN(n5885) );
  NAND2_X1 U5361 ( .A1(mem_12__23_), .A2(n981), .ZN(n998) );
  NOR2_X2 U5362 ( .A1(mem_12__23_), .A2(n2853), .ZN(n5805) );
  NAND2_X1 U5363 ( .A1(mem_12__31_), .A2(n2953), .ZN(n989) );
  NOR2_X2 U5364 ( .A1(mem_12__31_), .A2(n2854), .ZN(n6125) );
  NAND2_X1 U5365 ( .A1(mem_12__30_), .A2(n981), .ZN(n990) );
  NOR2_X2 U5366 ( .A1(mem_12__30_), .A2(n2854), .ZN(n6085) );
  NAND2_X1 U5367 ( .A1(mem_12__29_), .A2(n981), .ZN(n992) );
  NOR2_X2 U5368 ( .A1(mem_12__29_), .A2(n2854), .ZN(n6045) );
  NAND2_X1 U5369 ( .A1(mem_12__26_), .A2(n981), .ZN(n995) );
  NOR2_X2 U5370 ( .A1(mem_12__26_), .A2(n2852), .ZN(n5925) );
  NAND2_X4 U5371 ( .A1(n4583), .A2(n4582), .ZN(n4592) );
  NAND2_X1 U5372 ( .A1(mem_28__26_), .A2(n3020), .ZN(n424) );
  NOR2_X2 U5373 ( .A1(mem_28__26_), .A2(n2852), .ZN(n5943) );
  NAND2_X4 U5374 ( .A1(n4394), .A2(n4393), .ZN(n4403) );
  NAND2_X4 U5375 ( .A1(n4205), .A2(n4204), .ZN(n4214) );
  INV_X4 U5376 ( .A(n2630), .ZN(n2631) );
  MUX2_X2 U5377 ( .A(n4545), .B(n4544), .S(n3113), .Z(n4546) );
  MUX2_X2 U5378 ( .A(n4293), .B(n4292), .S(n3114), .Z(n4294) );
  MUX2_X2 U5379 ( .A(n4167), .B(n4166), .S(n3114), .Z(n4168) );
  MUX2_X2 U5380 ( .A(n4676), .B(n4675), .S(n3113), .Z(n4677) );
  NAND2_X1 U5381 ( .A1(mem_14__30_), .A2(n2960), .ZN(n923) );
  NOR2_X2 U5382 ( .A1(mem_14__30_), .A2(n2874), .ZN(n6087) );
  NAND2_X1 U5383 ( .A1(mem_14__28_), .A2(n2961), .ZN(n926) );
  NOR2_X2 U5384 ( .A1(mem_14__28_), .A2(n2873), .ZN(n6007) );
  NAND2_X1 U5385 ( .A1(mem_14__26_), .A2(n914), .ZN(n928) );
  NOR2_X2 U5386 ( .A1(mem_14__26_), .A2(n2874), .ZN(n5927) );
  NAND2_X1 U5387 ( .A1(mem_14__25_), .A2(n914), .ZN(n929) );
  NOR2_X2 U5388 ( .A1(mem_14__25_), .A2(n2873), .ZN(n5887) );
  NAND2_X1 U5389 ( .A1(mem_14__23_), .A2(n914), .ZN(n931) );
  NOR2_X2 U5390 ( .A1(mem_14__23_), .A2(n2873), .ZN(n5807) );
  NAND2_X1 U5391 ( .A1(mem_14__31_), .A2(n2961), .ZN(n922) );
  NOR2_X2 U5392 ( .A1(mem_14__31_), .A2(n2874), .ZN(n6127) );
  NAND2_X1 U5393 ( .A1(mem_14__29_), .A2(n914), .ZN(n925) );
  NOR2_X2 U5394 ( .A1(mem_14__29_), .A2(n2874), .ZN(n6047) );
  NAND2_X4 U5395 ( .A1(n4646), .A2(n4645), .ZN(n4655) );
  NAND2_X4 U5396 ( .A1(n4142), .A2(n4141), .ZN(n4151) );
  NAND2_X4 U5397 ( .A1(n4520), .A2(n4519), .ZN(n4529) );
  NAND2_X4 U5398 ( .A1(n4457), .A2(n4456), .ZN(n4466) );
  NAND2_X4 U5399 ( .A1(n4268), .A2(n4267), .ZN(n4277) );
  NAND2_X1 U5400 ( .A1(mem_30__26_), .A2(n3031), .ZN(n325) );
  NOR2_X2 U5401 ( .A1(mem_30__26_), .A2(n6146), .ZN(n5945) );
  NAND2_X1 U5402 ( .A1(mem_11__27_), .A2(n2949), .ZN(n1028) );
  NOR2_X2 U5403 ( .A1(mem_11__27_), .A2(n2857), .ZN(n5964) );
  NAND2_X1 U5404 ( .A1(mem_11__24_), .A2(n2947), .ZN(n1031) );
  NOR2_X2 U5405 ( .A1(mem_11__24_), .A2(n2856), .ZN(n5844) );
  NAND2_X4 U5406 ( .A1(n4588), .A2(n4587), .ZN(n4591) );
  NAND2_X1 U5407 ( .A1(mem_11__30_), .A2(n2948), .ZN(n1024) );
  NOR2_X1 U5408 ( .A1(mem_11__30_), .A2(n2856), .ZN(n6084) );
  NAND2_X1 U5409 ( .A1(mem_11__28_), .A2(n2949), .ZN(n1027) );
  NOR2_X1 U5410 ( .A1(mem_11__28_), .A2(n2857), .ZN(n6004) );
  NAND2_X1 U5411 ( .A1(mem_11__26_), .A2(n1015), .ZN(n1029) );
  NOR2_X1 U5412 ( .A1(mem_11__26_), .A2(n2857), .ZN(n5924) );
  NAND2_X1 U5413 ( .A1(mem_11__25_), .A2(n1015), .ZN(n1030) );
  NOR2_X1 U5414 ( .A1(mem_11__25_), .A2(n2856), .ZN(n5884) );
  NAND2_X1 U5415 ( .A1(mem_11__23_), .A2(n1015), .ZN(n1032) );
  NOR2_X1 U5416 ( .A1(mem_11__23_), .A2(n2856), .ZN(n5804) );
  NAND2_X1 U5417 ( .A1(mem_11__31_), .A2(n2949), .ZN(n1023) );
  NOR2_X1 U5418 ( .A1(mem_11__31_), .A2(n2857), .ZN(n6124) );
  NAND2_X1 U5419 ( .A1(mem_11__29_), .A2(n1015), .ZN(n1026) );
  NOR2_X1 U5420 ( .A1(mem_11__29_), .A2(n2856), .ZN(n6044) );
  NAND2_X4 U5421 ( .A1(n4525), .A2(n4524), .ZN(n4528) );
  NAND2_X4 U5422 ( .A1(n4462), .A2(n4461), .ZN(n4465) );
  INV_X4 U5423 ( .A(n2632), .ZN(n2633) );
  NAND2_X4 U5424 ( .A1(n4273), .A2(n4272), .ZN(n4276) );
  NAND2_X4 U5425 ( .A1(n4651), .A2(n4650), .ZN(n4654) );
  NAND2_X1 U5426 ( .A1(mem_15__27_), .A2(n2965), .ZN(n893) );
  OAI21_X1 U5427 ( .B1(mem_15__27_), .B2(n2862), .A(n2860), .ZN(n5969) );
  NAND2_X1 U5428 ( .A1(mem_15__24_), .A2(n2963), .ZN(n896) );
  OAI21_X1 U5429 ( .B1(mem_15__24_), .B2(n2863), .A(n2859), .ZN(n5849) );
  NAND2_X1 U5430 ( .A1(mem_23__30_), .A2(n3000), .ZN(n588) );
  OAI21_X1 U5431 ( .B1(mem_23__30_), .B2(n2863), .A(n2858), .ZN(n6099) );
  NAND2_X1 U5432 ( .A1(mem_10__27_), .A2(n2945), .ZN(n1061) );
  NOR3_X1 U5433 ( .A1(n3087), .A2(n3065), .A3(mem_10__27_), .ZN(n5966) );
  NAND2_X1 U5434 ( .A1(n2943), .A2(mem_10__24_), .ZN(n1064) );
  NOR3_X1 U5435 ( .A1(n3088), .A2(n3065), .A3(mem_10__24_), .ZN(n5846) );
  NAND2_X1 U5436 ( .A1(mem_23__27_), .A2(n2998), .ZN(n592) );
  OAI21_X1 U5437 ( .B1(mem_23__27_), .B2(n2862), .A(n2860), .ZN(n5979) );
  NAND2_X1 U5438 ( .A1(mem_23__24_), .A2(n2999), .ZN(n595) );
  OAI21_X1 U5439 ( .B1(mem_23__24_), .B2(n2863), .A(n2859), .ZN(n5859) );
  NAND2_X1 U5440 ( .A1(mem_18__30_), .A2(n2977), .ZN(n790) );
  NOR3_X1 U5441 ( .A1(n3086), .A2(n3066), .A3(mem_18__30_), .ZN(n6096) );
  NAND2_X1 U5442 ( .A1(mem_18__27_), .A2(n2975), .ZN(n794) );
  NOR3_X1 U5443 ( .A1(n3087), .A2(n3065), .A3(mem_18__27_), .ZN(n5976) );
  NAND2_X1 U5444 ( .A1(mem_18__24_), .A2(n2976), .ZN(n797) );
  NOR3_X1 U5445 ( .A1(n3088), .A2(n3065), .A3(mem_18__24_), .ZN(n5856) );
  NAND2_X1 U5446 ( .A1(mem_15__30_), .A2(n2964), .ZN(n889) );
  OAI21_X1 U5447 ( .B1(mem_15__30_), .B2(n2863), .A(n2860), .ZN(n6089) );
  NAND2_X1 U5448 ( .A1(mem_15__28_), .A2(n2965), .ZN(n892) );
  OAI21_X1 U5449 ( .B1(mem_15__28_), .B2(n2862), .A(n2860), .ZN(n6009) );
  NAND2_X1 U5450 ( .A1(mem_15__26_), .A2(n880), .ZN(n894) );
  OAI21_X1 U5451 ( .B1(mem_15__26_), .B2(n2862), .A(n2860), .ZN(n5929) );
  NAND2_X1 U5452 ( .A1(n880), .A2(mem_15__25_), .ZN(n895) );
  OAI21_X1 U5453 ( .B1(mem_15__25_), .B2(n2863), .A(n2859), .ZN(n5889) );
  NAND2_X1 U5454 ( .A1(mem_15__23_), .A2(n880), .ZN(n897) );
  OAI21_X1 U5455 ( .B1(mem_15__23_), .B2(n2863), .A(n2859), .ZN(n5809) );
  NAND2_X1 U5456 ( .A1(mem_15__31_), .A2(n2965), .ZN(n888) );
  OAI21_X1 U5457 ( .B1(mem_15__31_), .B2(n2863), .A(n2860), .ZN(n6129) );
  NAND2_X1 U5458 ( .A1(mem_15__29_), .A2(n880), .ZN(n891) );
  OAI21_X1 U5459 ( .B1(mem_15__29_), .B2(n2863), .A(n2858), .ZN(n6049) );
  INV_X4 U5460 ( .A(n2634), .ZN(n2635) );
  INV_X4 U5461 ( .A(n2636), .ZN(n2637) );
  NAND2_X1 U5462 ( .A1(mem_10__28_), .A2(n2944), .ZN(n1060) );
  NOR3_X1 U5463 ( .A1(n3087), .A2(n3066), .A3(mem_10__28_), .ZN(n6006) );
  NAND2_X1 U5464 ( .A1(n2945), .A2(mem_10__26_), .ZN(n1062) );
  NOR3_X1 U5465 ( .A1(n3087), .A2(n3065), .A3(mem_10__26_), .ZN(n5926) );
  NAND2_X1 U5466 ( .A1(mem_10__25_), .A2(n1048), .ZN(n1063) );
  NOR3_X1 U5467 ( .A1(n3088), .A2(n3065), .A3(mem_10__25_), .ZN(n5886) );
  NAND2_X1 U5468 ( .A1(mem_10__23_), .A2(n1048), .ZN(n1065) );
  NOR3_X1 U5469 ( .A1(n3088), .A2(n3065), .A3(mem_10__23_), .ZN(n5806) );
  NAND2_X1 U5470 ( .A1(mem_23__31_), .A2(n3000), .ZN(n587) );
  OAI21_X1 U5471 ( .B1(mem_23__31_), .B2(n2863), .A(n2858), .ZN(n6139) );
  NAND2_X1 U5472 ( .A1(mem_23__29_), .A2(n3000), .ZN(n590) );
  OAI21_X1 U5473 ( .B1(mem_23__29_), .B2(n2863), .A(n2858), .ZN(n6059) );
  NAND2_X1 U5474 ( .A1(mem_23__28_), .A2(n579), .ZN(n591) );
  OAI21_X1 U5475 ( .B1(mem_23__28_), .B2(n2862), .A(n2860), .ZN(n6019) );
  NAND2_X1 U5476 ( .A1(mem_31__26_), .A2(n3035), .ZN(n291) );
  OAI21_X2 U5477 ( .B1(mem_31__26_), .B2(n2862), .A(n2860), .ZN(n5947) );
  NAND2_X1 U5478 ( .A1(mem_23__25_), .A2(n579), .ZN(n594) );
  OAI21_X1 U5479 ( .B1(mem_23__25_), .B2(n2862), .A(n2860), .ZN(n5899) );
  NAND2_X1 U5480 ( .A1(mem_23__23_), .A2(n579), .ZN(n596) );
  OAI21_X1 U5481 ( .B1(mem_23__23_), .B2(n2863), .A(n2859), .ZN(n5819) );
  NAND2_X1 U5482 ( .A1(mem_10__30_), .A2(n1048), .ZN(n1057) );
  NOR3_X1 U5483 ( .A1(n3086), .A2(n3066), .A3(mem_10__30_), .ZN(n6086) );
  NAND2_X1 U5484 ( .A1(mem_10__31_), .A2(n2945), .ZN(n1056) );
  NOR3_X1 U5485 ( .A1(n3086), .A2(n3067), .A3(mem_10__31_), .ZN(n6126) );
  NAND2_X1 U5486 ( .A1(mem_10__29_), .A2(n1048), .ZN(n1059) );
  NOR3_X1 U5487 ( .A1(n3087), .A2(n3066), .A3(mem_10__29_), .ZN(n6046) );
  INV_X4 U5488 ( .A(n2638), .ZN(n2639) );
  NAND2_X1 U5489 ( .A1(mem_18__23_), .A2(n2977), .ZN(n798) );
  NOR3_X1 U5490 ( .A1(n3088), .A2(n3065), .A3(mem_18__23_), .ZN(n5816) );
  INV_X4 U5491 ( .A(n2640), .ZN(n2641) );
  INV_X4 U5492 ( .A(n2642), .ZN(n2643) );
  INV_X4 U5493 ( .A(n2644), .ZN(n2645) );
  INV_X4 U5494 ( .A(n2646), .ZN(n2647) );
  NAND2_X1 U5495 ( .A1(mem_18__31_), .A2(n2977), .ZN(n789) );
  NOR3_X1 U5496 ( .A1(n3086), .A2(n3067), .A3(mem_18__31_), .ZN(n6136) );
  INV_X4 U5497 ( .A(n2648), .ZN(n2649) );
  INV_X4 U5498 ( .A(n2650), .ZN(n2651) );
  INV_X4 U5499 ( .A(n2652), .ZN(n2653) );
  INV_X4 U5500 ( .A(n2654), .ZN(n2655) );
  INV_X4 U5501 ( .A(n2656), .ZN(n2657) );
  INV_X4 U5502 ( .A(n2658), .ZN(n2659) );
  INV_X4 U5503 ( .A(n2660), .ZN(n2661) );
  INV_X4 U5504 ( .A(n2662), .ZN(n2663) );
  INV_X4 U5505 ( .A(n2664), .ZN(n2665) );
  INV_X4 U5506 ( .A(n2666), .ZN(n2667) );
  INV_X4 U5507 ( .A(n2668), .ZN(n2669) );
  INV_X4 U5508 ( .A(n2670), .ZN(n2671) );
  INV_X4 U5509 ( .A(n2672), .ZN(n2673) );
  INV_X4 U5510 ( .A(n2674), .ZN(n2675) );
  INV_X4 U5511 ( .A(n2676), .ZN(n2677) );
  INV_X4 U5512 ( .A(n2678), .ZN(n2679) );
  INV_X4 U5513 ( .A(n2680), .ZN(n2681) );
  INV_X4 U5514 ( .A(n2682), .ZN(n2683) );
  INV_X4 U5515 ( .A(n2684), .ZN(n2685) );
  NAND2_X1 U5516 ( .A1(mem_31__28_), .A2(n3035), .ZN(n289) );
  OAI21_X2 U5517 ( .B1(mem_31__28_), .B2(n2862), .A(n2860), .ZN(n6027) );
  NAND2_X1 U5518 ( .A1(mem_31__25_), .A2(n3035), .ZN(n292) );
  OAI21_X2 U5519 ( .B1(mem_31__25_), .B2(n2862), .A(n2860), .ZN(n5907) );
  INV_X4 U5520 ( .A(n2686), .ZN(n2687) );
  INV_X4 U5521 ( .A(n2688), .ZN(n2689) );
  NAND2_X1 U5522 ( .A1(mem_23__26_), .A2(n579), .ZN(n593) );
  OAI21_X2 U5523 ( .B1(mem_23__26_), .B2(n2862), .A(n2860), .ZN(n5939) );
  INV_X4 U5524 ( .A(n2690), .ZN(n2691) );
  INV_X4 U5525 ( .A(n2692), .ZN(n2693) );
  INV_X4 U5526 ( .A(n2694), .ZN(n2695) );
  INV_X4 U5527 ( .A(n2696), .ZN(n2697) );
  INV_X4 U5528 ( .A(n2698), .ZN(n2699) );
  INV_X4 U5529 ( .A(n2700), .ZN(n2701) );
  INV_X4 U5530 ( .A(n2702), .ZN(n2703) );
  NAND2_X1 U5531 ( .A1(mem_19__26_), .A2(n747), .ZN(n761) );
  NOR2_X2 U5532 ( .A1(mem_19__26_), .A2(n2857), .ZN(n5934) );
  INV_X4 U5533 ( .A(n2704), .ZN(n2705) );
  INV_X4 U5534 ( .A(n2706), .ZN(n2707) );
  NAND2_X1 U5535 ( .A1(mem_31__23_), .A2(n3035), .ZN(n294) );
  OAI21_X2 U5536 ( .B1(mem_31__23_), .B2(n2863), .A(n2859), .ZN(n5827) );
  INV_X4 U5537 ( .A(n2708), .ZN(n2709) );
  INV_X4 U5538 ( .A(n2710), .ZN(n2711) );
  INV_X4 U5539 ( .A(n2712), .ZN(n2713) );
  INV_X4 U5540 ( .A(n2714), .ZN(n2715) );
  INV_X4 U5541 ( .A(n2716), .ZN(n2717) );
  NAND2_X1 U5542 ( .A1(mem_31__27_), .A2(n3035), .ZN(n290) );
  OAI21_X2 U5543 ( .B1(mem_31__27_), .B2(n2862), .A(n2860), .ZN(n5987) );
  NAND2_X1 U5544 ( .A1(mem_31__24_), .A2(n3035), .ZN(n293) );
  OAI21_X2 U5545 ( .B1(mem_31__24_), .B2(n2862), .A(n2859), .ZN(n5867) );
  INV_X4 U5546 ( .A(n2718), .ZN(n2719) );
  NAND2_X1 U5547 ( .A1(mem_22__26_), .A2(n2996), .ZN(n627) );
  NOR2_X1 U5548 ( .A1(mem_22__26_), .A2(n2874), .ZN(n5937) );
  INV_X4 U5549 ( .A(n2720), .ZN(n2721) );
  INV_X4 U5550 ( .A(n2722), .ZN(n2723) );
  INV_X4 U5551 ( .A(n2724), .ZN(n2725) );
  INV_X4 U5552 ( .A(n2726), .ZN(n2727) );
  INV_X4 U5553 ( .A(n2728), .ZN(n2729) );
  INV_X4 U5554 ( .A(n2730), .ZN(n2731) );
  INV_X4 U5555 ( .A(n2732), .ZN(n2733) );
  NAND2_X1 U5556 ( .A1(mem_26__24_), .A2(n3012), .ZN(n495) );
  NOR3_X1 U5557 ( .A1(n3088), .A2(n3066), .A3(mem_26__24_), .ZN(n5864) );
  INV_X4 U5558 ( .A(n2734), .ZN(n2735) );
  INV_X4 U5559 ( .A(n2736), .ZN(n2737) );
  INV_X4 U5560 ( .A(n2738), .ZN(n2739) );
  INV_X4 U5561 ( .A(n2740), .ZN(n2741) );
  INV_X4 U5562 ( .A(n2742), .ZN(n2743) );
  INV_X4 U5563 ( .A(n2744), .ZN(n2745) );
  INV_X4 U5564 ( .A(n2746), .ZN(n2747) );
  NAND2_X1 U5565 ( .A1(mem_26__23_), .A2(n3010), .ZN(n496) );
  NOR3_X1 U5566 ( .A1(n3087), .A2(n3065), .A3(mem_26__23_), .ZN(n5824) );
  INV_X4 U5567 ( .A(n2748), .ZN(n2749) );
  NAND2_X1 U5568 ( .A1(mem_26__31_), .A2(n3012), .ZN(n487) );
  NOR3_X1 U5569 ( .A1(n3088), .A2(n3067), .A3(mem_26__31_), .ZN(n6144) );
  NOR2_X4 U5570 ( .A1(n3137), .A2(n3155), .ZN(n2750) );
  NOR2_X1 U5571 ( .A1(n5164), .A2(n5749), .ZN(n5165) );
  NOR2_X1 U5572 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  INV_X4 U5573 ( .A(n3083), .ZN(n3081) );
  MUX2_X1 U5574 ( .A(n5871), .B(n5870), .S(n3063), .Z(n5872) );
  INV_X4 U5575 ( .A(n6145), .ZN(n2864) );
  INV_X4 U5576 ( .A(n3083), .ZN(n3082) );
  NOR2_X4 U5577 ( .A1(n3137), .A2(n3155), .ZN(n2751) );
  INV_X4 U5578 ( .A(n3136), .ZN(n3134) );
  NOR2_X2 U5579 ( .A1(n2762), .A2(n4469), .ZN(n4470) );
  NOR2_X2 U5580 ( .A1(n2761), .A2(n4280), .ZN(n4281) );
  NAND2_X4 U5581 ( .A1(n4408), .A2(n4407), .ZN(n4417) );
  NAND2_X4 U5582 ( .A1(n4219), .A2(n4218), .ZN(n4228) );
  NOR2_X2 U5583 ( .A1(n4158), .A2(n4157), .ZN(n4161) );
  INV_X4 U5584 ( .A(n3135), .ZN(n3125) );
  INV_X4 U5585 ( .A(n3124), .ZN(n3139) );
  INV_X4 U5586 ( .A(n3124), .ZN(n3138) );
  INV_X4 U5587 ( .A(n3135), .ZN(n3123) );
  NAND2_X4 U5588 ( .A1(n4330), .A2(n4331), .ZN(n4340) );
  MUX2_X1 U5589 ( .A(n4355), .B(n4356), .S(n3118), .Z(n4357) );
  INV_X4 U5590 ( .A(n3117), .ZN(n3114) );
  INV_X4 U5591 ( .A(rs2[3]), .ZN(n3118) );
  NOR2_X2 U5592 ( .A1(n2762), .A2(n4154), .ZN(n4155) );
  NAND2_X4 U5593 ( .A1(n4470), .A2(n4471), .ZN(n4480) );
  NOR2_X2 U5594 ( .A1(n2761), .A2(n4406), .ZN(n4407) );
  NAND2_X4 U5595 ( .A1(n4281), .A2(n4282), .ZN(n4291) );
  MUX2_X1 U5596 ( .A(n3415), .B(n3414), .S(n3116), .Z(n3416) );
  AOI211_X2 U5597 ( .C1(n3413), .C2(n3412), .A(n2626), .B(n2501), .ZN(n3414)
         );
  INV_X8 U5598 ( .A(n4657), .ZN(n2790) );
  INV_X2 U5599 ( .A(n3378), .ZN(n3379) );
  MUX2_X1 U5600 ( .A(n3375), .B(n3374), .S(n3116), .Z(n3376) );
  AOI211_X2 U5601 ( .C1(n3373), .C2(n3372), .A(n2627), .B(n2502), .ZN(n3374)
         );
  NOR2_X2 U5602 ( .A1(n2762), .A2(n4217), .ZN(n4218) );
  INV_X16 U5603 ( .A(n4660), .ZN(n2802) );
  AOI211_X2 U5604 ( .C1(n5829), .C2(n5828), .A(n2500), .B(n2625), .ZN(n5830)
         );
  NAND2_X4 U5605 ( .A1(n3067), .A2(rs1[1]), .ZN(n5749) );
  INV_X32 U5606 ( .A(n2789), .ZN(n2800) );
  INV_X32 U5607 ( .A(n2802), .ZN(n2801) );
  INV_X32 U5608 ( .A(rs2[1]), .ZN(n3155) );
  INV_X32 U5609 ( .A(n3164), .ZN(n3160) );
  INV_X32 U5610 ( .A(rs2[0]), .ZN(n3164) );
  NAND2_X2 U5611 ( .A1(n3160), .A2(n3135), .ZN(n4665) );
  NAND2_X2 U5612 ( .A1(n2751), .A2(n3160), .ZN(n4660) );
  NAND2_X2 U5613 ( .A1(n3155), .A2(n3135), .ZN(n4050) );
  NAND2_X2 U5614 ( .A1(n3160), .A2(n3155), .ZN(n4656) );
  NAND2_X2 U5615 ( .A1(n2750), .A2(n3164), .ZN(n4657) );
  MUX2_X2 U5616 ( .A(n3182), .B(n3181), .S(n3113), .Z(n3202) );
  MUX2_X2 U5617 ( .A(n3200), .B(n3199), .S(n3116), .Z(n3201) );
  MUX2_X2 U5618 ( .A(n3202), .B(n3201), .S(n3111), .Z(n3203) );
  INV_X4 U5619 ( .A(n3203), .ZN(n3207) );
  INV_X4 U5620 ( .A(regWr), .ZN(n3204) );
  NOR2_X4 U5621 ( .A1(n6171), .A2(n3204), .ZN(n4684) );
  MUX2_X2 U5622 ( .A(n3207), .B(wData[0]), .S(n2351), .Z(N193) );
  NAND2_X2 U5623 ( .A1(n3208), .A2(n3145), .ZN(n3209) );
  NAND2_X2 U5624 ( .A1(n3209), .A2(n2628), .ZN(n3212) );
  NAND2_X2 U5625 ( .A1(rs2[1]), .A2(n3160), .ZN(n3222) );
  NAND2_X2 U5626 ( .A1(rs2[1]), .A2(n3164), .ZN(n3223) );
  NAND2_X2 U5627 ( .A1(n3217), .A2(n3152), .ZN(n3218) );
  NAND2_X2 U5628 ( .A1(n3218), .A2(n2629), .ZN(n3221) );
  MUX2_X2 U5629 ( .A(n3229), .B(n3228), .S(n3115), .Z(n3259) );
  NAND2_X2 U5630 ( .A1(rs2[4]), .A2(n2354), .ZN(n3258) );
  NAND3_X2 U5631 ( .A1(n2373), .A2(n3152), .A3(n3234), .ZN(n3256) );
  OAI211_X2 U5632 ( .C1(n3238), .C2(n3237), .A(n3236), .B(n3235), .ZN(n3239)
         );
  NAND2_X2 U5633 ( .A1(n3239), .A2(n3151), .ZN(n3248) );
  NAND2_X2 U5634 ( .A1(n3242), .A2(n3164), .ZN(n3245) );
  NAND4_X2 U5635 ( .A1(n3113), .A2(n2354), .A3(n3248), .A4(n3247), .ZN(n3255)
         );
  OAI221_X2 U5636 ( .B1(mem_7__1_), .B2(n3163), .C1(mem_6__1_), .C2(n3160), 
        .A(rs2[1]), .ZN(n3250) );
  NAND4_X2 U5637 ( .A1(n2376), .A2(n2353), .A3(n3250), .A4(n3249), .ZN(n3254)
         );
  INV_X4 U5638 ( .A(n3258), .ZN(n3252) );
  NAND4_X2 U5639 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3257)
         );
  MUX2_X2 U5640 ( .A(n3277), .B(n3276), .S(n3115), .Z(n3297) );
  MUX2_X2 U5641 ( .A(n3295), .B(n3294), .S(n3115), .Z(n3296) );
  MUX2_X2 U5642 ( .A(n3297), .B(n3296), .S(n3111), .Z(n3298) );
  INV_X4 U5643 ( .A(n3298), .ZN(n3299) );
  MUX2_X2 U5644 ( .A(n3299), .B(wData[2]), .S(n2349), .Z(N195) );
  MUX2_X2 U5645 ( .A(n3317), .B(n3316), .S(n3115), .Z(n3337) );
  NOR3_X4 U5646 ( .A1(n3158), .A2(mem_26__3_), .A3(n3126), .ZN(n3328) );
  NOR2_X4 U5647 ( .A1(mem_27__3_), .A2(n2834), .ZN(n3326) );
  NOR3_X4 U5648 ( .A1(n3328), .A2(n3327), .A3(n3326), .ZN(n3333) );
  NOR3_X4 U5649 ( .A1(n3331), .A2(n3330), .A3(n3329), .ZN(n3332) );
  MUX2_X2 U5650 ( .A(n3335), .B(n3334), .S(n3116), .Z(n3336) );
  MUX2_X2 U5651 ( .A(n3337), .B(n3336), .S(rs2[4]), .Z(n3338) );
  INV_X4 U5652 ( .A(n3338), .ZN(n3339) );
  MUX2_X2 U5653 ( .A(n3339), .B(wData[3]), .S(n2349), .Z(N196) );
  MUX2_X2 U5654 ( .A(n3357), .B(n3356), .S(n3116), .Z(n3377) );
  OAI21_X4 U5655 ( .B1(mem_23__4_), .B2(n2809), .A(n2754), .ZN(n3363) );
  NOR2_X4 U5656 ( .A1(mem_21__4_), .A2(n2775), .ZN(n3362) );
  NOR2_X4 U5657 ( .A1(mem_22__4_), .A2(n2791), .ZN(n3361) );
  NOR3_X4 U5658 ( .A1(n3363), .A2(n3362), .A3(n3361), .ZN(n3364) );
  NOR2_X4 U5659 ( .A1(mem_27__4_), .A2(n2832), .ZN(n3366) );
  NOR3_X4 U5660 ( .A1(n3371), .A2(n3370), .A3(n3369), .ZN(n3372) );
  MUX2_X2 U5661 ( .A(n3377), .B(n3376), .S(n3111), .Z(n3378) );
  MUX2_X2 U5662 ( .A(n3379), .B(wData[4]), .S(n2350), .Z(N197) );
  MUX2_X2 U5663 ( .A(n3397), .B(n3396), .S(n3116), .Z(n3417) );
  NOR3_X4 U5664 ( .A1(n3403), .A2(n3402), .A3(n3401), .ZN(n3404) );
  NOR3_X4 U5665 ( .A1(n3158), .A2(mem_26__5_), .A3(n3126), .ZN(n3408) );
  NOR2_X4 U5666 ( .A1(mem_28__5_), .A2(n2318), .ZN(n3407) );
  NOR2_X4 U5667 ( .A1(mem_27__5_), .A2(n2832), .ZN(n3406) );
  NOR3_X4 U5668 ( .A1(n3408), .A2(n3407), .A3(n3406), .ZN(n3413) );
  NOR3_X4 U5669 ( .A1(n3411), .A2(n3410), .A3(n3409), .ZN(n3412) );
  MUX2_X2 U5670 ( .A(n3417), .B(n3416), .S(n3111), .Z(n3418) );
  INV_X4 U5671 ( .A(n3418), .ZN(n3419) );
  MUX2_X2 U5672 ( .A(n3419), .B(wData[5]), .S(n2351), .Z(N198) );
  NOR3_X4 U5673 ( .A1(n3433), .A2(n3432), .A3(n3431), .ZN(n3434) );
  MUX2_X2 U5674 ( .A(n3437), .B(n3436), .S(n3116), .Z(n3457) );
  NOR3_X4 U5675 ( .A1(n3158), .A2(mem_18__6_), .A3(n3127), .ZN(n3440) );
  NOR2_X4 U5676 ( .A1(mem_20__6_), .A2(n2319), .ZN(n3439) );
  NOR2_X4 U5677 ( .A1(mem_19__6_), .A2(n2832), .ZN(n3438) );
  NOR3_X4 U5678 ( .A1(n3440), .A2(n3439), .A3(n3438), .ZN(n3445) );
  NOR3_X4 U5679 ( .A1(n3443), .A2(n3442), .A3(n3441), .ZN(n3444) );
  NOR2_X4 U5680 ( .A1(mem_27__6_), .A2(n2832), .ZN(n3446) );
  NOR3_X4 U5681 ( .A1(n3448), .A2(n3447), .A3(n3446), .ZN(n3453) );
  OAI21_X4 U5682 ( .B1(mem_31__6_), .B2(n2808), .A(n2754), .ZN(n3451) );
  NOR3_X4 U5683 ( .A1(n3451), .A2(n3450), .A3(n3449), .ZN(n3452) );
  MUX2_X2 U5684 ( .A(n3455), .B(n3454), .S(n3115), .Z(n3456) );
  MUX2_X2 U5685 ( .A(n3457), .B(n3456), .S(n3111), .Z(n3458) );
  INV_X4 U5686 ( .A(n3458), .ZN(n3459) );
  MUX2_X2 U5687 ( .A(n3459), .B(wData[6]), .S(n2350), .Z(N199) );
  MUX2_X2 U5688 ( .A(n3477), .B(n3476), .S(n3116), .Z(n3497) );
  NOR2_X4 U5689 ( .A1(mem_27__7_), .A2(n2833), .ZN(n3486) );
  MUX2_X2 U5690 ( .A(n3495), .B(n3494), .S(n3116), .Z(n3496) );
  MUX2_X2 U5691 ( .A(n3497), .B(n3496), .S(n3111), .Z(n3498) );
  INV_X4 U5692 ( .A(n3498), .ZN(n3499) );
  MUX2_X2 U5693 ( .A(n3499), .B(wData[7]), .S(n2349), .Z(N200) );
  MUX2_X2 U5694 ( .A(n3517), .B(n3516), .S(n3116), .Z(n3537) );
  NOR3_X4 U5695 ( .A1(n3157), .A2(mem_26__8_), .A3(n3127), .ZN(n3528) );
  NOR2_X4 U5696 ( .A1(mem_28__8_), .A2(n2320), .ZN(n3527) );
  NOR2_X4 U5697 ( .A1(mem_27__8_), .A2(n2833), .ZN(n3526) );
  NOR3_X4 U5698 ( .A1(n3528), .A2(n3527), .A3(n3526), .ZN(n3533) );
  MUX2_X2 U5699 ( .A(n3535), .B(n3534), .S(n3116), .Z(n3536) );
  MUX2_X2 U5700 ( .A(n3537), .B(n3536), .S(n3111), .Z(n3538) );
  INV_X4 U5701 ( .A(n3538), .ZN(n3539) );
  MUX2_X2 U5702 ( .A(n3539), .B(wData[8]), .S(n2350), .Z(N201) );
  MUX2_X2 U5703 ( .A(n3557), .B(n3556), .S(n3115), .Z(n3577) );
  NOR3_X4 U5704 ( .A1(n3157), .A2(mem_18__9_), .A3(n3128), .ZN(n3560) );
  NOR2_X4 U5705 ( .A1(mem_20__9_), .A2(n2321), .ZN(n3559) );
  NOR2_X4 U5706 ( .A1(mem_19__9_), .A2(n2833), .ZN(n3558) );
  NOR3_X4 U5707 ( .A1(n3560), .A2(n3559), .A3(n3558), .ZN(n3565) );
  NOR2_X4 U5708 ( .A1(mem_27__9_), .A2(n2833), .ZN(n3566) );
  NOR3_X4 U5709 ( .A1(n3568), .A2(n3567), .A3(n3566), .ZN(n3573) );
  MUX2_X2 U5710 ( .A(n3575), .B(n3574), .S(n3115), .Z(n3576) );
  MUX2_X2 U5711 ( .A(n3577), .B(n3576), .S(n3111), .Z(n3578) );
  INV_X4 U5712 ( .A(n3578), .ZN(n3579) );
  MUX2_X2 U5713 ( .A(n3579), .B(wData[9]), .S(n2349), .Z(N202) );
  MUX2_X2 U5714 ( .A(n3597), .B(n3596), .S(n3115), .Z(n3617) );
  NOR3_X4 U5715 ( .A1(n3608), .A2(n3607), .A3(n3606), .ZN(n3613) );
  MUX2_X2 U5716 ( .A(n3615), .B(n3614), .S(n3115), .Z(n3616) );
  MUX2_X2 U5717 ( .A(n3617), .B(n3616), .S(n3111), .Z(n3618) );
  INV_X4 U5718 ( .A(n3618), .ZN(n3619) );
  MUX2_X2 U5719 ( .A(n3619), .B(wData[10]), .S(n2351), .Z(N203) );
  MUX2_X2 U5720 ( .A(n3637), .B(n3636), .S(n3115), .Z(n3657) );
  NOR3_X4 U5721 ( .A1(n3648), .A2(n3647), .A3(n3646), .ZN(n3653) );
  OAI21_X4 U5722 ( .B1(mem_31__11_), .B2(n2807), .A(n2756), .ZN(n3651) );
  NOR2_X4 U5723 ( .A1(mem_29__11_), .A2(n2777), .ZN(n3650) );
  NOR2_X4 U5724 ( .A1(mem_30__11_), .A2(n2792), .ZN(n3649) );
  NOR3_X4 U5725 ( .A1(n3651), .A2(n3650), .A3(n3649), .ZN(n3652) );
  MUX2_X2 U5726 ( .A(n3655), .B(n3654), .S(n3115), .Z(n3656) );
  MUX2_X2 U5727 ( .A(n3657), .B(n3656), .S(n3111), .Z(n3658) );
  INV_X4 U5728 ( .A(n3658), .ZN(n3659) );
  MUX2_X2 U5729 ( .A(n3659), .B(wData[11]), .S(n2351), .Z(N204) );
  MUX2_X2 U5730 ( .A(mem_20__12_), .B(mem_21__12_), .S(n3159), .Z(n3661) );
  MUX2_X2 U5731 ( .A(mem_22__12_), .B(mem_23__12_), .S(n3159), .Z(n3660) );
  MUX2_X2 U5732 ( .A(n3661), .B(n3660), .S(rs2[1]), .Z(n3663) );
  NAND2_X2 U5733 ( .A1(n2354), .A2(n2376), .ZN(n3662) );
  MUX2_X2 U5734 ( .A(mem_28__12_), .B(mem_29__12_), .S(n3159), .Z(n3665) );
  MUX2_X2 U5735 ( .A(mem_30__12_), .B(mem_31__12_), .S(n3159), .Z(n3664) );
  MUX2_X2 U5736 ( .A(n3665), .B(n3664), .S(rs2[1]), .Z(n3667) );
  NAND2_X2 U5737 ( .A1(n2353), .A2(n2418), .ZN(n3666) );
  MUX2_X2 U5738 ( .A(mem_24__12_), .B(mem_25__12_), .S(n3159), .Z(n3671) );
  MUX2_X2 U5739 ( .A(mem_26__12_), .B(mem_27__12_), .S(n3159), .Z(n3670) );
  MUX2_X2 U5740 ( .A(n3671), .B(n3670), .S(rs2[1]), .Z(n3673) );
  NAND2_X2 U5741 ( .A1(n2352), .A2(n2624), .ZN(n3672) );
  NAND2_X2 U5742 ( .A1(n2373), .A2(n3112), .ZN(n4076) );
  NAND2_X2 U5743 ( .A1(n3677), .A2(n3676), .ZN(n3700) );
  MUX2_X2 U5744 ( .A(mem_8__12_), .B(mem_9__12_), .S(n3159), .Z(n3679) );
  MUX2_X2 U5745 ( .A(mem_10__12_), .B(mem_11__12_), .S(n3159), .Z(n3678) );
  MUX2_X2 U5746 ( .A(n3679), .B(n3678), .S(rs2[1]), .Z(n3689) );
  NAND2_X2 U5747 ( .A1(n2352), .A2(n4083), .ZN(n3688) );
  MUX2_X2 U5748 ( .A(mem_16__12_), .B(mem_17__12_), .S(n3159), .Z(n3681) );
  MUX2_X2 U5749 ( .A(mem_18__12_), .B(mem_19__12_), .S(n3159), .Z(n3680) );
  MUX2_X2 U5750 ( .A(n3681), .B(n3680), .S(rs2[1]), .Z(n3687) );
  NAND2_X2 U5751 ( .A1(n2355), .A2(n2370), .ZN(n3686) );
  MUX2_X2 U5752 ( .A(mem_12__12_), .B(mem_13__12_), .S(n3159), .Z(n3683) );
  MUX2_X2 U5753 ( .A(mem_14__12_), .B(mem_15__12_), .S(n3159), .Z(n3682) );
  MUX2_X2 U5754 ( .A(n3683), .B(n3682), .S(rs2[1]), .Z(n3685) );
  NAND2_X2 U5755 ( .A1(n2355), .A2(n2380), .ZN(n3684) );
  OAI222_X2 U5756 ( .A1(n3689), .A2(n3688), .B1(n3687), .B2(n3686), .C1(n3685), 
        .C2(n3684), .ZN(n3699) );
  NAND2_X2 U5757 ( .A1(n2370), .A2(n3112), .ZN(n4094) );
  MUX2_X2 U5758 ( .A(mem_0__12_), .B(mem_1__12_), .S(n3159), .Z(n3691) );
  MUX2_X2 U5759 ( .A(mem_2__12_), .B(mem_3__12_), .S(n3159), .Z(n3690) );
  MUX2_X2 U5760 ( .A(n3691), .B(n3690), .S(rs2[1]), .Z(n3696) );
  NAND2_X2 U5761 ( .A1(n2376), .A2(n3112), .ZN(n4098) );
  MUX2_X2 U5762 ( .A(mem_4__12_), .B(mem_5__12_), .S(n3159), .Z(n3693) );
  MUX2_X2 U5763 ( .A(mem_6__12_), .B(mem_7__12_), .S(n3159), .Z(n3692) );
  MUX2_X2 U5764 ( .A(n3693), .B(n3692), .S(rs2[1]), .Z(n3694) );
  AOI22_X2 U5765 ( .A1(n3697), .A2(n3696), .B1(n3695), .B2(n3694), .ZN(n3698)
         );
  MUX2_X2 U5766 ( .A(n3718), .B(n3717), .S(n3115), .Z(n3738) );
  NOR3_X4 U5767 ( .A1(n3157), .A2(mem_26__13_), .A3(n3129), .ZN(n3729) );
  NOR2_X4 U5768 ( .A1(mem_28__13_), .A2(n2318), .ZN(n3728) );
  NOR2_X4 U5769 ( .A1(mem_27__13_), .A2(n2834), .ZN(n3727) );
  NOR3_X4 U5770 ( .A1(n3729), .A2(n3728), .A3(n3727), .ZN(n3734) );
  MUX2_X2 U5771 ( .A(n3736), .B(n3735), .S(n3115), .Z(n3737) );
  MUX2_X2 U5772 ( .A(n3738), .B(n3737), .S(n3111), .Z(n3739) );
  INV_X4 U5773 ( .A(n3739), .ZN(n3740) );
  MUX2_X2 U5774 ( .A(n3740), .B(wData[13]), .S(n2349), .Z(N206) );
  MUX2_X2 U5775 ( .A(n3758), .B(n3757), .S(n3115), .Z(n3778) );
  NOR2_X4 U5776 ( .A1(mem_27__14_), .A2(n2837), .ZN(n3767) );
  NOR3_X4 U5777 ( .A1(n3769), .A2(n3768), .A3(n3767), .ZN(n3774) );
  MUX2_X2 U5778 ( .A(n3776), .B(n3775), .S(n3115), .Z(n3777) );
  MUX2_X2 U5779 ( .A(n3778), .B(n3777), .S(n3111), .Z(n3779) );
  INV_X4 U5780 ( .A(n3779), .ZN(n3780) );
  MUX2_X2 U5781 ( .A(n3780), .B(wData[14]), .S(n2349), .Z(N207) );
  MUX2_X2 U5782 ( .A(n3798), .B(n3797), .S(n3116), .Z(n3818) );
  NOR3_X4 U5783 ( .A1(n3158), .A2(mem_18__15_), .A3(n3129), .ZN(n3801) );
  NOR2_X4 U5784 ( .A1(mem_19__15_), .A2(n2833), .ZN(n3799) );
  NOR3_X4 U5785 ( .A1(n3801), .A2(n3800), .A3(n3799), .ZN(n3806) );
  NOR3_X4 U5786 ( .A1(n3156), .A2(mem_26__15_), .A3(n3129), .ZN(n3809) );
  NOR2_X4 U5787 ( .A1(mem_28__15_), .A2(n2320), .ZN(n3808) );
  NOR2_X4 U5788 ( .A1(mem_27__15_), .A2(n2838), .ZN(n3807) );
  NOR3_X4 U5789 ( .A1(n3809), .A2(n3808), .A3(n3807), .ZN(n3814) );
  MUX2_X2 U5790 ( .A(n3816), .B(n3815), .S(n3116), .Z(n3817) );
  MUX2_X2 U5791 ( .A(n3818), .B(n3817), .S(n3111), .Z(n3819) );
  INV_X4 U5792 ( .A(n3819), .ZN(n3820) );
  MUX2_X2 U5793 ( .A(n3820), .B(wData[15]), .S(n2350), .Z(N208) );
  MUX2_X2 U5794 ( .A(n3838), .B(n3837), .S(n3116), .Z(n3858) );
  NOR3_X4 U5795 ( .A1(n3156), .A2(mem_18__16_), .A3(n3129), .ZN(n3841) );
  NOR2_X4 U5796 ( .A1(mem_20__16_), .A2(n2318), .ZN(n3840) );
  NOR2_X4 U5797 ( .A1(mem_19__16_), .A2(n2834), .ZN(n3839) );
  NOR3_X4 U5798 ( .A1(n3841), .A2(n3840), .A3(n3839), .ZN(n3846) );
  NOR3_X4 U5799 ( .A1(n3156), .A2(mem_26__16_), .A3(n3130), .ZN(n3849) );
  NOR2_X4 U5800 ( .A1(mem_27__16_), .A2(n2836), .ZN(n3847) );
  NOR3_X4 U5801 ( .A1(n3849), .A2(n3848), .A3(n3847), .ZN(n3854) );
  OAI21_X4 U5802 ( .B1(mem_31__16_), .B2(n2806), .A(n2757), .ZN(n3852) );
  MUX2_X2 U5803 ( .A(n3856), .B(n3855), .S(n3116), .Z(n3857) );
  MUX2_X2 U5804 ( .A(n3858), .B(n3857), .S(n3111), .Z(n3859) );
  INV_X4 U5805 ( .A(n3859), .ZN(n3860) );
  MUX2_X2 U5806 ( .A(n3860), .B(wData[16]), .S(n2350), .Z(N209) );
  MUX2_X2 U5807 ( .A(n3878), .B(n3877), .S(n3116), .Z(n3898) );
  OAI21_X4 U5808 ( .B1(mem_23__17_), .B2(n2806), .A(n2758), .ZN(n3884) );
  NOR2_X4 U5809 ( .A1(mem_21__17_), .A2(n2778), .ZN(n3883) );
  NOR2_X4 U5810 ( .A1(mem_22__17_), .A2(n2794), .ZN(n3882) );
  NOR3_X4 U5811 ( .A1(n3884), .A2(n3883), .A3(n3882), .ZN(n3885) );
  NOR3_X4 U5812 ( .A1(n3156), .A2(mem_26__17_), .A3(n3130), .ZN(n3889) );
  NOR2_X4 U5813 ( .A1(mem_28__17_), .A2(n2319), .ZN(n3888) );
  NOR2_X4 U5814 ( .A1(mem_27__17_), .A2(n2838), .ZN(n3887) );
  NOR3_X4 U5815 ( .A1(n3889), .A2(n3888), .A3(n3887), .ZN(n3894) );
  OAI21_X4 U5816 ( .B1(mem_31__17_), .B2(n2806), .A(n2758), .ZN(n3892) );
  NOR3_X4 U5817 ( .A1(n3892), .A2(n3891), .A3(n3890), .ZN(n3893) );
  MUX2_X2 U5818 ( .A(n3896), .B(n3895), .S(n3116), .Z(n3897) );
  MUX2_X2 U5819 ( .A(n3898), .B(n3897), .S(n3111), .Z(n3899) );
  INV_X4 U5820 ( .A(n3899), .ZN(n3900) );
  MUX2_X2 U5821 ( .A(n3900), .B(wData[17]), .S(n2349), .Z(N210) );
  OAI21_X4 U5822 ( .B1(mem_15__18_), .B2(n2806), .A(n2758), .ZN(n3914) );
  NOR2_X4 U5823 ( .A1(mem_13__18_), .A2(n2778), .ZN(n3913) );
  NOR2_X4 U5824 ( .A1(mem_14__18_), .A2(n2794), .ZN(n3912) );
  NOR3_X4 U5825 ( .A1(n3914), .A2(n3913), .A3(n3912), .ZN(n3915) );
  MUX2_X2 U5826 ( .A(n3918), .B(n3917), .S(n3116), .Z(n3938) );
  OAI21_X4 U5827 ( .B1(mem_23__18_), .B2(n2806), .A(n2758), .ZN(n3924) );
  NOR2_X4 U5828 ( .A1(mem_21__18_), .A2(n2778), .ZN(n3923) );
  NOR2_X4 U5829 ( .A1(mem_22__18_), .A2(n2794), .ZN(n3922) );
  NOR3_X4 U5830 ( .A1(n3924), .A2(n3923), .A3(n3922), .ZN(n3925) );
  OAI21_X4 U5831 ( .B1(mem_31__18_), .B2(n2806), .A(n2758), .ZN(n3932) );
  NOR3_X4 U5832 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3933) );
  MUX2_X2 U5833 ( .A(n3936), .B(n3935), .S(n3116), .Z(n3937) );
  MUX2_X2 U5834 ( .A(n3938), .B(n3937), .S(n3111), .Z(n3939) );
  INV_X4 U5835 ( .A(n3939), .ZN(n3940) );
  MUX2_X2 U5836 ( .A(n3940), .B(wData[18]), .S(n2350), .Z(N211) );
  OAI21_X4 U5837 ( .B1(mem_15__19_), .B2(n2805), .A(n2758), .ZN(n3954) );
  NOR2_X4 U5838 ( .A1(mem_13__19_), .A2(n2778), .ZN(n3953) );
  NOR2_X4 U5839 ( .A1(mem_14__19_), .A2(n2794), .ZN(n3952) );
  NOR3_X4 U5840 ( .A1(n3954), .A2(n3953), .A3(n3952), .ZN(n3955) );
  MUX2_X2 U5841 ( .A(n3958), .B(n3957), .S(n3116), .Z(n3978) );
  OAI21_X4 U5842 ( .B1(mem_31__19_), .B2(n2805), .A(n2758), .ZN(n3972) );
  NOR3_X4 U5843 ( .A1(n3972), .A2(n3971), .A3(n3970), .ZN(n3973) );
  MUX2_X2 U5844 ( .A(n3976), .B(n3975), .S(n3116), .Z(n3977) );
  MUX2_X2 U5845 ( .A(n3978), .B(n3977), .S(n3111), .Z(n3979) );
  INV_X4 U5846 ( .A(n3979), .ZN(n3980) );
  MUX2_X2 U5847 ( .A(n3980), .B(wData[19]), .S(n2351), .Z(N212) );
  MUX2_X2 U5848 ( .A(n3998), .B(n3997), .S(n3114), .Z(n4018) );
  OAI21_X4 U5849 ( .B1(mem_23__20_), .B2(n2805), .A(n2759), .ZN(n4004) );
  NOR2_X4 U5850 ( .A1(mem_21__20_), .A2(n2779), .ZN(n4003) );
  NOR2_X4 U5851 ( .A1(mem_22__20_), .A2(n2795), .ZN(n4002) );
  NOR3_X4 U5852 ( .A1(n4004), .A2(n4003), .A3(n4002), .ZN(n4005) );
  NOR3_X4 U5853 ( .A1(n4012), .A2(n4011), .A3(n4010), .ZN(n4013) );
  MUX2_X2 U5854 ( .A(n4016), .B(n4015), .S(n3114), .Z(n4017) );
  MUX2_X2 U5855 ( .A(n4018), .B(n4017), .S(n3111), .Z(n4019) );
  INV_X4 U5856 ( .A(n4019), .ZN(n4020) );
  MUX2_X2 U5857 ( .A(n4020), .B(wData[20]), .S(n2351), .Z(N213) );
  MUX2_X2 U5858 ( .A(n4038), .B(n4037), .S(n3114), .Z(n4059) );
  OAI21_X4 U5859 ( .B1(mem_31__21_), .B2(n2805), .A(n2759), .ZN(n4053) );
  NOR3_X4 U5860 ( .A1(n4053), .A2(n4052), .A3(n4051), .ZN(n4054) );
  MUX2_X2 U5861 ( .A(n4057), .B(n4056), .S(n3114), .Z(n4058) );
  MUX2_X2 U5862 ( .A(n4059), .B(n4058), .S(n3111), .Z(n4060) );
  INV_X4 U5863 ( .A(n4060), .ZN(n4061) );
  MUX2_X2 U5864 ( .A(n4061), .B(wData[21]), .S(n2349), .Z(N214) );
  MUX2_X2 U5865 ( .A(mem_20__22_), .B(mem_21__22_), .S(n3159), .Z(n4063) );
  MUX2_X2 U5866 ( .A(mem_22__22_), .B(mem_23__22_), .S(n3159), .Z(n4062) );
  MUX2_X2 U5867 ( .A(n4063), .B(n4062), .S(rs2[1]), .Z(n4065) );
  NAND2_X2 U5868 ( .A1(n2353), .A2(n2376), .ZN(n4064) );
  MUX2_X2 U5869 ( .A(mem_28__22_), .B(mem_29__22_), .S(n3160), .Z(n4067) );
  MUX2_X2 U5870 ( .A(mem_30__22_), .B(mem_31__22_), .S(n3159), .Z(n4066) );
  MUX2_X2 U5871 ( .A(n4067), .B(n4066), .S(rs2[1]), .Z(n4069) );
  NAND2_X2 U5872 ( .A1(n2354), .A2(n2418), .ZN(n4068) );
  MUX2_X2 U5873 ( .A(mem_24__22_), .B(mem_25__22_), .S(n3160), .Z(n4073) );
  MUX2_X2 U5874 ( .A(mem_26__22_), .B(mem_27__22_), .S(n3159), .Z(n4072) );
  MUX2_X2 U5875 ( .A(n4073), .B(n4072), .S(rs2[1]), .Z(n4075) );
  NAND2_X2 U5876 ( .A1(n2356), .A2(n2624), .ZN(n4074) );
  NAND2_X2 U5877 ( .A1(n4080), .A2(n4079), .ZN(n4107) );
  MUX2_X2 U5878 ( .A(mem_8__22_), .B(mem_9__22_), .S(n3160), .Z(n4082) );
  MUX2_X2 U5879 ( .A(mem_10__22_), .B(mem_11__22_), .S(n3160), .Z(n4081) );
  MUX2_X2 U5880 ( .A(n4082), .B(n4081), .S(rs2[1]), .Z(n4093) );
  NAND2_X2 U5881 ( .A1(n2355), .A2(n4083), .ZN(n4092) );
  MUX2_X2 U5882 ( .A(mem_16__22_), .B(mem_17__22_), .S(n3160), .Z(n4085) );
  MUX2_X2 U5883 ( .A(mem_18__22_), .B(mem_19__22_), .S(n3159), .Z(n4084) );
  MUX2_X2 U5884 ( .A(n4085), .B(n4084), .S(rs2[1]), .Z(n4091) );
  NAND2_X2 U5885 ( .A1(n2352), .A2(n2370), .ZN(n4090) );
  MUX2_X2 U5886 ( .A(mem_12__22_), .B(mem_13__22_), .S(n3160), .Z(n4087) );
  MUX2_X2 U5887 ( .A(mem_14__22_), .B(mem_15__22_), .S(n3160), .Z(n4086) );
  MUX2_X2 U5888 ( .A(n4087), .B(n4086), .S(rs2[1]), .Z(n4089) );
  NAND2_X2 U5889 ( .A1(n2353), .A2(n2380), .ZN(n4088) );
  OAI222_X2 U5890 ( .A1(n4093), .A2(n4092), .B1(n4091), .B2(n4090), .C1(n4089), 
        .C2(n4088), .ZN(n4106) );
  MUX2_X2 U5891 ( .A(mem_0__22_), .B(mem_1__22_), .S(n3160), .Z(n4096) );
  MUX2_X2 U5892 ( .A(mem_2__22_), .B(mem_3__22_), .S(n3160), .Z(n4095) );
  MUX2_X2 U5893 ( .A(n4096), .B(n4095), .S(rs2[1]), .Z(n4103) );
  MUX2_X2 U5894 ( .A(mem_4__22_), .B(mem_5__22_), .S(n3160), .Z(n4100) );
  MUX2_X2 U5895 ( .A(mem_6__22_), .B(mem_7__22_), .S(n3160), .Z(n4099) );
  MUX2_X2 U5896 ( .A(n4100), .B(n4099), .S(rs2[1]), .Z(n4101) );
  AOI22_X2 U5897 ( .A1(n4104), .A2(n4103), .B1(n4102), .B2(n4101), .ZN(n4105)
         );
  NAND2_X2 U5898 ( .A1(n4112), .A2(n4111), .ZN(n4121) );
  NAND2_X2 U5899 ( .A1(n4115), .A2(n3164), .ZN(n4116) );
  NAND2_X2 U5900 ( .A1(n4117), .A2(n4116), .ZN(n4120) );
  OAI211_X2 U5901 ( .C1(n4121), .C2(n4120), .A(n4119), .B(n4118), .ZN(n4137)
         );
  NOR2_X4 U5902 ( .A1(mem_15__23_), .A2(n2804), .ZN(n4124) );
  NOR2_X4 U5903 ( .A1(n2762), .A2(n4124), .ZN(n4125) );
  NAND2_X2 U5904 ( .A1(n4129), .A2(n3164), .ZN(n4130) );
  NAND3_X4 U5905 ( .A1(n2280), .A2(mem_8__23_), .A3(n3142), .ZN(n4133) );
  NAND3_X4 U5906 ( .A1(n2784), .A2(mem_9__23_), .A3(n3142), .ZN(n4132) );
  OAI211_X2 U5907 ( .C1(n4135), .C2(n4134), .A(n4133), .B(n4132), .ZN(n4136)
         );
  MUX2_X2 U5908 ( .A(n4137), .B(n4136), .S(n3114), .Z(n4169) );
  NOR2_X4 U5909 ( .A1(mem_18__23_), .A2(n3132), .ZN(n4145) );
  NAND2_X2 U5910 ( .A1(n4145), .A2(n3161), .ZN(n4146) );
  NAND3_X4 U5911 ( .A1(n2284), .A2(mem_16__23_), .A3(n3142), .ZN(n4149) );
  NOR2_X4 U5912 ( .A1(n2715), .A2(n2779), .ZN(n4153) );
  NOR2_X4 U5913 ( .A1(n2731), .A2(n2795), .ZN(n4152) );
  NAND2_X2 U5914 ( .A1(n4155), .A2(n4156), .ZN(n4165) );
  NOR2_X4 U5915 ( .A1(n2697), .A2(n2321), .ZN(n4158) );
  NOR2_X4 U5916 ( .A1(n2717), .A2(n2835), .ZN(n4157) );
  NAND2_X2 U5917 ( .A1(n4159), .A2(n3162), .ZN(n4160) );
  NAND2_X2 U5918 ( .A1(n4161), .A2(n4160), .ZN(n4164) );
  OAI211_X2 U5919 ( .C1(n4165), .C2(n4164), .A(n4163), .B(n4162), .ZN(n4166)
         );
  MUX2_X2 U5920 ( .A(n4169), .B(n4168), .S(n3111), .Z(n4170) );
  NOR2_X4 U5922 ( .A1(mem_7__24_), .A2(n2804), .ZN(n4173) );
  NOR2_X4 U5923 ( .A1(n2762), .A2(n4173), .ZN(n4174) );
  NAND2_X2 U5924 ( .A1(n4175), .A2(n4174), .ZN(n4184) );
  NAND2_X2 U5925 ( .A1(n4178), .A2(n3162), .ZN(n4179) );
  NAND2_X2 U5926 ( .A1(n4180), .A2(n4179), .ZN(n4183) );
  OAI211_X2 U5927 ( .C1(n4184), .C2(n4183), .A(n4182), .B(n4181), .ZN(n4200)
         );
  NOR2_X4 U5928 ( .A1(mem_13__24_), .A2(n2780), .ZN(n4186) );
  NOR2_X4 U5929 ( .A1(mem_14__24_), .A2(n2796), .ZN(n4185) );
  NOR2_X4 U5930 ( .A1(n4186), .A2(n4185), .ZN(n4189) );
  NOR2_X4 U5931 ( .A1(mem_15__24_), .A2(n2804), .ZN(n4187) );
  NOR2_X4 U5932 ( .A1(n2762), .A2(n4187), .ZN(n4188) );
  NOR2_X4 U5933 ( .A1(mem_11__24_), .A2(n2836), .ZN(n4190) );
  NOR2_X4 U5934 ( .A1(mem_10__24_), .A2(n3132), .ZN(n4192) );
  NAND2_X2 U5935 ( .A1(n4192), .A2(n3162), .ZN(n4193) );
  OAI211_X2 U5936 ( .C1(n4198), .C2(n4197), .A(n4196), .B(n4195), .ZN(n4199)
         );
  MUX2_X2 U5937 ( .A(n4200), .B(n4199), .S(n3114), .Z(n4232) );
  NOR2_X4 U5938 ( .A1(mem_18__24_), .A2(n3132), .ZN(n4208) );
  NAND2_X2 U5939 ( .A1(n4208), .A2(n3161), .ZN(n4209) );
  NAND3_X4 U5940 ( .A1(n2283), .A2(mem_16__24_), .A3(n3143), .ZN(n4212) );
  NAND2_X2 U5941 ( .A1(n4222), .A2(n3161), .ZN(n4223) );
  NAND2_X2 U5942 ( .A1(n4224), .A2(n4223), .ZN(n4227) );
  OAI211_X2 U5943 ( .C1(n4228), .C2(n4227), .A(n4226), .B(n4225), .ZN(n4229)
         );
  MUX2_X2 U5944 ( .A(n4232), .B(n4231), .S(n3111), .Z(n4233) );
  MUX2_X2 U5945 ( .A(n4233), .B(wData[24]), .S(n2350), .Z(N217) );
  NAND2_X2 U5946 ( .A1(n4238), .A2(n4237), .ZN(n4247) );
  NAND2_X2 U5947 ( .A1(n4241), .A2(n3162), .ZN(n4242) );
  NAND2_X2 U5948 ( .A1(n4243), .A2(n4242), .ZN(n4246) );
  OAI211_X2 U5949 ( .C1(n4247), .C2(n4246), .A(n4245), .B(n4244), .ZN(n4263)
         );
  NOR2_X4 U5950 ( .A1(mem_13__25_), .A2(n2780), .ZN(n4249) );
  NOR2_X4 U5951 ( .A1(mem_15__25_), .A2(n2804), .ZN(n4250) );
  NAND2_X2 U5952 ( .A1(n4252), .A2(n4251), .ZN(n4261) );
  NOR2_X4 U5953 ( .A1(mem_10__25_), .A2(n3132), .ZN(n4255) );
  OAI211_X2 U5954 ( .C1(n4261), .C2(n4260), .A(n4259), .B(n4258), .ZN(n4262)
         );
  MUX2_X2 U5955 ( .A(n4263), .B(n4262), .S(n3113), .Z(n4295) );
  NOR2_X4 U5956 ( .A1(mem_22__25_), .A2(n2796), .ZN(n4264) );
  NOR2_X4 U5957 ( .A1(n4265), .A2(n4264), .ZN(n4268) );
  NOR2_X4 U5958 ( .A1(mem_23__25_), .A2(n2804), .ZN(n4266) );
  NOR2_X4 U5959 ( .A1(n2762), .A2(n4266), .ZN(n4267) );
  NOR2_X4 U5960 ( .A1(mem_20__25_), .A2(n2320), .ZN(n4270) );
  NAND2_X2 U5961 ( .A1(n4271), .A2(n3162), .ZN(n4272) );
  NAND3_X4 U5962 ( .A1(n2278), .A2(mem_16__25_), .A3(n3144), .ZN(n4275) );
  OAI211_X2 U5963 ( .C1(n4277), .C2(n4276), .A(n4275), .B(n4274), .ZN(n4293)
         );
  NOR2_X4 U5964 ( .A1(n2689), .A2(n2780), .ZN(n4279) );
  NOR2_X4 U5965 ( .A1(n2721), .A2(n2796), .ZN(n4278) );
  NOR2_X4 U5966 ( .A1(n4279), .A2(n4278), .ZN(n4282) );
  NOR2_X4 U5967 ( .A1(n2637), .A2(n2804), .ZN(n4280) );
  NOR2_X4 U5968 ( .A1(n2705), .A2(n2836), .ZN(n4283) );
  NAND2_X2 U5969 ( .A1(n4285), .A2(n3161), .ZN(n4286) );
  OAI211_X2 U5970 ( .C1(n4291), .C2(n4290), .A(n4289), .B(n4288), .ZN(n4292)
         );
  MUX2_X2 U5971 ( .A(n4295), .B(n4294), .S(n3111), .Z(n4296) );
  MUX2_X2 U5972 ( .A(n4296), .B(wData[25]), .S(n2350), .Z(N218) );
  NAND2_X2 U5973 ( .A1(n4301), .A2(n4300), .ZN(n4310) );
  NAND2_X2 U5974 ( .A1(n4304), .A2(n3161), .ZN(n4305) );
  NAND2_X2 U5975 ( .A1(n4306), .A2(n4305), .ZN(n4309) );
  OAI211_X2 U5976 ( .C1(n4310), .C2(n4309), .A(n4308), .B(n4307), .ZN(n4326)
         );
  NOR2_X4 U5977 ( .A1(mem_13__26_), .A2(n2780), .ZN(n4312) );
  NOR2_X4 U5978 ( .A1(mem_14__26_), .A2(n2796), .ZN(n4311) );
  NOR2_X4 U5979 ( .A1(n4312), .A2(n4311), .ZN(n4315) );
  NOR2_X4 U5980 ( .A1(mem_15__26_), .A2(n2803), .ZN(n4313) );
  NAND2_X2 U5981 ( .A1(n4315), .A2(n4314), .ZN(n4324) );
  NOR2_X4 U5982 ( .A1(mem_10__26_), .A2(n3132), .ZN(n4318) );
  NAND2_X2 U5983 ( .A1(n4318), .A2(n3162), .ZN(n4319) );
  OAI211_X2 U5984 ( .C1(n4324), .C2(n4323), .A(n4322), .B(n4321), .ZN(n4325)
         );
  MUX2_X2 U5985 ( .A(n4326), .B(n4325), .S(n3114), .Z(n4358) );
  NOR2_X4 U5986 ( .A1(n2691), .A2(n2780), .ZN(n4328) );
  NAND2_X2 U5987 ( .A1(n4334), .A2(n3162), .ZN(n4335) );
  OAI211_X2 U5988 ( .C1(n4340), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4356)
         );
  NOR2_X4 U5989 ( .A1(mem_29__26_), .A2(n2780), .ZN(n4342) );
  NOR2_X4 U5990 ( .A1(mem_30__26_), .A2(n2796), .ZN(n4341) );
  NAND2_X2 U5991 ( .A1(n4345), .A2(n4344), .ZN(n4354) );
  NAND2_X2 U5992 ( .A1(n4348), .A2(n3161), .ZN(n4349) );
  NAND2_X2 U5993 ( .A1(n4350), .A2(n4349), .ZN(n4353) );
  OAI211_X2 U5994 ( .C1(n4354), .C2(n4353), .A(n4352), .B(n4351), .ZN(n4355)
         );
  MUX2_X2 U5995 ( .A(n4358), .B(n4357), .S(n3111), .Z(n4359) );
  NAND2_X2 U5997 ( .A1(n4364), .A2(n4363), .ZN(n4373) );
  NAND2_X2 U5998 ( .A1(n4367), .A2(n3161), .ZN(n4368) );
  NAND2_X2 U5999 ( .A1(n4369), .A2(n4368), .ZN(n4372) );
  OAI211_X2 U6000 ( .C1(n4373), .C2(n4372), .A(n4371), .B(n4370), .ZN(n4389)
         );
  NOR2_X4 U6001 ( .A1(mem_15__27_), .A2(n2803), .ZN(n4376) );
  NAND2_X2 U6002 ( .A1(n4378), .A2(n4377), .ZN(n4387) );
  NOR2_X4 U6003 ( .A1(mem_10__27_), .A2(n3133), .ZN(n4381) );
  NAND3_X4 U6004 ( .A1(n2279), .A2(mem_8__27_), .A3(n3145), .ZN(n4385) );
  NAND3_X4 U6005 ( .A1(n2771), .A2(mem_9__27_), .A3(n3145), .ZN(n4384) );
  OAI211_X2 U6006 ( .C1(n4387), .C2(n4386), .A(n4385), .B(n4384), .ZN(n4388)
         );
  MUX2_X2 U6007 ( .A(n4389), .B(n4388), .S(n3113), .Z(n4421) );
  NOR2_X4 U6008 ( .A1(mem_23__27_), .A2(n2803), .ZN(n4392) );
  NOR2_X4 U6009 ( .A1(mem_20__27_), .A2(n2321), .ZN(n4396) );
  NOR2_X4 U6010 ( .A1(mem_18__27_), .A2(n3133), .ZN(n4397) );
  NAND2_X2 U6011 ( .A1(n4397), .A2(n3162), .ZN(n4398) );
  OAI211_X2 U6012 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4419)
         );
  NAND2_X2 U6013 ( .A1(n4411), .A2(n3161), .ZN(n4412) );
  OAI211_X2 U6014 ( .C1(n4417), .C2(n4416), .A(n4415), .B(n4414), .ZN(n4418)
         );
  MUX2_X2 U6015 ( .A(n4421), .B(n4420), .S(n3111), .Z(n4422) );
  MUX2_X2 U6016 ( .A(n4422), .B(wData[27]), .S(n2351), .Z(N220) );
  NAND2_X2 U6017 ( .A1(n4427), .A2(n4426), .ZN(n4436) );
  NAND2_X2 U6018 ( .A1(n4430), .A2(n3161), .ZN(n4431) );
  NAND2_X2 U6019 ( .A1(n4432), .A2(n4431), .ZN(n4435) );
  OAI211_X2 U6020 ( .C1(n4436), .C2(n4435), .A(n4434), .B(n4433), .ZN(n4452)
         );
  NAND2_X2 U6021 ( .A1(n4441), .A2(n4440), .ZN(n4450) );
  NOR2_X4 U6022 ( .A1(mem_11__28_), .A2(n2837), .ZN(n4442) );
  NOR2_X4 U6023 ( .A1(mem_10__28_), .A2(n3133), .ZN(n4444) );
  OAI211_X2 U6024 ( .C1(n4450), .C2(n4449), .A(n4448), .B(n4447), .ZN(n4451)
         );
  MUX2_X2 U6025 ( .A(n4452), .B(n4451), .S(n3113), .Z(n4484) );
  NOR2_X4 U6026 ( .A1(mem_23__28_), .A2(n2803), .ZN(n4455) );
  NOR2_X4 U6027 ( .A1(mem_20__28_), .A2(n2319), .ZN(n4459) );
  NOR2_X4 U6028 ( .A1(mem_19__28_), .A2(n2837), .ZN(n4458) );
  NOR2_X4 U6029 ( .A1(n4459), .A2(n4458), .ZN(n4462) );
  NAND2_X2 U6030 ( .A1(n4460), .A2(n3163), .ZN(n4461) );
  NAND3_X4 U6031 ( .A1(n2277), .A2(mem_16__28_), .A3(n3146), .ZN(n4464) );
  NOR2_X4 U6032 ( .A1(n2687), .A2(n2781), .ZN(n4468) );
  NOR2_X4 U6033 ( .A1(n2635), .A2(n2803), .ZN(n4469) );
  NOR2_X4 U6034 ( .A1(n2703), .A2(n2837), .ZN(n4472) );
  NAND2_X2 U6035 ( .A1(n4474), .A2(n3161), .ZN(n4475) );
  OAI211_X2 U6036 ( .C1(n4480), .C2(n4479), .A(n4478), .B(n4477), .ZN(n4481)
         );
  MUX2_X2 U6037 ( .A(n4484), .B(n4483), .S(n3111), .Z(n4485) );
  MUX2_X2 U6038 ( .A(n4485), .B(wData[28]), .S(n2351), .Z(N221) );
  NAND2_X2 U6039 ( .A1(n4490), .A2(n4489), .ZN(n4499) );
  NAND2_X2 U6040 ( .A1(n4493), .A2(n3163), .ZN(n4494) );
  NAND2_X2 U6041 ( .A1(n4495), .A2(n4494), .ZN(n4498) );
  OAI211_X2 U6042 ( .C1(n4499), .C2(n4498), .A(n4497), .B(n4496), .ZN(n4515)
         );
  NOR2_X4 U6043 ( .A1(mem_15__29_), .A2(n2810), .ZN(n4502) );
  NOR2_X4 U6044 ( .A1(n2762), .A2(n4502), .ZN(n4503) );
  NOR2_X4 U6045 ( .A1(mem_11__29_), .A2(n2837), .ZN(n4505) );
  NOR2_X4 U6046 ( .A1(mem_10__29_), .A2(n3134), .ZN(n4507) );
  NAND2_X2 U6047 ( .A1(n4507), .A2(n3163), .ZN(n4508) );
  NAND2_X2 U6048 ( .A1(n4509), .A2(n4508), .ZN(n4512) );
  OAI211_X2 U6049 ( .C1(n4513), .C2(n4512), .A(n4511), .B(n4510), .ZN(n4514)
         );
  MUX2_X2 U6050 ( .A(n4515), .B(n4514), .S(n3113), .Z(n4547) );
  NOR2_X4 U6051 ( .A1(mem_23__29_), .A2(n2809), .ZN(n4518) );
  NOR2_X4 U6052 ( .A1(mem_20__29_), .A2(n2321), .ZN(n4522) );
  NOR2_X4 U6053 ( .A1(mem_19__29_), .A2(n2837), .ZN(n4521) );
  NOR2_X4 U6054 ( .A1(n4522), .A2(n4521), .ZN(n4525) );
  NAND2_X2 U6055 ( .A1(n4523), .A2(n3163), .ZN(n4524) );
  NAND3_X4 U6056 ( .A1(n2261), .A2(mem_16__29_), .A3(n3146), .ZN(n4527) );
  OAI211_X2 U6057 ( .C1(n4529), .C2(n4528), .A(n4527), .B(n4526), .ZN(n4545)
         );
  NOR2_X4 U6058 ( .A1(n2679), .A2(n2781), .ZN(n4531) );
  NAND2_X2 U6059 ( .A1(n4534), .A2(n4533), .ZN(n4543) );
  NOR2_X4 U6060 ( .A1(n2707), .A2(n2837), .ZN(n4535) );
  NAND2_X2 U6061 ( .A1(n4537), .A2(n3163), .ZN(n4538) );
  OAI211_X2 U6062 ( .C1(n4543), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4544)
         );
  MUX2_X2 U6063 ( .A(n4547), .B(n4546), .S(n3111), .Z(n4548) );
  MUX2_X2 U6064 ( .A(n4548), .B(wData[29]), .S(n2349), .Z(N222) );
  NAND2_X2 U6065 ( .A1(n4556), .A2(n3163), .ZN(n4557) );
  NAND2_X2 U6066 ( .A1(n4558), .A2(n4557), .ZN(n4561) );
  OAI211_X2 U6067 ( .C1(n4562), .C2(n4561), .A(n4560), .B(n4559), .ZN(n4578)
         );
  NOR2_X4 U6068 ( .A1(mem_15__30_), .A2(n2810), .ZN(n4565) );
  NOR2_X4 U6069 ( .A1(mem_10__30_), .A2(n3134), .ZN(n4570) );
  NAND2_X2 U6070 ( .A1(n4570), .A2(n3163), .ZN(n4571) );
  OAI211_X2 U6071 ( .C1(n4576), .C2(n4575), .A(n4574), .B(n4573), .ZN(n4577)
         );
  MUX2_X2 U6072 ( .A(n4578), .B(n4577), .S(n3113), .Z(n4610) );
  NOR2_X4 U6073 ( .A1(mem_23__30_), .A2(n2807), .ZN(n4581) );
  NOR2_X4 U6074 ( .A1(mem_20__30_), .A2(n2322), .ZN(n4585) );
  NOR2_X4 U6075 ( .A1(mem_18__30_), .A2(n3134), .ZN(n4586) );
  NAND2_X2 U6076 ( .A1(n4586), .A2(n3163), .ZN(n4587) );
  OAI211_X2 U6077 ( .C1(n4592), .C2(n4591), .A(n4590), .B(n4589), .ZN(n4608)
         );
  NAND2_X2 U6078 ( .A1(n4597), .A2(n4596), .ZN(n4606) );
  NAND2_X2 U6079 ( .A1(n4600), .A2(n3163), .ZN(n4601) );
  NAND2_X2 U6080 ( .A1(n4602), .A2(n4601), .ZN(n4605) );
  OAI211_X2 U6081 ( .C1(n4606), .C2(n4605), .A(n4604), .B(n4603), .ZN(n4607)
         );
  MUX2_X2 U6082 ( .A(n4608), .B(n4607), .S(n3113), .Z(n4609) );
  MUX2_X2 U6083 ( .A(n4610), .B(n4609), .S(n3111), .Z(n4611) );
  MUX2_X2 U6084 ( .A(n4611), .B(wData[30]), .S(n2351), .Z(N223) );
  NAND2_X2 U6085 ( .A1(n4619), .A2(n3163), .ZN(n4620) );
  NAND2_X2 U6086 ( .A1(n4621), .A2(n4620), .ZN(n4624) );
  OAI211_X2 U6087 ( .C1(n4625), .C2(n4624), .A(n4623), .B(n4622), .ZN(n4641)
         );
  NOR2_X4 U6088 ( .A1(mem_13__31_), .A2(n2782), .ZN(n4627) );
  NOR2_X4 U6089 ( .A1(mem_15__31_), .A2(n2810), .ZN(n4628) );
  NOR2_X4 U6090 ( .A1(mem_10__31_), .A2(n3134), .ZN(n4633) );
  NAND2_X2 U6091 ( .A1(n4633), .A2(n3163), .ZN(n4634) );
  OAI211_X2 U6092 ( .C1(n4639), .C2(n4638), .A(n4637), .B(n4636), .ZN(n4640)
         );
  MUX2_X2 U6093 ( .A(n4641), .B(n4640), .S(n3113), .Z(n4678) );
  NOR2_X4 U6094 ( .A1(mem_23__31_), .A2(n2805), .ZN(n4644) );
  NOR2_X4 U6095 ( .A1(mem_20__31_), .A2(n2319), .ZN(n4648) );
  NOR2_X4 U6096 ( .A1(mem_19__31_), .A2(n2838), .ZN(n4647) );
  NOR2_X4 U6097 ( .A1(n4648), .A2(n4647), .ZN(n4651) );
  NOR2_X4 U6098 ( .A1(mem_18__31_), .A2(n3134), .ZN(n4649) );
  NAND2_X2 U6099 ( .A1(n4649), .A2(n3163), .ZN(n4650) );
  NAND3_X4 U6100 ( .A1(n2298), .A2(mem_16__31_), .A3(n3144), .ZN(n4653) );
  NAND3_X4 U6101 ( .A1(n2772), .A2(mem_17__31_), .A3(n3146), .ZN(n4652) );
  OAI211_X2 U6102 ( .C1(n4655), .C2(n4654), .A(n4653), .B(n4652), .ZN(n4676)
         );
  NAND2_X2 U6103 ( .A1(n4663), .A2(n4662), .ZN(n4674) );
  NAND2_X2 U6104 ( .A1(n4668), .A2(n3163), .ZN(n4669) );
  OAI211_X2 U6105 ( .C1(n4674), .C2(n4673), .A(n4672), .B(n4671), .ZN(n4675)
         );
  MUX2_X2 U6106 ( .A(n4678), .B(n4677), .S(n3111), .Z(n4679) );
  MUX2_X2 U6107 ( .A(n4679), .B(wData[31]), .S(n2350), .Z(N224) );
  MUX2_X2 U6108 ( .A(mem_28__0_), .B(mem_29__0_), .S(n3088), .Z(n4680) );
  INV_X4 U6109 ( .A(n4680), .ZN(n4683) );
  MUX2_X2 U6110 ( .A(mem_30__0_), .B(mem_31__0_), .S(n3099), .Z(n4681) );
  INV_X4 U6111 ( .A(n4681), .ZN(n4682) );
  MUX2_X2 U6112 ( .A(n4683), .B(n4682), .S(n3078), .Z(n4685) );
  NAND4_X2 U6113 ( .A1(n4685), .A2(n2334), .A3(n3059), .A4(n2374), .ZN(n4695)
         );
  MUX2_X2 U6114 ( .A(mem_24__0_), .B(mem_25__0_), .S(n3099), .Z(n4686) );
  INV_X4 U6115 ( .A(n4686), .ZN(n4689) );
  MUX2_X2 U6116 ( .A(mem_26__0_), .B(mem_27__0_), .S(n3099), .Z(n4687) );
  INV_X4 U6117 ( .A(n4687), .ZN(n4688) );
  MUX2_X2 U6118 ( .A(n4689), .B(n4688), .S(n3080), .Z(n4690) );
  NAND4_X2 U6119 ( .A1(n4690), .A2(n2339), .A3(n3061), .A4(n2503), .ZN(n4694)
         );
  NAND3_X2 U6120 ( .A1(n2339), .A2(n3064), .A3(n3062), .ZN(n4691) );
  NAND3_X2 U6121 ( .A1(n4695), .A2(n4694), .A3(n4693), .ZN(n4729) );
  MUX2_X2 U6122 ( .A(mem_12__0_), .B(mem_13__0_), .S(n3099), .Z(n4696) );
  INV_X4 U6123 ( .A(n4696), .ZN(n4699) );
  MUX2_X2 U6124 ( .A(mem_14__0_), .B(mem_15__0_), .S(n3099), .Z(n4697) );
  INV_X4 U6125 ( .A(n4697), .ZN(n4698) );
  MUX2_X2 U6126 ( .A(n4699), .B(n4698), .S(n3077), .Z(n4700) );
  NAND3_X2 U6127 ( .A1(n4700), .A2(n2338), .A3(n2504), .ZN(n4719) );
  MUX2_X2 U6128 ( .A(mem_16__0_), .B(mem_17__0_), .S(n3098), .Z(n4701) );
  INV_X4 U6129 ( .A(n4701), .ZN(n4704) );
  MUX2_X2 U6130 ( .A(mem_18__0_), .B(mem_19__0_), .S(n3098), .Z(n4702) );
  INV_X4 U6131 ( .A(n4702), .ZN(n4703) );
  MUX2_X2 U6132 ( .A(n4704), .B(n4703), .S(n3078), .Z(n4705) );
  NAND3_X2 U6133 ( .A1(n4705), .A2(n2345), .A3(n2364), .ZN(n4718) );
  MUX2_X2 U6134 ( .A(mem_20__0_), .B(mem_21__0_), .S(n3098), .Z(n4706) );
  INV_X4 U6135 ( .A(n4706), .ZN(n4709) );
  MUX2_X2 U6136 ( .A(mem_22__0_), .B(mem_23__0_), .S(n3098), .Z(n4707) );
  INV_X4 U6137 ( .A(n4707), .ZN(n4708) );
  MUX2_X2 U6138 ( .A(n4709), .B(n4708), .S(n3080), .Z(n4710) );
  NAND3_X2 U6139 ( .A1(n4710), .A2(n2343), .A3(n2366), .ZN(n4717) );
  MUX2_X2 U6140 ( .A(mem_8__0_), .B(mem_9__0_), .S(n3098), .Z(n4711) );
  INV_X4 U6141 ( .A(n4711), .ZN(n4714) );
  MUX2_X2 U6142 ( .A(mem_10__0_), .B(mem_11__0_), .S(n3098), .Z(n4712) );
  INV_X4 U6143 ( .A(n4712), .ZN(n4713) );
  MUX2_X2 U6144 ( .A(n4714), .B(n4713), .S(n3079), .Z(n4715) );
  NAND3_X2 U6145 ( .A1(n4715), .A2(n2346), .A3(n2367), .ZN(n4716) );
  NAND4_X2 U6146 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4728)
         );
  MUX2_X2 U6147 ( .A(mem_0__0_), .B(mem_1__0_), .S(n3098), .Z(n4721) );
  MUX2_X2 U6148 ( .A(mem_2__0_), .B(mem_3__0_), .S(n3098), .Z(n4720) );
  MUX2_X2 U6149 ( .A(n4721), .B(n4720), .S(n3077), .Z(n4722) );
  NAND3_X2 U6150 ( .A1(n4722), .A2(n2346), .A3(n2368), .ZN(n4727) );
  MUX2_X2 U6151 ( .A(mem_4__0_), .B(mem_5__0_), .S(n3098), .Z(n4724) );
  MUX2_X2 U6152 ( .A(mem_6__0_), .B(mem_7__0_), .S(n3098), .Z(n4723) );
  MUX2_X2 U6153 ( .A(n4724), .B(n4723), .S(n3080), .Z(n4725) );
  NAND3_X2 U6154 ( .A1(n4725), .A2(n2343), .A3(n2369), .ZN(n4726) );
  OAI211_X2 U6155 ( .C1(n4729), .C2(n4728), .A(n4727), .B(n4726), .ZN(n7226)
         );
  MUX2_X2 U6156 ( .A(mem_28__1_), .B(mem_29__1_), .S(n3098), .Z(n4730) );
  INV_X4 U6157 ( .A(n4730), .ZN(n4733) );
  MUX2_X2 U6158 ( .A(mem_30__1_), .B(mem_31__1_), .S(n3098), .Z(n4731) );
  INV_X4 U6159 ( .A(n4731), .ZN(n4732) );
  MUX2_X2 U6160 ( .A(n4733), .B(n4732), .S(n3079), .Z(n4734) );
  NAND4_X2 U6161 ( .A1(n4734), .A2(n2327), .A3(n3059), .A4(n2374), .ZN(n4743)
         );
  MUX2_X2 U6162 ( .A(mem_24__1_), .B(mem_25__1_), .S(n3098), .Z(n4735) );
  INV_X4 U6163 ( .A(n4735), .ZN(n4738) );
  MUX2_X2 U6164 ( .A(mem_26__1_), .B(mem_27__1_), .S(n3098), .Z(n4736) );
  INV_X4 U6165 ( .A(n4736), .ZN(n4737) );
  MUX2_X2 U6166 ( .A(n4738), .B(n4737), .S(n3077), .Z(n4739) );
  NAND4_X2 U6167 ( .A1(n4739), .A2(n2338), .A3(n3061), .A4(n2503), .ZN(n4742)
         );
  NAND3_X2 U6168 ( .A1(n4743), .A2(n4742), .A3(n4741), .ZN(n4777) );
  MUX2_X2 U6169 ( .A(mem_12__1_), .B(mem_13__1_), .S(n3098), .Z(n4744) );
  INV_X4 U6170 ( .A(n4744), .ZN(n4747) );
  MUX2_X2 U6171 ( .A(mem_14__1_), .B(mem_15__1_), .S(n3098), .Z(n4745) );
  INV_X4 U6172 ( .A(n4745), .ZN(n4746) );
  MUX2_X2 U6173 ( .A(n4747), .B(n4746), .S(n3078), .Z(n4748) );
  NAND3_X2 U6174 ( .A1(n4748), .A2(n2329), .A3(n2504), .ZN(n4767) );
  MUX2_X2 U6175 ( .A(mem_16__1_), .B(mem_17__1_), .S(n3098), .Z(n4749) );
  INV_X4 U6176 ( .A(n4749), .ZN(n4752) );
  MUX2_X2 U6177 ( .A(mem_18__1_), .B(mem_19__1_), .S(n3098), .Z(n4750) );
  INV_X4 U6178 ( .A(n4750), .ZN(n4751) );
  MUX2_X2 U6179 ( .A(n4752), .B(n4751), .S(n3079), .Z(n4753) );
  NAND3_X2 U6180 ( .A1(n4753), .A2(n2330), .A3(n2364), .ZN(n4766) );
  MUX2_X2 U6181 ( .A(mem_20__1_), .B(mem_21__1_), .S(n3098), .Z(n4754) );
  INV_X4 U6182 ( .A(n4754), .ZN(n4757) );
  MUX2_X2 U6183 ( .A(mem_22__1_), .B(mem_23__1_), .S(n3098), .Z(n4755) );
  INV_X4 U6184 ( .A(n4755), .ZN(n4756) );
  MUX2_X2 U6185 ( .A(n4757), .B(n4756), .S(n3081), .Z(n4758) );
  NAND3_X2 U6186 ( .A1(n4758), .A2(n2342), .A3(n2366), .ZN(n4765) );
  MUX2_X2 U6187 ( .A(mem_8__1_), .B(mem_9__1_), .S(n3098), .Z(n4759) );
  INV_X4 U6188 ( .A(n4759), .ZN(n4762) );
  MUX2_X2 U6189 ( .A(mem_10__1_), .B(mem_11__1_), .S(n3097), .Z(n4760) );
  INV_X4 U6190 ( .A(n4760), .ZN(n4761) );
  MUX2_X2 U6191 ( .A(n4762), .B(n4761), .S(n3078), .Z(n4763) );
  NAND3_X2 U6192 ( .A1(n4763), .A2(n2336), .A3(n2367), .ZN(n4764) );
  NAND4_X2 U6193 ( .A1(n4767), .A2(n4766), .A3(n4765), .A4(n4764), .ZN(n4776)
         );
  MUX2_X2 U6194 ( .A(mem_0__1_), .B(mem_1__1_), .S(n3097), .Z(n4769) );
  MUX2_X2 U6195 ( .A(mem_2__1_), .B(mem_3__1_), .S(n3097), .Z(n4768) );
  MUX2_X2 U6196 ( .A(n4769), .B(n4768), .S(n3081), .Z(n4770) );
  NAND3_X2 U6197 ( .A1(n4770), .A2(n2346), .A3(n2368), .ZN(n4775) );
  MUX2_X2 U6198 ( .A(mem_4__1_), .B(mem_5__1_), .S(n3097), .Z(n4772) );
  MUX2_X2 U6199 ( .A(mem_6__1_), .B(mem_7__1_), .S(n3097), .Z(n4771) );
  MUX2_X2 U6200 ( .A(n4772), .B(n4771), .S(n3081), .Z(n4773) );
  NAND3_X2 U6201 ( .A1(n4773), .A2(n2340), .A3(n2369), .ZN(n4774) );
  OAI211_X2 U6202 ( .C1(n4777), .C2(n4776), .A(n4775), .B(n4774), .ZN(n7225)
         );
  MUX2_X2 U6203 ( .A(mem_28__2_), .B(mem_29__2_), .S(n3097), .Z(n4778) );
  INV_X4 U6204 ( .A(n4778), .ZN(n4781) );
  MUX2_X2 U6205 ( .A(mem_30__2_), .B(mem_31__2_), .S(n3097), .Z(n4779) );
  INV_X4 U6206 ( .A(n4779), .ZN(n4780) );
  MUX2_X2 U6207 ( .A(n4781), .B(n4780), .S(n3081), .Z(n4782) );
  NAND4_X2 U6208 ( .A1(n4782), .A2(n2336), .A3(n3059), .A4(n2374), .ZN(n4791)
         );
  MUX2_X2 U6209 ( .A(mem_24__2_), .B(mem_25__2_), .S(n3097), .Z(n4783) );
  INV_X4 U6210 ( .A(n4783), .ZN(n4786) );
  MUX2_X2 U6211 ( .A(mem_26__2_), .B(mem_27__2_), .S(n3097), .Z(n4784) );
  INV_X4 U6212 ( .A(n4784), .ZN(n4785) );
  MUX2_X2 U6213 ( .A(n4786), .B(n4785), .S(n3081), .Z(n4787) );
  NAND4_X2 U6214 ( .A1(n4787), .A2(n2345), .A3(n3061), .A4(n2503), .ZN(n4790)
         );
  NAND3_X2 U6215 ( .A1(n4791), .A2(n4790), .A3(n4789), .ZN(n4825) );
  MUX2_X2 U6216 ( .A(mem_12__2_), .B(mem_13__2_), .S(n3097), .Z(n4792) );
  INV_X4 U6217 ( .A(n4792), .ZN(n4795) );
  MUX2_X2 U6218 ( .A(mem_14__2_), .B(mem_15__2_), .S(n3097), .Z(n4793) );
  INV_X4 U6219 ( .A(n4793), .ZN(n4794) );
  MUX2_X2 U6220 ( .A(n4795), .B(n4794), .S(n3081), .Z(n4796) );
  NAND3_X2 U6221 ( .A1(n4796), .A2(n2327), .A3(n2504), .ZN(n4815) );
  MUX2_X2 U6222 ( .A(mem_16__2_), .B(mem_17__2_), .S(n3097), .Z(n4797) );
  INV_X4 U6223 ( .A(n4797), .ZN(n4800) );
  MUX2_X2 U6224 ( .A(mem_18__2_), .B(mem_19__2_), .S(n3097), .Z(n4798) );
  INV_X4 U6225 ( .A(n4798), .ZN(n4799) );
  MUX2_X2 U6226 ( .A(n4800), .B(n4799), .S(n3081), .Z(n4801) );
  NAND3_X2 U6227 ( .A1(n4801), .A2(n2331), .A3(n2364), .ZN(n4814) );
  MUX2_X2 U6228 ( .A(mem_20__2_), .B(mem_21__2_), .S(n3097), .Z(n4802) );
  INV_X4 U6229 ( .A(n4802), .ZN(n4805) );
  MUX2_X2 U6230 ( .A(mem_22__2_), .B(mem_23__2_), .S(n3097), .Z(n4803) );
  INV_X4 U6231 ( .A(n4803), .ZN(n4804) );
  MUX2_X2 U6232 ( .A(n4805), .B(n4804), .S(n3081), .Z(n4806) );
  NAND3_X2 U6233 ( .A1(n4806), .A2(n2335), .A3(n2366), .ZN(n4813) );
  MUX2_X2 U6234 ( .A(mem_8__2_), .B(mem_9__2_), .S(n3097), .Z(n4807) );
  INV_X4 U6235 ( .A(n4807), .ZN(n4810) );
  MUX2_X2 U6236 ( .A(mem_10__2_), .B(mem_11__2_), .S(n3097), .Z(n4808) );
  INV_X4 U6237 ( .A(n4808), .ZN(n4809) );
  MUX2_X2 U6238 ( .A(n4810), .B(n4809), .S(n3081), .Z(n4811) );
  NAND3_X2 U6239 ( .A1(n4811), .A2(n2340), .A3(n2367), .ZN(n4812) );
  NAND4_X2 U6240 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4824)
         );
  MUX2_X2 U6241 ( .A(mem_0__2_), .B(mem_1__2_), .S(n3097), .Z(n4817) );
  MUX2_X2 U6242 ( .A(mem_2__2_), .B(mem_3__2_), .S(n3097), .Z(n4816) );
  MUX2_X2 U6243 ( .A(n4817), .B(n4816), .S(n3081), .Z(n4818) );
  NAND3_X2 U6244 ( .A1(n4818), .A2(n2344), .A3(n2368), .ZN(n4823) );
  MUX2_X2 U6245 ( .A(mem_4__2_), .B(mem_5__2_), .S(n3097), .Z(n4820) );
  MUX2_X2 U6246 ( .A(mem_6__2_), .B(mem_7__2_), .S(n3097), .Z(n4819) );
  MUX2_X2 U6247 ( .A(n4820), .B(n4819), .S(n3081), .Z(n4821) );
  NAND3_X2 U6248 ( .A1(n4821), .A2(n2342), .A3(n2369), .ZN(n4822) );
  OAI211_X2 U6249 ( .C1(n4825), .C2(n4824), .A(n4823), .B(n4822), .ZN(n7224)
         );
  MUX2_X2 U6250 ( .A(mem_28__3_), .B(mem_29__3_), .S(n3096), .Z(n4826) );
  INV_X4 U6251 ( .A(n4826), .ZN(n4829) );
  MUX2_X2 U6252 ( .A(mem_30__3_), .B(mem_31__3_), .S(n3096), .Z(n4827) );
  INV_X4 U6253 ( .A(n4827), .ZN(n4828) );
  MUX2_X2 U6254 ( .A(n4829), .B(n4828), .S(n3081), .Z(n4830) );
  NAND4_X2 U6255 ( .A1(n4830), .A2(n2334), .A3(n3061), .A4(n2374), .ZN(n4839)
         );
  MUX2_X2 U6256 ( .A(mem_24__3_), .B(mem_25__3_), .S(n3096), .Z(n4831) );
  INV_X4 U6257 ( .A(n4831), .ZN(n4834) );
  MUX2_X2 U6258 ( .A(mem_26__3_), .B(mem_27__3_), .S(n3096), .Z(n4832) );
  INV_X4 U6259 ( .A(n4832), .ZN(n4833) );
  MUX2_X2 U6260 ( .A(n4834), .B(n4833), .S(n3081), .Z(n4835) );
  NAND4_X2 U6261 ( .A1(n4835), .A2(n2343), .A3(n3061), .A4(n2503), .ZN(n4838)
         );
  NAND3_X2 U6262 ( .A1(n4839), .A2(n4838), .A3(n4837), .ZN(n4873) );
  MUX2_X2 U6263 ( .A(mem_12__3_), .B(mem_13__3_), .S(n3096), .Z(n4840) );
  INV_X4 U6264 ( .A(n4840), .ZN(n4843) );
  MUX2_X2 U6265 ( .A(mem_14__3_), .B(mem_15__3_), .S(n3096), .Z(n4841) );
  INV_X4 U6266 ( .A(n4841), .ZN(n4842) );
  MUX2_X2 U6267 ( .A(n4843), .B(n4842), .S(n3081), .Z(n4844) );
  NAND3_X2 U6268 ( .A1(n4844), .A2(n2346), .A3(n2504), .ZN(n4863) );
  MUX2_X2 U6269 ( .A(mem_16__3_), .B(mem_17__3_), .S(n3096), .Z(n4845) );
  INV_X4 U6270 ( .A(n4845), .ZN(n4848) );
  MUX2_X2 U6271 ( .A(mem_18__3_), .B(mem_19__3_), .S(n3096), .Z(n4846) );
  INV_X4 U6272 ( .A(n4846), .ZN(n4847) );
  MUX2_X2 U6273 ( .A(n4848), .B(n4847), .S(n3080), .Z(n4849) );
  NAND3_X2 U6274 ( .A1(n4849), .A2(n2332), .A3(n2364), .ZN(n4862) );
  MUX2_X2 U6275 ( .A(mem_20__3_), .B(mem_21__3_), .S(n3096), .Z(n4850) );
  INV_X4 U6276 ( .A(n4850), .ZN(n4853) );
  MUX2_X2 U6277 ( .A(mem_22__3_), .B(mem_23__3_), .S(n3096), .Z(n4851) );
  INV_X4 U6278 ( .A(n4851), .ZN(n4852) );
  MUX2_X2 U6279 ( .A(n4853), .B(n4852), .S(n3081), .Z(n4854) );
  NAND3_X2 U6280 ( .A1(n4854), .A2(n2336), .A3(n2366), .ZN(n4861) );
  MUX2_X2 U6281 ( .A(mem_8__3_), .B(mem_9__3_), .S(n3096), .Z(n4855) );
  INV_X4 U6282 ( .A(n4855), .ZN(n4858) );
  MUX2_X2 U6283 ( .A(mem_10__3_), .B(mem_11__3_), .S(n3096), .Z(n4856) );
  INV_X4 U6284 ( .A(n4856), .ZN(n4857) );
  MUX2_X2 U6285 ( .A(n4858), .B(n4857), .S(n3081), .Z(n4859) );
  NAND3_X2 U6286 ( .A1(n4859), .A2(n2341), .A3(n2367), .ZN(n4860) );
  NAND4_X2 U6287 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n4872)
         );
  MUX2_X2 U6288 ( .A(mem_0__3_), .B(mem_1__3_), .S(n3096), .Z(n4865) );
  MUX2_X2 U6289 ( .A(mem_2__3_), .B(mem_3__3_), .S(n3096), .Z(n4864) );
  MUX2_X2 U6290 ( .A(n4865), .B(n4864), .S(n3080), .Z(n4866) );
  NAND3_X2 U6291 ( .A1(n4866), .A2(n2345), .A3(n2368), .ZN(n4871) );
  MUX2_X2 U6292 ( .A(mem_4__3_), .B(mem_5__3_), .S(n3096), .Z(n4868) );
  MUX2_X2 U6293 ( .A(mem_6__3_), .B(mem_7__3_), .S(n3096), .Z(n4867) );
  MUX2_X2 U6294 ( .A(n4868), .B(n4867), .S(n3080), .Z(n4869) );
  NAND3_X2 U6295 ( .A1(n4869), .A2(n2341), .A3(n2369), .ZN(n4870) );
  OAI211_X2 U6296 ( .C1(n4873), .C2(n4872), .A(n4871), .B(n4870), .ZN(n7223)
         );
  MUX2_X2 U6297 ( .A(mem_28__4_), .B(mem_29__4_), .S(n3096), .Z(n4874) );
  INV_X4 U6298 ( .A(n4874), .ZN(n4877) );
  MUX2_X2 U6299 ( .A(mem_30__4_), .B(mem_31__4_), .S(n3096), .Z(n4875) );
  INV_X4 U6300 ( .A(n4875), .ZN(n4876) );
  MUX2_X2 U6301 ( .A(n4877), .B(n4876), .S(n3080), .Z(n4878) );
  NAND4_X2 U6302 ( .A1(n4878), .A2(n2331), .A3(n3061), .A4(n2374), .ZN(n4887)
         );
  MUX2_X2 U6303 ( .A(mem_24__4_), .B(mem_25__4_), .S(n3096), .Z(n4879) );
  INV_X4 U6304 ( .A(n4879), .ZN(n4882) );
  MUX2_X2 U6305 ( .A(mem_26__4_), .B(mem_27__4_), .S(n3096), .Z(n4880) );
  INV_X4 U6306 ( .A(n4880), .ZN(n4881) );
  MUX2_X2 U6307 ( .A(n4882), .B(n4881), .S(n3080), .Z(n4883) );
  NAND4_X2 U6308 ( .A1(n4883), .A2(n2343), .A3(n3061), .A4(n2503), .ZN(n4886)
         );
  NAND3_X2 U6309 ( .A1(n4887), .A2(n4886), .A3(n4885), .ZN(n4921) );
  MUX2_X2 U6310 ( .A(mem_12__4_), .B(mem_13__4_), .S(n3095), .Z(n4888) );
  INV_X4 U6311 ( .A(n4888), .ZN(n4891) );
  MUX2_X2 U6312 ( .A(mem_14__4_), .B(mem_15__4_), .S(n3095), .Z(n4889) );
  INV_X4 U6313 ( .A(n4889), .ZN(n4890) );
  MUX2_X2 U6314 ( .A(n4891), .B(n4890), .S(n3080), .Z(n4892) );
  NAND3_X2 U6315 ( .A1(n4892), .A2(n2337), .A3(n2504), .ZN(n4911) );
  MUX2_X2 U6316 ( .A(mem_16__4_), .B(mem_17__4_), .S(n3095), .Z(n4893) );
  INV_X4 U6317 ( .A(n4893), .ZN(n4896) );
  MUX2_X2 U6318 ( .A(mem_18__4_), .B(mem_19__4_), .S(n3095), .Z(n4894) );
  INV_X4 U6319 ( .A(n4894), .ZN(n4895) );
  MUX2_X2 U6320 ( .A(n4896), .B(n4895), .S(n3080), .Z(n4897) );
  NAND3_X2 U6321 ( .A1(n4897), .A2(n2346), .A3(n2364), .ZN(n4910) );
  MUX2_X2 U6322 ( .A(mem_20__4_), .B(mem_21__4_), .S(n3095), .Z(n4898) );
  INV_X4 U6323 ( .A(n4898), .ZN(n4901) );
  MUX2_X2 U6324 ( .A(mem_22__4_), .B(mem_23__4_), .S(n3095), .Z(n4899) );
  INV_X4 U6325 ( .A(n4899), .ZN(n4900) );
  MUX2_X2 U6326 ( .A(n4901), .B(n4900), .S(n3080), .Z(n4902) );
  NAND3_X2 U6327 ( .A1(n4902), .A2(n2331), .A3(n2366), .ZN(n4909) );
  MUX2_X2 U6328 ( .A(mem_8__4_), .B(mem_9__4_), .S(n3095), .Z(n4903) );
  INV_X4 U6329 ( .A(n4903), .ZN(n4906) );
  MUX2_X2 U6330 ( .A(mem_10__4_), .B(mem_11__4_), .S(n3095), .Z(n4904) );
  INV_X4 U6331 ( .A(n4904), .ZN(n4905) );
  MUX2_X2 U6332 ( .A(n4906), .B(n4905), .S(n3080), .Z(n4907) );
  NAND3_X2 U6333 ( .A1(n4907), .A2(n2327), .A3(n2367), .ZN(n4908) );
  NAND4_X2 U6334 ( .A1(n4911), .A2(n4910), .A3(n4909), .A4(n4908), .ZN(n4920)
         );
  MUX2_X2 U6335 ( .A(mem_0__4_), .B(mem_1__4_), .S(n3095), .Z(n4913) );
  MUX2_X2 U6336 ( .A(mem_2__4_), .B(mem_3__4_), .S(n3095), .Z(n4912) );
  MUX2_X2 U6337 ( .A(n4913), .B(n4912), .S(n3080), .Z(n4914) );
  NAND3_X2 U6338 ( .A1(n4914), .A2(n2338), .A3(n2368), .ZN(n4919) );
  MUX2_X2 U6339 ( .A(mem_4__4_), .B(mem_5__4_), .S(n3095), .Z(n4916) );
  MUX2_X2 U6340 ( .A(mem_6__4_), .B(mem_7__4_), .S(n3095), .Z(n4915) );
  MUX2_X2 U6341 ( .A(n4916), .B(n4915), .S(n3080), .Z(n4917) );
  NAND3_X2 U6342 ( .A1(n4917), .A2(n2340), .A3(n2369), .ZN(n4918) );
  OAI211_X2 U6343 ( .C1(n4921), .C2(n4920), .A(n4919), .B(n4918), .ZN(n7222)
         );
  MUX2_X2 U6344 ( .A(mem_28__5_), .B(mem_29__5_), .S(n3095), .Z(n4922) );
  INV_X4 U6345 ( .A(n4922), .ZN(n4925) );
  MUX2_X2 U6346 ( .A(mem_30__5_), .B(mem_31__5_), .S(n3095), .Z(n4923) );
  INV_X4 U6347 ( .A(n4923), .ZN(n4924) );
  MUX2_X2 U6348 ( .A(n4925), .B(n4924), .S(n3080), .Z(n4926) );
  NAND4_X2 U6349 ( .A1(n4926), .A2(n2327), .A3(n3061), .A4(n2374), .ZN(n4935)
         );
  MUX2_X2 U6350 ( .A(mem_24__5_), .B(mem_25__5_), .S(n3095), .Z(n4927) );
  INV_X4 U6351 ( .A(n4927), .ZN(n4930) );
  MUX2_X2 U6352 ( .A(mem_26__5_), .B(mem_27__5_), .S(n3095), .Z(n4928) );
  INV_X4 U6353 ( .A(n4928), .ZN(n4929) );
  MUX2_X2 U6354 ( .A(n4930), .B(n4929), .S(n3080), .Z(n4931) );
  NAND4_X2 U6355 ( .A1(n4931), .A2(n2337), .A3(n3061), .A4(n2503), .ZN(n4934)
         );
  NAND3_X2 U6356 ( .A1(n4935), .A2(n4934), .A3(n4933), .ZN(n4969) );
  MUX2_X2 U6357 ( .A(mem_12__5_), .B(mem_13__5_), .S(n3095), .Z(n4936) );
  INV_X4 U6358 ( .A(n4936), .ZN(n4939) );
  MUX2_X2 U6359 ( .A(mem_14__5_), .B(mem_15__5_), .S(n3095), .Z(n4937) );
  INV_X4 U6360 ( .A(n4937), .ZN(n4938) );
  MUX2_X2 U6361 ( .A(n4939), .B(n4938), .S(n3080), .Z(n4940) );
  NAND3_X2 U6362 ( .A1(n4940), .A2(n2338), .A3(n2504), .ZN(n4959) );
  MUX2_X2 U6363 ( .A(mem_16__5_), .B(mem_17__5_), .S(n3095), .Z(n4941) );
  INV_X4 U6364 ( .A(n4941), .ZN(n4944) );
  MUX2_X2 U6365 ( .A(mem_18__5_), .B(mem_19__5_), .S(n3095), .Z(n4942) );
  INV_X4 U6366 ( .A(n4942), .ZN(n4943) );
  MUX2_X2 U6367 ( .A(n4944), .B(n4943), .S(n3080), .Z(n4945) );
  NAND3_X2 U6368 ( .A1(n4945), .A2(n2329), .A3(n2364), .ZN(n4958) );
  MUX2_X2 U6369 ( .A(mem_20__5_), .B(mem_21__5_), .S(n3095), .Z(n4946) );
  INV_X4 U6370 ( .A(n4946), .ZN(n4949) );
  MUX2_X2 U6371 ( .A(mem_22__5_), .B(mem_23__5_), .S(n3102), .Z(n4947) );
  INV_X4 U6372 ( .A(n4947), .ZN(n4948) );
  MUX2_X2 U6373 ( .A(n4949), .B(n4948), .S(n3079), .Z(n4950) );
  NAND3_X2 U6374 ( .A1(n4950), .A2(n2332), .A3(n2366), .ZN(n4957) );
  MUX2_X2 U6375 ( .A(mem_8__5_), .B(mem_9__5_), .S(n3102), .Z(n4951) );
  INV_X4 U6376 ( .A(n4951), .ZN(n4954) );
  MUX2_X2 U6377 ( .A(mem_10__5_), .B(mem_11__5_), .S(n3101), .Z(n4952) );
  INV_X4 U6378 ( .A(n4952), .ZN(n4953) );
  MUX2_X2 U6379 ( .A(n4954), .B(n4953), .S(n3080), .Z(n4955) );
  NAND3_X2 U6380 ( .A1(n4955), .A2(n2345), .A3(n2367), .ZN(n4956) );
  NAND4_X2 U6381 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4968)
         );
  MUX2_X2 U6382 ( .A(mem_0__5_), .B(mem_1__5_), .S(n3101), .Z(n4961) );
  MUX2_X2 U6383 ( .A(mem_2__5_), .B(mem_3__5_), .S(n3101), .Z(n4960) );
  MUX2_X2 U6384 ( .A(n4961), .B(n4960), .S(n3079), .Z(n4962) );
  NAND3_X2 U6385 ( .A1(n4962), .A2(n2337), .A3(n2368), .ZN(n4967) );
  MUX2_X2 U6386 ( .A(mem_4__5_), .B(mem_5__5_), .S(n3102), .Z(n4964) );
  MUX2_X2 U6387 ( .A(mem_6__5_), .B(mem_7__5_), .S(n3101), .Z(n4963) );
  MUX2_X2 U6388 ( .A(n4964), .B(n4963), .S(n3079), .Z(n4965) );
  NAND3_X2 U6389 ( .A1(n4965), .A2(n2341), .A3(n2369), .ZN(n4966) );
  OAI211_X2 U6390 ( .C1(n4969), .C2(n4968), .A(n4967), .B(n4966), .ZN(n7221)
         );
  MUX2_X2 U6391 ( .A(mem_28__6_), .B(mem_29__6_), .S(n3102), .Z(n4970) );
  INV_X4 U6392 ( .A(n4970), .ZN(n4973) );
  MUX2_X2 U6393 ( .A(mem_30__6_), .B(mem_31__6_), .S(n3102), .Z(n4971) );
  INV_X4 U6394 ( .A(n4971), .ZN(n4972) );
  MUX2_X2 U6395 ( .A(n4973), .B(n4972), .S(n3079), .Z(n4974) );
  NAND4_X2 U6396 ( .A1(n4974), .A2(n2341), .A3(n3061), .A4(n2374), .ZN(n4983)
         );
  MUX2_X2 U6397 ( .A(mem_24__6_), .B(mem_25__6_), .S(n3098), .Z(n4975) );
  INV_X4 U6398 ( .A(n4975), .ZN(n4978) );
  MUX2_X2 U6399 ( .A(mem_26__6_), .B(mem_27__6_), .S(n3101), .Z(n4976) );
  INV_X4 U6400 ( .A(n4976), .ZN(n4977) );
  MUX2_X2 U6401 ( .A(n4978), .B(n4977), .S(n3079), .Z(n4979) );
  NAND4_X2 U6402 ( .A1(n4979), .A2(n2338), .A3(n3061), .A4(n2503), .ZN(n4982)
         );
  NAND3_X2 U6403 ( .A1(n4983), .A2(n4982), .A3(n4981), .ZN(n5017) );
  MUX2_X2 U6404 ( .A(mem_12__6_), .B(mem_13__6_), .S(n3096), .Z(n4984) );
  INV_X4 U6405 ( .A(n4984), .ZN(n4987) );
  MUX2_X2 U6406 ( .A(mem_14__6_), .B(mem_15__6_), .S(n3103), .Z(n4985) );
  INV_X4 U6407 ( .A(n4985), .ZN(n4986) );
  MUX2_X2 U6408 ( .A(n4987), .B(n4986), .S(n3079), .Z(n4988) );
  NAND3_X2 U6409 ( .A1(n4988), .A2(n2334), .A3(n2504), .ZN(n5007) );
  MUX2_X2 U6410 ( .A(mem_16__6_), .B(mem_17__6_), .S(n3103), .Z(n4989) );
  INV_X4 U6411 ( .A(n4989), .ZN(n4992) );
  MUX2_X2 U6412 ( .A(mem_18__6_), .B(mem_19__6_), .S(n3103), .Z(n4990) );
  INV_X4 U6413 ( .A(n4990), .ZN(n4991) );
  MUX2_X2 U6414 ( .A(n4992), .B(n4991), .S(n3079), .Z(n4993) );
  NAND3_X2 U6415 ( .A1(n4993), .A2(n2331), .A3(n2364), .ZN(n5006) );
  MUX2_X2 U6416 ( .A(mem_20__6_), .B(mem_21__6_), .S(n3103), .Z(n4994) );
  INV_X4 U6417 ( .A(n4994), .ZN(n4997) );
  MUX2_X2 U6418 ( .A(mem_22__6_), .B(mem_23__6_), .S(n3103), .Z(n4995) );
  INV_X4 U6419 ( .A(n4995), .ZN(n4996) );
  MUX2_X2 U6420 ( .A(n4997), .B(n4996), .S(n3079), .Z(n4998) );
  NAND3_X2 U6421 ( .A1(n4998), .A2(n2333), .A3(n2366), .ZN(n5005) );
  MUX2_X2 U6422 ( .A(mem_8__6_), .B(mem_9__6_), .S(n3103), .Z(n4999) );
  INV_X4 U6423 ( .A(n4999), .ZN(n5002) );
  MUX2_X2 U6424 ( .A(mem_10__6_), .B(mem_11__6_), .S(n3103), .Z(n5000) );
  INV_X4 U6425 ( .A(n5000), .ZN(n5001) );
  MUX2_X2 U6426 ( .A(n5002), .B(n5001), .S(n3079), .Z(n5003) );
  NAND3_X2 U6427 ( .A1(n5003), .A2(n2344), .A3(n2367), .ZN(n5004) );
  NAND4_X2 U6428 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5016)
         );
  MUX2_X2 U6429 ( .A(mem_0__6_), .B(mem_1__6_), .S(n3103), .Z(n5009) );
  MUX2_X2 U6430 ( .A(mem_2__6_), .B(mem_3__6_), .S(n3103), .Z(n5008) );
  MUX2_X2 U6431 ( .A(n5009), .B(n5008), .S(n3079), .Z(n5010) );
  NAND3_X2 U6432 ( .A1(n5010), .A2(n2336), .A3(n2368), .ZN(n5015) );
  MUX2_X2 U6433 ( .A(mem_4__6_), .B(mem_5__6_), .S(n3103), .Z(n5012) );
  MUX2_X2 U6434 ( .A(mem_6__6_), .B(mem_7__6_), .S(n3103), .Z(n5011) );
  MUX2_X2 U6435 ( .A(n5012), .B(n5011), .S(n3079), .Z(n5013) );
  NAND3_X2 U6436 ( .A1(n5013), .A2(n2342), .A3(n2369), .ZN(n5014) );
  OAI211_X2 U6437 ( .C1(n5017), .C2(n5016), .A(n5015), .B(n5014), .ZN(n7220)
         );
  MUX2_X2 U6438 ( .A(mem_28__7_), .B(mem_29__7_), .S(n3103), .Z(n5018) );
  INV_X4 U6439 ( .A(n5018), .ZN(n5021) );
  MUX2_X2 U6440 ( .A(mem_30__7_), .B(mem_31__7_), .S(n3103), .Z(n5019) );
  INV_X4 U6441 ( .A(n5019), .ZN(n5020) );
  MUX2_X2 U6442 ( .A(n5021), .B(n5020), .S(n3079), .Z(n5022) );
  NAND4_X2 U6443 ( .A1(n5022), .A2(n2345), .A3(n3061), .A4(n2374), .ZN(n5031)
         );
  MUX2_X2 U6444 ( .A(mem_24__7_), .B(mem_25__7_), .S(n3103), .Z(n5023) );
  INV_X4 U6445 ( .A(n5023), .ZN(n5026) );
  MUX2_X2 U6446 ( .A(mem_26__7_), .B(mem_27__7_), .S(n3103), .Z(n5024) );
  INV_X4 U6447 ( .A(n5024), .ZN(n5025) );
  MUX2_X2 U6448 ( .A(n5026), .B(n5025), .S(n3079), .Z(n5027) );
  NAND4_X2 U6449 ( .A1(n5027), .A2(n2338), .A3(n3061), .A4(n2503), .ZN(n5030)
         );
  NAND3_X2 U6450 ( .A1(n5031), .A2(n5030), .A3(n5029), .ZN(n5065) );
  MUX2_X2 U6451 ( .A(mem_12__7_), .B(mem_13__7_), .S(n3103), .Z(n5032) );
  INV_X4 U6452 ( .A(n5032), .ZN(n5035) );
  MUX2_X2 U6453 ( .A(mem_14__7_), .B(mem_15__7_), .S(n3102), .Z(n5033) );
  INV_X4 U6454 ( .A(n5033), .ZN(n5034) );
  MUX2_X2 U6455 ( .A(n5035), .B(n5034), .S(n3079), .Z(n5036) );
  NAND3_X2 U6456 ( .A1(n5036), .A2(n2338), .A3(n2504), .ZN(n5055) );
  MUX2_X2 U6457 ( .A(mem_16__7_), .B(mem_17__7_), .S(n3103), .Z(n5037) );
  INV_X4 U6458 ( .A(n5037), .ZN(n5040) );
  MUX2_X2 U6459 ( .A(mem_18__7_), .B(mem_19__7_), .S(n3103), .Z(n5038) );
  INV_X4 U6460 ( .A(n5038), .ZN(n5039) );
  MUX2_X2 U6461 ( .A(n5040), .B(n5039), .S(n3078), .Z(n5041) );
  NAND3_X2 U6462 ( .A1(n5041), .A2(n2333), .A3(n2364), .ZN(n5054) );
  MUX2_X2 U6463 ( .A(mem_20__7_), .B(mem_21__7_), .S(n3103), .Z(n5042) );
  INV_X4 U6464 ( .A(n5042), .ZN(n5045) );
  MUX2_X2 U6465 ( .A(mem_22__7_), .B(mem_23__7_), .S(n3102), .Z(n5043) );
  INV_X4 U6466 ( .A(n5043), .ZN(n5044) );
  MUX2_X2 U6467 ( .A(n5045), .B(n5044), .S(n3079), .Z(n5046) );
  NAND3_X2 U6468 ( .A1(n5046), .A2(n2341), .A3(n2366), .ZN(n5053) );
  MUX2_X2 U6469 ( .A(mem_8__7_), .B(mem_9__7_), .S(n3102), .Z(n5047) );
  INV_X4 U6470 ( .A(n5047), .ZN(n5050) );
  MUX2_X2 U6471 ( .A(mem_10__7_), .B(mem_11__7_), .S(n3102), .Z(n5048) );
  INV_X4 U6472 ( .A(n5048), .ZN(n5049) );
  MUX2_X2 U6473 ( .A(n5050), .B(n5049), .S(n3079), .Z(n5051) );
  NAND3_X2 U6474 ( .A1(n5051), .A2(n2328), .A3(n2367), .ZN(n5052) );
  NAND4_X2 U6475 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n5064)
         );
  MUX2_X2 U6476 ( .A(mem_0__7_), .B(mem_1__7_), .S(n3102), .Z(n5057) );
  MUX2_X2 U6477 ( .A(mem_2__7_), .B(mem_3__7_), .S(n3102), .Z(n5056) );
  MUX2_X2 U6478 ( .A(n5057), .B(n5056), .S(n3078), .Z(n5058) );
  NAND3_X2 U6479 ( .A1(n5058), .A2(n2335), .A3(n2368), .ZN(n5063) );
  MUX2_X2 U6480 ( .A(mem_4__7_), .B(mem_5__7_), .S(n3102), .Z(n5060) );
  MUX2_X2 U6481 ( .A(mem_6__7_), .B(mem_7__7_), .S(n3102), .Z(n5059) );
  MUX2_X2 U6482 ( .A(n5060), .B(n5059), .S(n3078), .Z(n5061) );
  NAND3_X2 U6483 ( .A1(n5061), .A2(n2342), .A3(n2369), .ZN(n5062) );
  OAI211_X2 U6484 ( .C1(n5065), .C2(n5064), .A(n5063), .B(n5062), .ZN(n7219)
         );
  MUX2_X2 U6485 ( .A(mem_28__8_), .B(mem_29__8_), .S(n3102), .Z(n5066) );
  INV_X4 U6486 ( .A(n5066), .ZN(n5069) );
  MUX2_X2 U6487 ( .A(mem_30__8_), .B(mem_31__8_), .S(n3102), .Z(n5067) );
  INV_X4 U6488 ( .A(n5067), .ZN(n5068) );
  MUX2_X2 U6489 ( .A(n5069), .B(n5068), .S(n3078), .Z(n5070) );
  NAND4_X2 U6490 ( .A1(n5070), .A2(n2336), .A3(n3061), .A4(n2374), .ZN(n5079)
         );
  MUX2_X2 U6491 ( .A(mem_24__8_), .B(mem_25__8_), .S(n3102), .Z(n5071) );
  INV_X4 U6492 ( .A(n5071), .ZN(n5074) );
  MUX2_X2 U6493 ( .A(mem_26__8_), .B(mem_27__8_), .S(n3102), .Z(n5072) );
  INV_X4 U6494 ( .A(n5072), .ZN(n5073) );
  MUX2_X2 U6495 ( .A(n5074), .B(n5073), .S(n3078), .Z(n5075) );
  NAND4_X2 U6496 ( .A1(n5075), .A2(n2339), .A3(n3061), .A4(n2503), .ZN(n5078)
         );
  NAND3_X2 U6497 ( .A1(n5079), .A2(n5078), .A3(n5077), .ZN(n5113) );
  MUX2_X2 U6498 ( .A(mem_12__8_), .B(mem_13__8_), .S(n3102), .Z(n5080) );
  INV_X4 U6499 ( .A(n5080), .ZN(n5083) );
  MUX2_X2 U6500 ( .A(mem_14__8_), .B(mem_15__8_), .S(n3102), .Z(n5081) );
  INV_X4 U6501 ( .A(n5081), .ZN(n5082) );
  MUX2_X2 U6502 ( .A(n5083), .B(n5082), .S(n3078), .Z(n5084) );
  NAND3_X2 U6503 ( .A1(n5084), .A2(n2339), .A3(n2504), .ZN(n5103) );
  MUX2_X2 U6504 ( .A(mem_16__8_), .B(mem_17__8_), .S(n3102), .Z(n5085) );
  INV_X4 U6505 ( .A(n5085), .ZN(n5088) );
  MUX2_X2 U6506 ( .A(mem_18__8_), .B(mem_19__8_), .S(n3102), .Z(n5086) );
  INV_X4 U6507 ( .A(n5086), .ZN(n5087) );
  MUX2_X2 U6508 ( .A(n5088), .B(n5087), .S(n3078), .Z(n5089) );
  NAND3_X2 U6509 ( .A1(n5089), .A2(n2334), .A3(n2364), .ZN(n5102) );
  MUX2_X2 U6510 ( .A(mem_20__8_), .B(mem_21__8_), .S(n3102), .Z(n5090) );
  INV_X4 U6511 ( .A(n5090), .ZN(n5093) );
  MUX2_X2 U6512 ( .A(mem_22__8_), .B(mem_23__8_), .S(n3102), .Z(n5091) );
  INV_X4 U6513 ( .A(n5091), .ZN(n5092) );
  MUX2_X2 U6514 ( .A(n5093), .B(n5092), .S(n3078), .Z(n5094) );
  NAND3_X2 U6515 ( .A1(n5094), .A2(n2329), .A3(n2366), .ZN(n5101) );
  MUX2_X2 U6516 ( .A(mem_8__8_), .B(mem_9__8_), .S(n3101), .Z(n5095) );
  INV_X4 U6517 ( .A(n5095), .ZN(n5098) );
  MUX2_X2 U6518 ( .A(mem_10__8_), .B(mem_11__8_), .S(n3102), .Z(n5096) );
  INV_X4 U6519 ( .A(n5096), .ZN(n5097) );
  MUX2_X2 U6520 ( .A(n5098), .B(n5097), .S(n3078), .Z(n5099) );
  NAND3_X2 U6521 ( .A1(n5099), .A2(n2333), .A3(n2367), .ZN(n5100) );
  NAND4_X2 U6522 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n5112)
         );
  MUX2_X2 U6523 ( .A(mem_0__8_), .B(mem_1__8_), .S(n3102), .Z(n5105) );
  MUX2_X2 U6524 ( .A(mem_2__8_), .B(mem_3__8_), .S(n3102), .Z(n5104) );
  MUX2_X2 U6525 ( .A(n5105), .B(n5104), .S(n3078), .Z(n5106) );
  NAND3_X2 U6526 ( .A1(n5106), .A2(n2336), .A3(n2368), .ZN(n5111) );
  MUX2_X2 U6527 ( .A(mem_4__8_), .B(mem_5__8_), .S(n3101), .Z(n5108) );
  MUX2_X2 U6528 ( .A(mem_6__8_), .B(mem_7__8_), .S(n3101), .Z(n5107) );
  MUX2_X2 U6529 ( .A(n5108), .B(n5107), .S(n3078), .Z(n5109) );
  NAND3_X2 U6530 ( .A1(n5109), .A2(n2341), .A3(n2369), .ZN(n5110) );
  OAI211_X2 U6531 ( .C1(n5113), .C2(n5112), .A(n5111), .B(n5110), .ZN(n7218)
         );
  MUX2_X2 U6532 ( .A(mem_28__9_), .B(mem_29__9_), .S(n3101), .Z(n5114) );
  INV_X4 U6533 ( .A(n5114), .ZN(n5117) );
  MUX2_X2 U6534 ( .A(mem_30__9_), .B(mem_31__9_), .S(n3101), .Z(n5115) );
  INV_X4 U6535 ( .A(n5115), .ZN(n5116) );
  MUX2_X2 U6536 ( .A(n5117), .B(n5116), .S(n3078), .Z(n5118) );
  NAND4_X2 U6537 ( .A1(n5118), .A2(n2346), .A3(n3061), .A4(n2374), .ZN(n5127)
         );
  MUX2_X2 U6538 ( .A(mem_24__9_), .B(mem_25__9_), .S(n3101), .Z(n5119) );
  INV_X4 U6539 ( .A(n5119), .ZN(n5122) );
  MUX2_X2 U6540 ( .A(mem_26__9_), .B(mem_27__9_), .S(n3101), .Z(n5120) );
  INV_X4 U6541 ( .A(n5120), .ZN(n5121) );
  MUX2_X2 U6542 ( .A(n5122), .B(n5121), .S(n3078), .Z(n5123) );
  NAND4_X2 U6543 ( .A1(n5123), .A2(n2330), .A3(n3061), .A4(n2503), .ZN(n5126)
         );
  NAND3_X2 U6544 ( .A1(n5127), .A2(n5126), .A3(n5125), .ZN(n5161) );
  MUX2_X2 U6545 ( .A(mem_12__9_), .B(mem_13__9_), .S(n3101), .Z(n5128) );
  INV_X4 U6546 ( .A(n5128), .ZN(n5131) );
  MUX2_X2 U6547 ( .A(mem_14__9_), .B(mem_15__9_), .S(n3101), .Z(n5129) );
  INV_X4 U6548 ( .A(n5129), .ZN(n5130) );
  MUX2_X2 U6549 ( .A(n5131), .B(n5130), .S(n3078), .Z(n5132) );
  NAND3_X2 U6550 ( .A1(n5132), .A2(n2340), .A3(n2504), .ZN(n5151) );
  MUX2_X2 U6551 ( .A(mem_16__9_), .B(mem_17__9_), .S(n3101), .Z(n5133) );
  INV_X4 U6552 ( .A(n5133), .ZN(n5136) );
  MUX2_X2 U6553 ( .A(mem_18__9_), .B(mem_19__9_), .S(n3101), .Z(n5134) );
  INV_X4 U6554 ( .A(n5134), .ZN(n5135) );
  MUX2_X2 U6555 ( .A(n5136), .B(n5135), .S(n3078), .Z(n5137) );
  NAND3_X2 U6556 ( .A1(n5137), .A2(n2335), .A3(n2364), .ZN(n5150) );
  MUX2_X2 U6557 ( .A(mem_20__9_), .B(mem_21__9_), .S(n3101), .Z(n5138) );
  INV_X4 U6558 ( .A(n5138), .ZN(n5141) );
  MUX2_X2 U6559 ( .A(mem_22__9_), .B(mem_23__9_), .S(n3101), .Z(n5139) );
  INV_X4 U6560 ( .A(n5139), .ZN(n5140) );
  MUX2_X2 U6561 ( .A(n5141), .B(n5140), .S(n3078), .Z(n5142) );
  NAND3_X2 U6562 ( .A1(n5142), .A2(n2330), .A3(n2366), .ZN(n5149) );
  MUX2_X2 U6563 ( .A(mem_8__9_), .B(mem_9__9_), .S(n3101), .Z(n5143) );
  INV_X4 U6564 ( .A(n5143), .ZN(n5146) );
  MUX2_X2 U6565 ( .A(mem_10__9_), .B(mem_11__9_), .S(n3101), .Z(n5144) );
  INV_X4 U6566 ( .A(n5144), .ZN(n5145) );
  MUX2_X2 U6567 ( .A(n5146), .B(n5145), .S(n3077), .Z(n5147) );
  NAND3_X2 U6568 ( .A1(n5147), .A2(n2334), .A3(n2367), .ZN(n5148) );
  NAND4_X2 U6569 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n5160)
         );
  MUX2_X2 U6570 ( .A(mem_0__9_), .B(mem_1__9_), .S(n3101), .Z(n5153) );
  MUX2_X2 U6571 ( .A(mem_2__9_), .B(mem_3__9_), .S(n3101), .Z(n5152) );
  MUX2_X2 U6572 ( .A(n5153), .B(n5152), .S(n3077), .Z(n5154) );
  NAND3_X2 U6573 ( .A1(n5154), .A2(n2345), .A3(n2368), .ZN(n5159) );
  MUX2_X2 U6574 ( .A(mem_4__9_), .B(mem_5__9_), .S(n3101), .Z(n5156) );
  MUX2_X2 U6575 ( .A(mem_6__9_), .B(mem_7__9_), .S(n3101), .Z(n5155) );
  MUX2_X2 U6576 ( .A(n5156), .B(n5155), .S(n3080), .Z(n5157) );
  NAND3_X2 U6577 ( .A1(n5157), .A2(n2343), .A3(n2369), .ZN(n5158) );
  OAI211_X2 U6578 ( .C1(n5161), .C2(n5160), .A(n5159), .B(n5158), .ZN(n7217)
         );
  MUX2_X2 U6579 ( .A(mem_8__10_), .B(mem_9__10_), .S(n3101), .Z(n5162) );
  NAND2_X2 U6580 ( .A1(n5163), .A2(n3062), .ZN(n5170) );
  MUX2_X2 U6581 ( .A(mem_14__10_), .B(mem_15__10_), .S(n3100), .Z(n5164) );
  NAND2_X2 U6582 ( .A1(n5165), .A2(n3062), .ZN(n5169) );
  MUX2_X2 U6583 ( .A(mem_10__10_), .B(mem_11__10_), .S(n3100), .Z(n5166) );
  NAND2_X2 U6584 ( .A1(n3081), .A2(n3070), .ZN(n5746) );
  NAND2_X2 U6585 ( .A1(n5167), .A2(n3062), .ZN(n5168) );
  NAND3_X2 U6586 ( .A1(n5170), .A2(n5169), .A3(n5168), .ZN(n5211) );
  MUX2_X2 U6587 ( .A(mem_30__10_), .B(mem_31__10_), .S(n3100), .Z(n5171) );
  NAND3_X2 U6588 ( .A1(n3063), .A2(n5171), .A3(n5798), .ZN(n5174) );
  MUX2_X2 U6589 ( .A(mem_28__10_), .B(mem_29__10_), .S(n3100), .Z(n5172) );
  NAND2_X2 U6590 ( .A1(n3067), .A2(n3084), .ZN(n5743) );
  INV_X4 U6591 ( .A(n5743), .ZN(n5756) );
  NAND3_X2 U6592 ( .A1(n3063), .A2(n5172), .A3(n5756), .ZN(n5173) );
  OAI22_X2 U6593 ( .A1(n3060), .A2(n3063), .B1(n2364), .B2(n3062), .ZN(n5758)
         );
  NAND3_X2 U6594 ( .A1(n5174), .A2(n5173), .A3(n5758), .ZN(n5192) );
  MUX2_X2 U6595 ( .A(mem_22__10_), .B(mem_23__10_), .S(n3100), .Z(n5175) );
  NAND3_X2 U6596 ( .A1(n3059), .A2(n5175), .A3(n2382), .ZN(n5182) );
  MUX2_X2 U6597 ( .A(mem_24__10_), .B(mem_25__10_), .S(n3100), .Z(n5176) );
  NAND3_X2 U6598 ( .A1(n3063), .A2(n5176), .A3(n2861), .ZN(n5181) );
  MUX2_X2 U6599 ( .A(mem_26__10_), .B(mem_27__10_), .S(n3100), .Z(n5177) );
  INV_X4 U6600 ( .A(n5746), .ZN(n5763) );
  NAND3_X2 U6601 ( .A1(n3063), .A2(n5177), .A3(n5763), .ZN(n5180) );
  MUX2_X2 U6602 ( .A(mem_20__10_), .B(mem_21__10_), .S(n3100), .Z(n5178) );
  NAND3_X2 U6603 ( .A1(n3061), .A2(n5178), .A3(n5765), .ZN(n5179) );
  NAND4_X2 U6604 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n5191)
         );
  MUX2_X2 U6605 ( .A(mem_16__10_), .B(mem_17__10_), .S(n3100), .Z(n5183) );
  NAND2_X2 U6606 ( .A1(n5184), .A2(n3064), .ZN(n5190) );
  MUX2_X2 U6607 ( .A(mem_18__10_), .B(mem_19__10_), .S(n3100), .Z(n5185) );
  MUX2_X2 U6608 ( .A(mem_12__10_), .B(mem_13__10_), .S(n3100), .Z(n5186) );
  OAI211_X2 U6609 ( .C1(n5192), .C2(n5191), .A(n5190), .B(n5189), .ZN(n5210)
         );
  NAND2_X2 U6610 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  NAND4_X2 U6611 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n5206)
         );
  NAND3_X2 U6612 ( .A1(n5207), .A2(n5206), .A3(n5205), .ZN(n5208) );
  NAND3_X2 U6613 ( .A1(n5208), .A2(n3064), .A3(n3062), .ZN(n5209) );
  MUX2_X2 U6614 ( .A(n5212), .B(wData[10]), .S(n2347), .Z(n7216) );
  MUX2_X2 U6615 ( .A(mem_28__11_), .B(mem_29__11_), .S(n3100), .Z(n5213) );
  INV_X4 U6616 ( .A(n5213), .ZN(n5216) );
  MUX2_X2 U6617 ( .A(mem_30__11_), .B(mem_31__11_), .S(n3100), .Z(n5214) );
  INV_X4 U6618 ( .A(n5214), .ZN(n5215) );
  MUX2_X2 U6619 ( .A(n5216), .B(n5215), .S(n3080), .Z(n5217) );
  NAND4_X2 U6620 ( .A1(n5217), .A2(n2342), .A3(n3060), .A4(n2374), .ZN(n5226)
         );
  MUX2_X2 U6621 ( .A(mem_24__11_), .B(mem_25__11_), .S(n3100), .Z(n5218) );
  INV_X4 U6622 ( .A(n5218), .ZN(n5221) );
  MUX2_X2 U6623 ( .A(mem_26__11_), .B(mem_27__11_), .S(n3100), .Z(n5219) );
  INV_X4 U6624 ( .A(n5219), .ZN(n5220) );
  MUX2_X2 U6625 ( .A(n5221), .B(n5220), .S(n3077), .Z(n5222) );
  NAND4_X2 U6626 ( .A1(n5222), .A2(n2335), .A3(n3060), .A4(n2503), .ZN(n5225)
         );
  NAND3_X2 U6627 ( .A1(n5226), .A2(n5225), .A3(n5224), .ZN(n5260) );
  MUX2_X2 U6628 ( .A(mem_12__11_), .B(mem_13__11_), .S(n3100), .Z(n5227) );
  INV_X4 U6629 ( .A(n5227), .ZN(n5230) );
  MUX2_X2 U6630 ( .A(mem_14__11_), .B(mem_15__11_), .S(n3100), .Z(n5228) );
  INV_X4 U6631 ( .A(n5228), .ZN(n5229) );
  MUX2_X2 U6632 ( .A(n5230), .B(n5229), .S(n3079), .Z(n5231) );
  NAND3_X2 U6633 ( .A1(n5231), .A2(n2337), .A3(n2504), .ZN(n5250) );
  MUX2_X2 U6634 ( .A(mem_16__11_), .B(mem_17__11_), .S(n3100), .Z(n5232) );
  INV_X4 U6635 ( .A(n5232), .ZN(n5235) );
  MUX2_X2 U6636 ( .A(mem_18__11_), .B(mem_19__11_), .S(n3100), .Z(n5233) );
  INV_X4 U6637 ( .A(n5233), .ZN(n5234) );
  MUX2_X2 U6638 ( .A(n5235), .B(n5234), .S(n3080), .Z(n5236) );
  NAND3_X2 U6639 ( .A1(n5236), .A2(n2331), .A3(n2364), .ZN(n5249) );
  MUX2_X2 U6640 ( .A(mem_20__11_), .B(mem_21__11_), .S(n3100), .Z(n5237) );
  INV_X4 U6641 ( .A(n5237), .ZN(n5240) );
  MUX2_X2 U6642 ( .A(mem_22__11_), .B(mem_23__11_), .S(n3100), .Z(n5238) );
  INV_X4 U6643 ( .A(n5238), .ZN(n5239) );
  MUX2_X2 U6644 ( .A(n5240), .B(n5239), .S(n3077), .Z(n5241) );
  NAND3_X2 U6645 ( .A1(n5241), .A2(n2346), .A3(n2366), .ZN(n5248) );
  MUX2_X2 U6646 ( .A(mem_8__11_), .B(mem_9__11_), .S(n3099), .Z(n5242) );
  INV_X4 U6647 ( .A(n5242), .ZN(n5245) );
  MUX2_X2 U6648 ( .A(mem_10__11_), .B(mem_11__11_), .S(n3099), .Z(n5243) );
  INV_X4 U6649 ( .A(n5243), .ZN(n5244) );
  MUX2_X2 U6650 ( .A(n5245), .B(n5244), .S(n3079), .Z(n5246) );
  NAND3_X2 U6651 ( .A1(n5246), .A2(n2343), .A3(n2367), .ZN(n5247) );
  NAND4_X2 U6652 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n5259)
         );
  MUX2_X2 U6653 ( .A(mem_0__11_), .B(mem_1__11_), .S(n3099), .Z(n5252) );
  MUX2_X2 U6654 ( .A(mem_2__11_), .B(mem_3__11_), .S(n3099), .Z(n5251) );
  MUX2_X2 U6655 ( .A(n5252), .B(n5251), .S(n3079), .Z(n5253) );
  NAND3_X2 U6656 ( .A1(n5253), .A2(n2328), .A3(n2368), .ZN(n5258) );
  MUX2_X2 U6657 ( .A(mem_4__11_), .B(mem_5__11_), .S(n3099), .Z(n5255) );
  MUX2_X2 U6658 ( .A(mem_6__11_), .B(mem_7__11_), .S(n3099), .Z(n5254) );
  MUX2_X2 U6659 ( .A(n5255), .B(n5254), .S(n3079), .Z(n5256) );
  NAND3_X2 U6660 ( .A1(n5256), .A2(n2341), .A3(n2369), .ZN(n5257) );
  OAI211_X2 U6661 ( .C1(n5260), .C2(n5259), .A(n5258), .B(n5257), .ZN(n7215)
         );
  MUX2_X2 U6662 ( .A(mem_28__12_), .B(mem_29__12_), .S(n3099), .Z(n5261) );
  INV_X4 U6663 ( .A(n5261), .ZN(n5264) );
  MUX2_X2 U6664 ( .A(mem_30__12_), .B(mem_31__12_), .S(n3099), .Z(n5262) );
  INV_X4 U6665 ( .A(n5262), .ZN(n5263) );
  MUX2_X2 U6666 ( .A(n5264), .B(n5263), .S(n3077), .Z(n5265) );
  NAND4_X2 U6667 ( .A1(n5265), .A2(n2332), .A3(n3060), .A4(n2374), .ZN(n5274)
         );
  MUX2_X2 U6668 ( .A(mem_24__12_), .B(mem_25__12_), .S(n3099), .Z(n5266) );
  INV_X4 U6669 ( .A(n5266), .ZN(n5269) );
  MUX2_X2 U6670 ( .A(mem_26__12_), .B(mem_27__12_), .S(n3099), .Z(n5267) );
  INV_X4 U6671 ( .A(n5267), .ZN(n5268) );
  MUX2_X2 U6672 ( .A(n5269), .B(n5268), .S(n3079), .Z(n5270) );
  NAND4_X2 U6673 ( .A1(n5270), .A2(n2344), .A3(n3060), .A4(n2503), .ZN(n5273)
         );
  NAND3_X2 U6674 ( .A1(n5274), .A2(n5273), .A3(n5272), .ZN(n5308) );
  MUX2_X2 U6675 ( .A(mem_12__12_), .B(mem_13__12_), .S(n3099), .Z(n5275) );
  INV_X4 U6676 ( .A(n5275), .ZN(n5278) );
  MUX2_X2 U6677 ( .A(mem_14__12_), .B(mem_15__12_), .S(n3099), .Z(n5276) );
  INV_X4 U6678 ( .A(n5276), .ZN(n5277) );
  MUX2_X2 U6679 ( .A(n5278), .B(n5277), .S(n3080), .Z(n5279) );
  NAND3_X2 U6680 ( .A1(n5279), .A2(n2338), .A3(n2504), .ZN(n5298) );
  MUX2_X2 U6681 ( .A(mem_16__12_), .B(mem_17__12_), .S(n3099), .Z(n5280) );
  INV_X4 U6682 ( .A(n5280), .ZN(n5283) );
  MUX2_X2 U6683 ( .A(mem_18__12_), .B(mem_19__12_), .S(n3099), .Z(n5281) );
  INV_X4 U6684 ( .A(n5281), .ZN(n5282) );
  MUX2_X2 U6685 ( .A(n5283), .B(n5282), .S(n3077), .Z(n5284) );
  NAND3_X2 U6686 ( .A1(n5284), .A2(n2332), .A3(n2364), .ZN(n5297) );
  MUX2_X2 U6687 ( .A(mem_20__12_), .B(mem_21__12_), .S(n3099), .Z(n5285) );
  INV_X4 U6688 ( .A(n5285), .ZN(n5288) );
  MUX2_X2 U6689 ( .A(mem_22__12_), .B(mem_23__12_), .S(n3099), .Z(n5286) );
  INV_X4 U6690 ( .A(n5286), .ZN(n5287) );
  MUX2_X2 U6691 ( .A(n5288), .B(n5287), .S(n3079), .Z(n5289) );
  NAND3_X2 U6692 ( .A1(n5289), .A2(n2330), .A3(n2366), .ZN(n5296) );
  MUX2_X2 U6693 ( .A(mem_8__12_), .B(mem_9__12_), .S(n3101), .Z(n5290) );
  INV_X4 U6694 ( .A(n5290), .ZN(n5293) );
  MUX2_X2 U6695 ( .A(mem_10__12_), .B(mem_11__12_), .S(n3092), .Z(n5291) );
  INV_X4 U6696 ( .A(n5291), .ZN(n5292) );
  MUX2_X2 U6697 ( .A(n5293), .B(n5292), .S(n3077), .Z(n5294) );
  NAND3_X2 U6698 ( .A1(n5294), .A2(n2327), .A3(n2367), .ZN(n5295) );
  NAND4_X2 U6699 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n5307)
         );
  MUX2_X2 U6700 ( .A(mem_0__12_), .B(mem_1__12_), .S(n3092), .Z(n5300) );
  MUX2_X2 U6701 ( .A(mem_2__12_), .B(mem_3__12_), .S(n3092), .Z(n5299) );
  MUX2_X2 U6702 ( .A(n5300), .B(n5299), .S(n3077), .Z(n5301) );
  NAND3_X2 U6703 ( .A1(n5301), .A2(n2335), .A3(n2368), .ZN(n5306) );
  MUX2_X2 U6704 ( .A(mem_4__12_), .B(mem_5__12_), .S(n3092), .Z(n5303) );
  MUX2_X2 U6705 ( .A(mem_6__12_), .B(mem_7__12_), .S(n3092), .Z(n5302) );
  MUX2_X2 U6706 ( .A(n5303), .B(n5302), .S(n3077), .Z(n5304) );
  NAND3_X2 U6707 ( .A1(n5304), .A2(n2331), .A3(n2369), .ZN(n5305) );
  OAI211_X2 U6708 ( .C1(n5308), .C2(n5307), .A(n5306), .B(n5305), .ZN(n7214)
         );
  MUX2_X2 U6709 ( .A(mem_28__13_), .B(mem_29__13_), .S(n3092), .Z(n5309) );
  INV_X4 U6710 ( .A(n5309), .ZN(n5312) );
  MUX2_X2 U6711 ( .A(mem_30__13_), .B(mem_31__13_), .S(n3092), .Z(n5310) );
  INV_X4 U6712 ( .A(n5310), .ZN(n5311) );
  MUX2_X2 U6713 ( .A(n5312), .B(n5311), .S(n3077), .Z(n5313) );
  NAND4_X2 U6714 ( .A1(n5313), .A2(n2329), .A3(n3060), .A4(n2374), .ZN(n5322)
         );
  MUX2_X2 U6715 ( .A(mem_24__13_), .B(mem_25__13_), .S(n3092), .Z(n5314) );
  INV_X4 U6716 ( .A(n5314), .ZN(n5317) );
  MUX2_X2 U6717 ( .A(mem_26__13_), .B(mem_27__13_), .S(n3092), .Z(n5315) );
  INV_X4 U6718 ( .A(n5315), .ZN(n5316) );
  MUX2_X2 U6719 ( .A(n5317), .B(n5316), .S(n3077), .Z(n5318) );
  NAND4_X2 U6720 ( .A1(n5318), .A2(n2341), .A3(n3060), .A4(n2503), .ZN(n5321)
         );
  NAND3_X2 U6721 ( .A1(n5322), .A2(n5321), .A3(n5320), .ZN(n5356) );
  MUX2_X2 U6722 ( .A(mem_12__13_), .B(mem_13__13_), .S(n3092), .Z(n5323) );
  INV_X4 U6723 ( .A(n5323), .ZN(n5326) );
  MUX2_X2 U6724 ( .A(mem_14__13_), .B(mem_15__13_), .S(n3092), .Z(n5324) );
  INV_X4 U6725 ( .A(n5324), .ZN(n5325) );
  MUX2_X2 U6726 ( .A(n5326), .B(n5325), .S(n3077), .Z(n5327) );
  NAND3_X2 U6727 ( .A1(n5327), .A2(n2328), .A3(n2504), .ZN(n5346) );
  MUX2_X2 U6728 ( .A(mem_16__13_), .B(mem_17__13_), .S(n3092), .Z(n5328) );
  INV_X4 U6729 ( .A(n5328), .ZN(n5331) );
  MUX2_X2 U6730 ( .A(mem_18__13_), .B(mem_19__13_), .S(n3092), .Z(n5329) );
  INV_X4 U6731 ( .A(n5329), .ZN(n5330) );
  MUX2_X2 U6732 ( .A(n5331), .B(n5330), .S(n3077), .Z(n5332) );
  NAND3_X2 U6733 ( .A1(n5332), .A2(n2343), .A3(n2364), .ZN(n5345) );
  MUX2_X2 U6734 ( .A(mem_20__13_), .B(mem_21__13_), .S(n3092), .Z(n5333) );
  INV_X4 U6735 ( .A(n5333), .ZN(n5336) );
  MUX2_X2 U6736 ( .A(mem_22__13_), .B(mem_23__13_), .S(n3091), .Z(n5334) );
  INV_X4 U6737 ( .A(n5334), .ZN(n5335) );
  MUX2_X2 U6738 ( .A(n5336), .B(n5335), .S(n3077), .Z(n5337) );
  NAND3_X2 U6739 ( .A1(n5337), .A2(n2345), .A3(n2366), .ZN(n5344) );
  MUX2_X2 U6740 ( .A(mem_8__13_), .B(mem_9__13_), .S(n3091), .Z(n5338) );
  INV_X4 U6741 ( .A(n5338), .ZN(n5341) );
  MUX2_X2 U6742 ( .A(mem_10__13_), .B(mem_11__13_), .S(n3091), .Z(n5339) );
  INV_X4 U6743 ( .A(n5339), .ZN(n5340) );
  MUX2_X2 U6744 ( .A(n5341), .B(n5340), .S(n3077), .Z(n5342) );
  NAND3_X2 U6745 ( .A1(n5342), .A2(n2328), .A3(n2367), .ZN(n5343) );
  NAND4_X2 U6746 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n5355)
         );
  MUX2_X2 U6747 ( .A(mem_0__13_), .B(mem_1__13_), .S(n3091), .Z(n5348) );
  MUX2_X2 U6748 ( .A(mem_2__13_), .B(mem_3__13_), .S(n3091), .Z(n5347) );
  MUX2_X2 U6749 ( .A(n5348), .B(n5347), .S(n3077), .Z(n5349) );
  NAND3_X2 U6750 ( .A1(n5349), .A2(n2335), .A3(n2368), .ZN(n5354) );
  MUX2_X2 U6751 ( .A(mem_4__13_), .B(mem_5__13_), .S(n3091), .Z(n5351) );
  MUX2_X2 U6752 ( .A(mem_6__13_), .B(mem_7__13_), .S(n3091), .Z(n5350) );
  MUX2_X2 U6753 ( .A(n5351), .B(n5350), .S(n3077), .Z(n5352) );
  NAND3_X2 U6754 ( .A1(n5352), .A2(n2329), .A3(n2369), .ZN(n5353) );
  OAI211_X2 U6755 ( .C1(n5356), .C2(n5355), .A(n5354), .B(n5353), .ZN(n7213)
         );
  MUX2_X2 U6756 ( .A(mem_28__14_), .B(mem_29__14_), .S(n3091), .Z(n5357) );
  INV_X4 U6757 ( .A(n5357), .ZN(n5360) );
  MUX2_X2 U6758 ( .A(mem_30__14_), .B(mem_31__14_), .S(n3091), .Z(n5358) );
  INV_X4 U6759 ( .A(n5358), .ZN(n5359) );
  MUX2_X2 U6760 ( .A(n5360), .B(n5359), .S(n3077), .Z(n5361) );
  NAND4_X2 U6761 ( .A1(n5361), .A2(n2335), .A3(n3060), .A4(n2374), .ZN(n5370)
         );
  MUX2_X2 U6762 ( .A(mem_24__14_), .B(mem_25__14_), .S(n3091), .Z(n5362) );
  INV_X4 U6763 ( .A(n5362), .ZN(n5365) );
  MUX2_X2 U6764 ( .A(mem_26__14_), .B(mem_27__14_), .S(n3091), .Z(n5363) );
  INV_X4 U6765 ( .A(n5363), .ZN(n5364) );
  MUX2_X2 U6766 ( .A(n5365), .B(n5364), .S(n3077), .Z(n5366) );
  NAND4_X2 U6767 ( .A1(n5366), .A2(n2340), .A3(n3060), .A4(n2503), .ZN(n5369)
         );
  NAND3_X2 U6768 ( .A1(n5370), .A2(n5369), .A3(n5368), .ZN(n5404) );
  MUX2_X2 U6769 ( .A(mem_12__14_), .B(mem_13__14_), .S(n3091), .Z(n5371) );
  INV_X4 U6770 ( .A(n5371), .ZN(n5374) );
  MUX2_X2 U6771 ( .A(mem_14__14_), .B(mem_15__14_), .S(n3091), .Z(n5372) );
  INV_X4 U6772 ( .A(n5372), .ZN(n5373) );
  MUX2_X2 U6773 ( .A(n5374), .B(n5373), .S(n3077), .Z(n5375) );
  NAND3_X2 U6774 ( .A1(n5375), .A2(n2340), .A3(n2504), .ZN(n5394) );
  MUX2_X2 U6775 ( .A(mem_16__14_), .B(mem_17__14_), .S(n3091), .Z(n5376) );
  INV_X4 U6776 ( .A(n5376), .ZN(n5379) );
  MUX2_X2 U6777 ( .A(mem_18__14_), .B(mem_19__14_), .S(n3091), .Z(n5377) );
  INV_X4 U6778 ( .A(n5377), .ZN(n5378) );
  MUX2_X2 U6779 ( .A(n5379), .B(n5378), .S(n3077), .Z(n5380) );
  NAND3_X2 U6780 ( .A1(n5380), .A2(n2332), .A3(n2364), .ZN(n5393) );
  MUX2_X2 U6781 ( .A(mem_20__14_), .B(mem_21__14_), .S(n3091), .Z(n5381) );
  INV_X4 U6782 ( .A(n5381), .ZN(n5384) );
  MUX2_X2 U6783 ( .A(mem_22__14_), .B(mem_23__14_), .S(n3091), .Z(n5382) );
  INV_X4 U6784 ( .A(n5382), .ZN(n5383) );
  MUX2_X2 U6785 ( .A(n5384), .B(n5383), .S(n3076), .Z(n5385) );
  NAND3_X2 U6786 ( .A1(n5385), .A2(n2330), .A3(n2366), .ZN(n5392) );
  MUX2_X2 U6787 ( .A(mem_8__14_), .B(mem_9__14_), .S(n3091), .Z(n5386) );
  INV_X4 U6788 ( .A(n5386), .ZN(n5389) );
  MUX2_X2 U6789 ( .A(mem_10__14_), .B(mem_11__14_), .S(n3091), .Z(n5387) );
  INV_X4 U6790 ( .A(n5387), .ZN(n5388) );
  MUX2_X2 U6791 ( .A(n5389), .B(n5388), .S(n3076), .Z(n5390) );
  NAND3_X2 U6792 ( .A1(n5390), .A2(n2335), .A3(n2367), .ZN(n5391) );
  NAND4_X2 U6793 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n5403)
         );
  MUX2_X2 U6794 ( .A(mem_0__14_), .B(mem_1__14_), .S(n3091), .Z(n5396) );
  MUX2_X2 U6795 ( .A(mem_2__14_), .B(mem_3__14_), .S(n3091), .Z(n5395) );
  MUX2_X2 U6796 ( .A(n5396), .B(n5395), .S(n3076), .Z(n5397) );
  NAND3_X2 U6797 ( .A1(n5397), .A2(n2330), .A3(n2368), .ZN(n5402) );
  MUX2_X2 U6798 ( .A(mem_4__14_), .B(mem_5__14_), .S(n3090), .Z(n5399) );
  MUX2_X2 U6799 ( .A(mem_6__14_), .B(mem_7__14_), .S(n3090), .Z(n5398) );
  MUX2_X2 U6800 ( .A(n5399), .B(n5398), .S(n3076), .Z(n5400) );
  NAND3_X2 U6801 ( .A1(n5400), .A2(n2328), .A3(n2369), .ZN(n5401) );
  OAI211_X2 U6802 ( .C1(n5404), .C2(n5403), .A(n5402), .B(n5401), .ZN(n7212)
         );
  MUX2_X2 U6803 ( .A(mem_28__15_), .B(mem_29__15_), .S(n3090), .Z(n5405) );
  INV_X4 U6804 ( .A(n5405), .ZN(n5408) );
  MUX2_X2 U6805 ( .A(mem_30__15_), .B(mem_31__15_), .S(n3090), .Z(n5406) );
  INV_X4 U6806 ( .A(n5406), .ZN(n5407) );
  MUX2_X2 U6807 ( .A(n5408), .B(n5407), .S(n3076), .Z(n5409) );
  NAND4_X2 U6808 ( .A1(n5409), .A2(n2332), .A3(n3060), .A4(n2374), .ZN(n5418)
         );
  MUX2_X2 U6809 ( .A(mem_24__15_), .B(mem_25__15_), .S(n3090), .Z(n5410) );
  INV_X4 U6810 ( .A(n5410), .ZN(n5413) );
  MUX2_X2 U6811 ( .A(mem_26__15_), .B(mem_27__15_), .S(n3090), .Z(n5411) );
  INV_X4 U6812 ( .A(n5411), .ZN(n5412) );
  MUX2_X2 U6813 ( .A(n5413), .B(n5412), .S(n3076), .Z(n5414) );
  NAND4_X2 U6814 ( .A1(n5414), .A2(n2343), .A3(n3060), .A4(n2503), .ZN(n5417)
         );
  NAND3_X2 U6815 ( .A1(n5418), .A2(n5417), .A3(n5416), .ZN(n5452) );
  MUX2_X2 U6816 ( .A(mem_12__15_), .B(mem_13__15_), .S(n3090), .Z(n5419) );
  INV_X4 U6817 ( .A(n5419), .ZN(n5422) );
  MUX2_X2 U6818 ( .A(mem_14__15_), .B(mem_15__15_), .S(n3090), .Z(n5420) );
  INV_X4 U6819 ( .A(n5420), .ZN(n5421) );
  MUX2_X2 U6820 ( .A(n5422), .B(n5421), .S(n3076), .Z(n5423) );
  NAND3_X2 U6821 ( .A1(n5423), .A2(n2337), .A3(n2504), .ZN(n5442) );
  MUX2_X2 U6822 ( .A(mem_16__15_), .B(mem_17__15_), .S(n3090), .Z(n5424) );
  INV_X4 U6823 ( .A(n5424), .ZN(n5427) );
  MUX2_X2 U6824 ( .A(mem_18__15_), .B(mem_19__15_), .S(n3090), .Z(n5425) );
  INV_X4 U6825 ( .A(n5425), .ZN(n5426) );
  MUX2_X2 U6826 ( .A(n5427), .B(n5426), .S(n3076), .Z(n5428) );
  NAND3_X2 U6827 ( .A1(n5428), .A2(n2344), .A3(n2364), .ZN(n5441) );
  MUX2_X2 U6828 ( .A(mem_20__15_), .B(mem_21__15_), .S(n3090), .Z(n5429) );
  INV_X4 U6829 ( .A(n5429), .ZN(n5432) );
  MUX2_X2 U6830 ( .A(mem_22__15_), .B(mem_23__15_), .S(n3090), .Z(n5430) );
  INV_X4 U6831 ( .A(n5430), .ZN(n5431) );
  MUX2_X2 U6832 ( .A(n5432), .B(n5431), .S(n3076), .Z(n5433) );
  NAND3_X2 U6833 ( .A1(n5433), .A2(n2339), .A3(n2366), .ZN(n5440) );
  MUX2_X2 U6834 ( .A(mem_8__15_), .B(mem_9__15_), .S(n3090), .Z(n5434) );
  INV_X4 U6835 ( .A(n5434), .ZN(n5437) );
  MUX2_X2 U6836 ( .A(mem_10__15_), .B(mem_11__15_), .S(n3090), .Z(n5435) );
  INV_X4 U6837 ( .A(n5435), .ZN(n5436) );
  MUX2_X2 U6838 ( .A(n5437), .B(n5436), .S(n3076), .Z(n5438) );
  NAND3_X2 U6839 ( .A1(n5438), .A2(n2331), .A3(n2367), .ZN(n5439) );
  NAND4_X2 U6840 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n5451)
         );
  MUX2_X2 U6841 ( .A(mem_0__15_), .B(mem_1__15_), .S(n3090), .Z(n5444) );
  MUX2_X2 U6842 ( .A(mem_2__15_), .B(mem_3__15_), .S(n3090), .Z(n5443) );
  MUX2_X2 U6843 ( .A(n5444), .B(n5443), .S(n3076), .Z(n5445) );
  NAND3_X2 U6844 ( .A1(n5445), .A2(n2345), .A3(n2368), .ZN(n5450) );
  MUX2_X2 U6845 ( .A(mem_4__15_), .B(mem_5__15_), .S(n3090), .Z(n5447) );
  MUX2_X2 U6846 ( .A(mem_6__15_), .B(mem_7__15_), .S(n3090), .Z(n5446) );
  MUX2_X2 U6847 ( .A(n5447), .B(n5446), .S(n3076), .Z(n5448) );
  NAND3_X2 U6848 ( .A1(n5448), .A2(n2331), .A3(n2369), .ZN(n5449) );
  OAI211_X2 U6849 ( .C1(n5452), .C2(n5451), .A(n5450), .B(n5449), .ZN(n7211)
         );
  MUX2_X2 U6850 ( .A(mem_28__16_), .B(mem_29__16_), .S(n3090), .Z(n5453) );
  INV_X4 U6851 ( .A(n5453), .ZN(n5456) );
  MUX2_X2 U6852 ( .A(mem_30__16_), .B(mem_31__16_), .S(n3090), .Z(n5454) );
  INV_X4 U6853 ( .A(n5454), .ZN(n5455) );
  MUX2_X2 U6854 ( .A(n5456), .B(n5455), .S(n3076), .Z(n5457) );
  NAND4_X2 U6855 ( .A1(n5457), .A2(n2331), .A3(n3060), .A4(n2374), .ZN(n5466)
         );
  MUX2_X2 U6856 ( .A(mem_24__16_), .B(mem_25__16_), .S(n3089), .Z(n5458) );
  INV_X4 U6857 ( .A(n5458), .ZN(n5461) );
  MUX2_X2 U6858 ( .A(mem_26__16_), .B(mem_27__16_), .S(n3089), .Z(n5459) );
  INV_X4 U6859 ( .A(n5459), .ZN(n5460) );
  MUX2_X2 U6860 ( .A(n5461), .B(n5460), .S(n3076), .Z(n5462) );
  NAND4_X2 U6861 ( .A1(n5462), .A2(n2337), .A3(n3060), .A4(n2503), .ZN(n5465)
         );
  NAND3_X2 U6862 ( .A1(n5466), .A2(n5465), .A3(n5464), .ZN(n5500) );
  MUX2_X2 U6863 ( .A(mem_12__16_), .B(mem_13__16_), .S(n3089), .Z(n5467) );
  INV_X4 U6864 ( .A(n5467), .ZN(n5470) );
  MUX2_X2 U6865 ( .A(mem_14__16_), .B(mem_15__16_), .S(n3089), .Z(n5468) );
  INV_X4 U6866 ( .A(n5468), .ZN(n5469) );
  MUX2_X2 U6867 ( .A(n5470), .B(n5469), .S(n3076), .Z(n5471) );
  NAND3_X2 U6868 ( .A1(n5471), .A2(n2329), .A3(n2504), .ZN(n5490) );
  MUX2_X2 U6869 ( .A(mem_16__16_), .B(mem_17__16_), .S(n3089), .Z(n5472) );
  INV_X4 U6870 ( .A(n5472), .ZN(n5475) );
  MUX2_X2 U6871 ( .A(mem_18__16_), .B(mem_19__16_), .S(n3089), .Z(n5473) );
  INV_X4 U6872 ( .A(n5473), .ZN(n5474) );
  MUX2_X2 U6873 ( .A(n5475), .B(n5474), .S(n3075), .Z(n5476) );
  NAND3_X2 U6874 ( .A1(n5476), .A2(n2336), .A3(n2364), .ZN(n5489) );
  MUX2_X2 U6875 ( .A(mem_20__16_), .B(mem_21__16_), .S(n3089), .Z(n5477) );
  INV_X4 U6876 ( .A(n5477), .ZN(n5480) );
  MUX2_X2 U6877 ( .A(mem_22__16_), .B(mem_23__16_), .S(n3089), .Z(n5478) );
  INV_X4 U6878 ( .A(n5478), .ZN(n5479) );
  MUX2_X2 U6879 ( .A(n5480), .B(n5479), .S(n3075), .Z(n5481) );
  NAND3_X2 U6880 ( .A1(n5481), .A2(n2340), .A3(n2366), .ZN(n5488) );
  MUX2_X2 U6881 ( .A(mem_8__16_), .B(mem_9__16_), .S(n3089), .Z(n5482) );
  INV_X4 U6882 ( .A(n5482), .ZN(n5485) );
  MUX2_X2 U6883 ( .A(mem_10__16_), .B(mem_11__16_), .S(n3089), .Z(n5483) );
  INV_X4 U6884 ( .A(n5483), .ZN(n5484) );
  MUX2_X2 U6885 ( .A(n5485), .B(n5484), .S(n3076), .Z(n5486) );
  NAND3_X2 U6886 ( .A1(n5486), .A2(n2327), .A3(n2367), .ZN(n5487) );
  NAND4_X2 U6887 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n5499)
         );
  MUX2_X2 U6888 ( .A(mem_0__16_), .B(mem_1__16_), .S(n3089), .Z(n5492) );
  MUX2_X2 U6889 ( .A(mem_2__16_), .B(mem_3__16_), .S(n3089), .Z(n5491) );
  MUX2_X2 U6890 ( .A(n5492), .B(n5491), .S(n3075), .Z(n5493) );
  NAND3_X2 U6891 ( .A1(n5493), .A2(n2340), .A3(n2368), .ZN(n5498) );
  MUX2_X2 U6892 ( .A(mem_4__16_), .B(mem_5__16_), .S(n3089), .Z(n5495) );
  MUX2_X2 U6893 ( .A(mem_6__16_), .B(mem_7__16_), .S(n3089), .Z(n5494) );
  MUX2_X2 U6894 ( .A(n5495), .B(n5494), .S(n3077), .Z(n5496) );
  NAND3_X2 U6895 ( .A1(n5496), .A2(n2330), .A3(n2369), .ZN(n5497) );
  OAI211_X2 U6896 ( .C1(n5500), .C2(n5499), .A(n5498), .B(n5497), .ZN(n7210)
         );
  MUX2_X2 U6897 ( .A(mem_28__17_), .B(mem_29__17_), .S(n3089), .Z(n5501) );
  INV_X4 U6898 ( .A(n5501), .ZN(n5504) );
  MUX2_X2 U6899 ( .A(mem_30__17_), .B(mem_31__17_), .S(n3089), .Z(n5502) );
  INV_X4 U6900 ( .A(n5502), .ZN(n5503) );
  MUX2_X2 U6901 ( .A(n5504), .B(n5503), .S(n3075), .Z(n5505) );
  NAND4_X2 U6902 ( .A1(n5505), .A2(n2344), .A3(n3060), .A4(n2374), .ZN(n5514)
         );
  MUX2_X2 U6903 ( .A(mem_24__17_), .B(mem_25__17_), .S(n3089), .Z(n5506) );
  INV_X4 U6904 ( .A(n5506), .ZN(n5509) );
  MUX2_X2 U6905 ( .A(mem_26__17_), .B(mem_27__17_), .S(n3089), .Z(n5507) );
  INV_X4 U6906 ( .A(n5507), .ZN(n5508) );
  MUX2_X2 U6907 ( .A(n5509), .B(n5508), .S(n3075), .Z(n5510) );
  NAND4_X2 U6908 ( .A1(n5510), .A2(n2336), .A3(n3060), .A4(n2503), .ZN(n5513)
         );
  NAND3_X2 U6909 ( .A1(n5514), .A2(n5513), .A3(n5512), .ZN(n5548) );
  MUX2_X2 U6910 ( .A(mem_12__17_), .B(mem_13__17_), .S(n3089), .Z(n5515) );
  INV_X4 U6911 ( .A(n5515), .ZN(n5518) );
  MUX2_X2 U6912 ( .A(mem_14__17_), .B(mem_15__17_), .S(n3089), .Z(n5516) );
  INV_X4 U6913 ( .A(n5516), .ZN(n5517) );
  MUX2_X2 U6914 ( .A(n5518), .B(n5517), .S(n3075), .Z(n5519) );
  NAND3_X2 U6915 ( .A1(n5519), .A2(n2328), .A3(n2504), .ZN(n5538) );
  MUX2_X2 U6916 ( .A(mem_16__17_), .B(mem_17__17_), .S(n3089), .Z(n5520) );
  INV_X4 U6917 ( .A(n5520), .ZN(n5523) );
  MUX2_X2 U6918 ( .A(mem_18__17_), .B(mem_19__17_), .S(n3088), .Z(n5521) );
  INV_X4 U6919 ( .A(n5521), .ZN(n5522) );
  MUX2_X2 U6920 ( .A(n5523), .B(n5522), .S(n3075), .Z(n5524) );
  NAND3_X2 U6921 ( .A1(n5524), .A2(n2339), .A3(n2364), .ZN(n5537) );
  MUX2_X2 U6922 ( .A(mem_20__17_), .B(mem_21__17_), .S(n3088), .Z(n5525) );
  INV_X4 U6923 ( .A(n5525), .ZN(n5528) );
  MUX2_X2 U6924 ( .A(mem_22__17_), .B(mem_23__17_), .S(n3090), .Z(n5526) );
  INV_X4 U6925 ( .A(n5526), .ZN(n5527) );
  MUX2_X2 U6926 ( .A(n5528), .B(n5527), .S(n3075), .Z(n5529) );
  NAND3_X2 U6927 ( .A1(n5529), .A2(n2329), .A3(n2366), .ZN(n5536) );
  MUX2_X2 U6928 ( .A(mem_8__17_), .B(mem_9__17_), .S(n3092), .Z(n5530) );
  INV_X4 U6929 ( .A(n5530), .ZN(n5533) );
  MUX2_X2 U6930 ( .A(mem_10__17_), .B(mem_11__17_), .S(n3092), .Z(n5531) );
  INV_X4 U6931 ( .A(n5531), .ZN(n5532) );
  MUX2_X2 U6932 ( .A(n5533), .B(n5532), .S(n3075), .Z(n5534) );
  NAND3_X2 U6933 ( .A1(n5534), .A2(n2344), .A3(n2367), .ZN(n5535) );
  NAND4_X2 U6934 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n5547)
         );
  MUX2_X2 U6935 ( .A(mem_0__17_), .B(mem_1__17_), .S(n3092), .Z(n5540) );
  MUX2_X2 U6936 ( .A(mem_2__17_), .B(mem_3__17_), .S(n3092), .Z(n5539) );
  MUX2_X2 U6937 ( .A(n5540), .B(n5539), .S(n3075), .Z(n5541) );
  NAND3_X2 U6938 ( .A1(n5541), .A2(n2339), .A3(n2368), .ZN(n5546) );
  MUX2_X2 U6939 ( .A(mem_4__17_), .B(mem_5__17_), .S(n3092), .Z(n5543) );
  MUX2_X2 U6940 ( .A(mem_6__17_), .B(mem_7__17_), .S(n3092), .Z(n5542) );
  MUX2_X2 U6941 ( .A(n5543), .B(n5542), .S(n3075), .Z(n5544) );
  NAND3_X2 U6942 ( .A1(n5544), .A2(n2329), .A3(n2369), .ZN(n5545) );
  OAI211_X2 U6943 ( .C1(n5548), .C2(n5547), .A(n5546), .B(n5545), .ZN(n7209)
         );
  MUX2_X2 U6944 ( .A(mem_28__18_), .B(mem_29__18_), .S(n3092), .Z(n5549) );
  INV_X4 U6945 ( .A(n5549), .ZN(n5552) );
  MUX2_X2 U6946 ( .A(mem_30__18_), .B(mem_31__18_), .S(n3093), .Z(n5550) );
  INV_X4 U6947 ( .A(n5550), .ZN(n5551) );
  MUX2_X2 U6948 ( .A(n5552), .B(n5551), .S(n3075), .Z(n5553) );
  NAND4_X2 U6949 ( .A1(n5553), .A2(n2337), .A3(n3060), .A4(n2374), .ZN(n5562)
         );
  MUX2_X2 U6950 ( .A(mem_24__18_), .B(mem_25__18_), .S(n3093), .Z(n5554) );
  INV_X4 U6951 ( .A(n5554), .ZN(n5557) );
  MUX2_X2 U6952 ( .A(mem_26__18_), .B(mem_27__18_), .S(n3093), .Z(n5555) );
  INV_X4 U6953 ( .A(n5555), .ZN(n5556) );
  MUX2_X2 U6954 ( .A(n5557), .B(n5556), .S(n3075), .Z(n5558) );
  NAND4_X2 U6955 ( .A1(n5558), .A2(n2340), .A3(n3060), .A4(n2503), .ZN(n5561)
         );
  NAND3_X2 U6956 ( .A1(n5562), .A2(n5561), .A3(n5560), .ZN(n5596) );
  MUX2_X2 U6957 ( .A(mem_12__18_), .B(mem_13__18_), .S(n3093), .Z(n5563) );
  INV_X4 U6958 ( .A(n5563), .ZN(n5566) );
  MUX2_X2 U6959 ( .A(mem_14__18_), .B(mem_15__18_), .S(n3093), .Z(n5564) );
  INV_X4 U6960 ( .A(n5564), .ZN(n5565) );
  MUX2_X2 U6961 ( .A(n5566), .B(n5565), .S(n3075), .Z(n5567) );
  NAND3_X2 U6962 ( .A1(n5567), .A2(n2327), .A3(n2504), .ZN(n5586) );
  MUX2_X2 U6963 ( .A(mem_16__18_), .B(mem_17__18_), .S(n3093), .Z(n5568) );
  INV_X4 U6964 ( .A(n5568), .ZN(n5571) );
  MUX2_X2 U6965 ( .A(mem_18__18_), .B(mem_19__18_), .S(n3093), .Z(n5569) );
  INV_X4 U6966 ( .A(n5569), .ZN(n5570) );
  MUX2_X2 U6967 ( .A(n5571), .B(n5570), .S(n3075), .Z(n5572) );
  NAND3_X2 U6968 ( .A1(n5572), .A2(n2338), .A3(n2364), .ZN(n5585) );
  MUX2_X2 U6969 ( .A(mem_20__18_), .B(mem_21__18_), .S(n3093), .Z(n5573) );
  INV_X4 U6970 ( .A(n5573), .ZN(n5576) );
  MUX2_X2 U6971 ( .A(mem_22__18_), .B(mem_23__18_), .S(n3093), .Z(n5574) );
  INV_X4 U6972 ( .A(n5574), .ZN(n5575) );
  MUX2_X2 U6973 ( .A(n5576), .B(n5575), .S(n3074), .Z(n5577) );
  NAND3_X2 U6974 ( .A1(n5577), .A2(n2330), .A3(n2366), .ZN(n5584) );
  MUX2_X2 U6975 ( .A(mem_8__18_), .B(mem_9__18_), .S(n3093), .Z(n5578) );
  INV_X4 U6976 ( .A(n5578), .ZN(n5581) );
  MUX2_X2 U6977 ( .A(mem_10__18_), .B(mem_11__18_), .S(n3093), .Z(n5579) );
  INV_X4 U6978 ( .A(n5579), .ZN(n5580) );
  MUX2_X2 U6979 ( .A(n5581), .B(n5580), .S(n3075), .Z(n5582) );
  NAND3_X2 U6980 ( .A1(n5582), .A2(n2346), .A3(n2367), .ZN(n5583) );
  NAND4_X2 U6981 ( .A1(n5586), .A2(n5585), .A3(n5584), .A4(n5583), .ZN(n5595)
         );
  MUX2_X2 U6982 ( .A(mem_0__18_), .B(mem_1__18_), .S(n3093), .Z(n5588) );
  MUX2_X2 U6983 ( .A(mem_2__18_), .B(mem_3__18_), .S(n3093), .Z(n5587) );
  MUX2_X2 U6984 ( .A(n5588), .B(n5587), .S(n3074), .Z(n5589) );
  NAND3_X2 U6985 ( .A1(n5589), .A2(n2334), .A3(n2368), .ZN(n5594) );
  MUX2_X2 U6986 ( .A(mem_4__18_), .B(mem_5__18_), .S(n3093), .Z(n5591) );
  MUX2_X2 U6987 ( .A(mem_6__18_), .B(mem_7__18_), .S(n3093), .Z(n5590) );
  MUX2_X2 U6988 ( .A(n5591), .B(n5590), .S(n3074), .Z(n5592) );
  NAND3_X2 U6989 ( .A1(n5592), .A2(n2344), .A3(n2369), .ZN(n5593) );
  OAI211_X2 U6990 ( .C1(n5596), .C2(n5595), .A(n5594), .B(n5593), .ZN(n7208)
         );
  MUX2_X2 U6991 ( .A(mem_28__19_), .B(mem_29__19_), .S(n3093), .Z(n5597) );
  INV_X4 U6992 ( .A(n5597), .ZN(n5600) );
  MUX2_X2 U6993 ( .A(mem_30__19_), .B(mem_31__19_), .S(n3101), .Z(n5598) );
  INV_X4 U6994 ( .A(n5598), .ZN(n5599) );
  MUX2_X2 U6995 ( .A(n5600), .B(n5599), .S(n3074), .Z(n5601) );
  NAND4_X2 U6996 ( .A1(n5601), .A2(n2333), .A3(n3059), .A4(n2374), .ZN(n5610)
         );
  MUX2_X2 U6997 ( .A(mem_24__19_), .B(mem_25__19_), .S(n3093), .Z(n5602) );
  INV_X4 U6998 ( .A(n5602), .ZN(n5605) );
  MUX2_X2 U6999 ( .A(mem_26__19_), .B(mem_27__19_), .S(n3093), .Z(n5603) );
  INV_X4 U7000 ( .A(n5603), .ZN(n5604) );
  MUX2_X2 U7001 ( .A(n5605), .B(n5604), .S(n3074), .Z(n5606) );
  NAND4_X2 U7002 ( .A1(n5606), .A2(n2342), .A3(n3059), .A4(n2503), .ZN(n5609)
         );
  NAND3_X2 U7003 ( .A1(n5610), .A2(n5609), .A3(n5608), .ZN(n5644) );
  MUX2_X2 U7004 ( .A(mem_12__19_), .B(mem_13__19_), .S(n3093), .Z(n5611) );
  INV_X4 U7005 ( .A(n5611), .ZN(n5614) );
  MUX2_X2 U7006 ( .A(mem_14__19_), .B(mem_15__19_), .S(n3093), .Z(n5612) );
  INV_X4 U7007 ( .A(n5612), .ZN(n5613) );
  MUX2_X2 U7008 ( .A(n5614), .B(n5613), .S(n3074), .Z(n5615) );
  NAND3_X2 U7009 ( .A1(n5615), .A2(n2337), .A3(n2504), .ZN(n5634) );
  MUX2_X2 U7010 ( .A(mem_16__19_), .B(mem_17__19_), .S(n3093), .Z(n5616) );
  INV_X4 U7011 ( .A(n5616), .ZN(n5619) );
  MUX2_X2 U7012 ( .A(mem_18__19_), .B(mem_19__19_), .S(n3094), .Z(n5617) );
  INV_X4 U7013 ( .A(n5617), .ZN(n5618) );
  MUX2_X2 U7014 ( .A(n5619), .B(n5618), .S(n3074), .Z(n5620) );
  NAND3_X2 U7015 ( .A1(n5620), .A2(n2328), .A3(n2364), .ZN(n5633) );
  MUX2_X2 U7016 ( .A(mem_20__19_), .B(mem_21__19_), .S(n3094), .Z(n5621) );
  INV_X4 U7017 ( .A(n5621), .ZN(n5624) );
  MUX2_X2 U7018 ( .A(mem_22__19_), .B(mem_23__19_), .S(n3094), .Z(n5622) );
  INV_X4 U7019 ( .A(n5622), .ZN(n5623) );
  MUX2_X2 U7020 ( .A(n5624), .B(n5623), .S(n3074), .Z(n5625) );
  NAND3_X2 U7021 ( .A1(n5625), .A2(n2344), .A3(n2366), .ZN(n5632) );
  MUX2_X2 U7022 ( .A(mem_8__19_), .B(mem_9__19_), .S(n3094), .Z(n5626) );
  INV_X4 U7023 ( .A(n5626), .ZN(n5629) );
  MUX2_X2 U7024 ( .A(mem_10__19_), .B(mem_11__19_), .S(n3094), .Z(n5627) );
  INV_X4 U7025 ( .A(n5627), .ZN(n5628) );
  MUX2_X2 U7026 ( .A(n5629), .B(n5628), .S(n3074), .Z(n5630) );
  NAND3_X2 U7027 ( .A1(n5630), .A2(n2345), .A3(n2367), .ZN(n5631) );
  NAND4_X2 U7028 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n5643)
         );
  MUX2_X2 U7029 ( .A(mem_0__19_), .B(mem_1__19_), .S(n3094), .Z(n5636) );
  MUX2_X2 U7030 ( .A(mem_2__19_), .B(mem_3__19_), .S(n3094), .Z(n5635) );
  MUX2_X2 U7031 ( .A(n5636), .B(n5635), .S(n3074), .Z(n5637) );
  NAND3_X2 U7032 ( .A1(n5637), .A2(n2333), .A3(n2368), .ZN(n5642) );
  MUX2_X2 U7033 ( .A(mem_4__19_), .B(mem_5__19_), .S(n3094), .Z(n5639) );
  MUX2_X2 U7034 ( .A(mem_6__19_), .B(mem_7__19_), .S(n3094), .Z(n5638) );
  MUX2_X2 U7035 ( .A(n5639), .B(n5638), .S(n3074), .Z(n5640) );
  NAND3_X2 U7036 ( .A1(n5640), .A2(n2343), .A3(n2369), .ZN(n5641) );
  OAI211_X2 U7037 ( .C1(n5644), .C2(n5643), .A(n5642), .B(n5641), .ZN(n7207)
         );
  MUX2_X2 U7038 ( .A(mem_28__20_), .B(mem_29__20_), .S(n3094), .Z(n5645) );
  INV_X4 U7039 ( .A(n5645), .ZN(n5648) );
  MUX2_X2 U7040 ( .A(mem_30__20_), .B(mem_31__20_), .S(n3094), .Z(n5646) );
  INV_X4 U7041 ( .A(n5646), .ZN(n5647) );
  MUX2_X2 U7042 ( .A(n5648), .B(n5647), .S(n3074), .Z(n5649) );
  NAND4_X2 U7043 ( .A1(n5649), .A2(n2333), .A3(n3059), .A4(n2374), .ZN(n5658)
         );
  MUX2_X2 U7044 ( .A(mem_24__20_), .B(mem_25__20_), .S(n3094), .Z(n5650) );
  INV_X4 U7045 ( .A(n5650), .ZN(n5653) );
  MUX2_X2 U7046 ( .A(mem_26__20_), .B(mem_27__20_), .S(n3094), .Z(n5651) );
  INV_X4 U7047 ( .A(n5651), .ZN(n5652) );
  MUX2_X2 U7048 ( .A(n5653), .B(n5652), .S(n3074), .Z(n5654) );
  NAND4_X2 U7049 ( .A1(n5654), .A2(n2344), .A3(n3060), .A4(n2503), .ZN(n5657)
         );
  NAND3_X2 U7050 ( .A1(n5658), .A2(n5657), .A3(n5656), .ZN(n5692) );
  MUX2_X2 U7051 ( .A(mem_12__20_), .B(mem_13__20_), .S(n3094), .Z(n5659) );
  INV_X4 U7052 ( .A(n5659), .ZN(n5662) );
  MUX2_X2 U7053 ( .A(mem_14__20_), .B(mem_15__20_), .S(n3094), .Z(n5660) );
  INV_X4 U7054 ( .A(n5660), .ZN(n5661) );
  MUX2_X2 U7055 ( .A(n5662), .B(n5661), .S(n3074), .Z(n5663) );
  NAND3_X2 U7056 ( .A1(n5663), .A2(n2333), .A3(n2504), .ZN(n5682) );
  MUX2_X2 U7057 ( .A(mem_16__20_), .B(mem_17__20_), .S(n3094), .Z(n5664) );
  INV_X4 U7058 ( .A(n5664), .ZN(n5667) );
  MUX2_X2 U7059 ( .A(mem_18__20_), .B(mem_19__20_), .S(n3094), .Z(n5665) );
  INV_X4 U7060 ( .A(n5665), .ZN(n5666) );
  MUX2_X2 U7061 ( .A(n5667), .B(n5666), .S(n3074), .Z(n5668) );
  NAND3_X2 U7062 ( .A1(n5668), .A2(n2329), .A3(n2364), .ZN(n5681) );
  MUX2_X2 U7063 ( .A(mem_20__20_), .B(mem_21__20_), .S(n3094), .Z(n5669) );
  INV_X4 U7064 ( .A(n5669), .ZN(n5672) );
  MUX2_X2 U7065 ( .A(mem_22__20_), .B(mem_23__20_), .S(n3094), .Z(n5670) );
  INV_X4 U7066 ( .A(n5670), .ZN(n5671) );
  MUX2_X2 U7067 ( .A(n5672), .B(n5671), .S(n3074), .Z(n5673) );
  NAND3_X2 U7068 ( .A1(n5673), .A2(n2332), .A3(n2366), .ZN(n5680) );
  MUX2_X2 U7069 ( .A(mem_8__20_), .B(mem_9__20_), .S(n3094), .Z(n5674) );
  INV_X4 U7070 ( .A(n5674), .ZN(n5677) );
  MUX2_X2 U7071 ( .A(mem_10__20_), .B(mem_11__20_), .S(n3094), .Z(n5675) );
  INV_X4 U7072 ( .A(n5675), .ZN(n5676) );
  MUX2_X2 U7073 ( .A(n5677), .B(n5676), .S(n3077), .Z(n5678) );
  NAND3_X2 U7074 ( .A1(n5678), .A2(n2339), .A3(n2367), .ZN(n5679) );
  NAND4_X2 U7075 ( .A1(n5682), .A2(n5681), .A3(n5680), .A4(n5679), .ZN(n5691)
         );
  MUX2_X2 U7076 ( .A(mem_0__20_), .B(mem_1__20_), .S(n3101), .Z(n5684) );
  MUX2_X2 U7077 ( .A(mem_2__20_), .B(mem_3__20_), .S(n3101), .Z(n5683) );
  MUX2_X2 U7078 ( .A(n5684), .B(n5683), .S(n3077), .Z(n5685) );
  NAND3_X2 U7079 ( .A1(n5685), .A2(n2339), .A3(n2368), .ZN(n5690) );
  MUX2_X2 U7080 ( .A(mem_4__20_), .B(mem_5__20_), .S(n3101), .Z(n5687) );
  MUX2_X2 U7081 ( .A(mem_6__20_), .B(mem_7__20_), .S(n3101), .Z(n5686) );
  MUX2_X2 U7082 ( .A(n5687), .B(n5686), .S(n3079), .Z(n5688) );
  NAND3_X2 U7083 ( .A1(n5688), .A2(n2332), .A3(n2369), .ZN(n5689) );
  OAI211_X2 U7084 ( .C1(n5692), .C2(n5691), .A(n5690), .B(n5689), .ZN(n7206)
         );
  MUX2_X2 U7085 ( .A(mem_28__21_), .B(mem_29__21_), .S(n3101), .Z(n5693) );
  INV_X4 U7086 ( .A(n5693), .ZN(n5696) );
  MUX2_X2 U7087 ( .A(mem_30__21_), .B(mem_31__21_), .S(n3101), .Z(n5694) );
  INV_X4 U7088 ( .A(n5694), .ZN(n5695) );
  MUX2_X2 U7089 ( .A(n5696), .B(n5695), .S(n3079), .Z(n5697) );
  NAND4_X2 U7090 ( .A1(n5697), .A2(n2328), .A3(n3059), .A4(n2374), .ZN(n5707)
         );
  MUX2_X2 U7091 ( .A(mem_24__21_), .B(mem_25__21_), .S(n3101), .Z(n5698) );
  INV_X4 U7092 ( .A(n5698), .ZN(n5701) );
  MUX2_X2 U7093 ( .A(mem_26__21_), .B(mem_27__21_), .S(n3101), .Z(n5699) );
  INV_X4 U7094 ( .A(n5699), .ZN(n5700) );
  MUX2_X2 U7095 ( .A(n5701), .B(n5700), .S(n3077), .Z(n5702) );
  NAND4_X2 U7096 ( .A1(n5702), .A2(n2346), .A3(n3059), .A4(n2503), .ZN(n5706)
         );
  NAND3_X2 U7097 ( .A1(n5707), .A2(n5706), .A3(n5705), .ZN(n5742) );
  MUX2_X2 U7098 ( .A(mem_12__21_), .B(mem_13__21_), .S(n3101), .Z(n5708) );
  INV_X4 U7099 ( .A(n5708), .ZN(n5711) );
  MUX2_X2 U7100 ( .A(mem_14__21_), .B(mem_15__21_), .S(n3101), .Z(n5709) );
  INV_X4 U7101 ( .A(n5709), .ZN(n5710) );
  MUX2_X2 U7102 ( .A(n5711), .B(n5710), .S(n3080), .Z(n5712) );
  NAND3_X2 U7103 ( .A1(n5712), .A2(n2334), .A3(n2504), .ZN(n5731) );
  MUX2_X2 U7104 ( .A(mem_16__21_), .B(mem_17__21_), .S(n3101), .Z(n5713) );
  INV_X4 U7105 ( .A(n5713), .ZN(n5716) );
  MUX2_X2 U7106 ( .A(mem_18__21_), .B(mem_19__21_), .S(n3101), .Z(n5714) );
  INV_X4 U7107 ( .A(n5714), .ZN(n5715) );
  MUX2_X2 U7108 ( .A(n5716), .B(n5715), .S(n3079), .Z(n5717) );
  NAND3_X2 U7109 ( .A1(n5717), .A2(n2330), .A3(n2364), .ZN(n5730) );
  MUX2_X2 U7110 ( .A(mem_20__21_), .B(mem_21__21_), .S(n3101), .Z(n5718) );
  INV_X4 U7111 ( .A(n5718), .ZN(n5721) );
  MUX2_X2 U7112 ( .A(mem_22__21_), .B(mem_23__21_), .S(n3101), .Z(n5719) );
  INV_X4 U7113 ( .A(n5719), .ZN(n5720) );
  MUX2_X2 U7114 ( .A(n5721), .B(n5720), .S(n3078), .Z(n5722) );
  NAND3_X2 U7115 ( .A1(n5722), .A2(n2331), .A3(n2366), .ZN(n5729) );
  MUX2_X2 U7116 ( .A(mem_8__21_), .B(mem_9__21_), .S(n3101), .Z(n5723) );
  INV_X4 U7117 ( .A(n5723), .ZN(n5726) );
  MUX2_X2 U7118 ( .A(mem_10__21_), .B(mem_11__21_), .S(n3101), .Z(n5724) );
  INV_X4 U7119 ( .A(n5724), .ZN(n5725) );
  MUX2_X2 U7120 ( .A(n5726), .B(n5725), .S(n3080), .Z(n5727) );
  NAND3_X2 U7121 ( .A1(n5727), .A2(n2342), .A3(n2367), .ZN(n5728) );
  NAND4_X2 U7122 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n5741)
         );
  MUX2_X2 U7123 ( .A(mem_0__21_), .B(mem_1__21_), .S(n3101), .Z(n5733) );
  MUX2_X2 U7124 ( .A(mem_2__21_), .B(mem_3__21_), .S(n3101), .Z(n5732) );
  MUX2_X2 U7125 ( .A(n5733), .B(n5732), .S(n3080), .Z(n5734) );
  NAND3_X2 U7126 ( .A1(n5734), .A2(n2327), .A3(n2368), .ZN(n5740) );
  MUX2_X2 U7127 ( .A(mem_4__21_), .B(mem_5__21_), .S(n3101), .Z(n5736) );
  MUX2_X2 U7128 ( .A(mem_6__21_), .B(mem_7__21_), .S(n3101), .Z(n5735) );
  MUX2_X2 U7129 ( .A(n5736), .B(n5735), .S(n3080), .Z(n5738) );
  NAND3_X2 U7130 ( .A1(n5738), .A2(n2342), .A3(n2369), .ZN(n5739) );
  OAI211_X2 U7131 ( .C1(n5742), .C2(n5741), .A(n5740), .B(n5739), .ZN(n7205)
         );
  MUX2_X2 U7132 ( .A(mem_12__22_), .B(mem_13__22_), .S(n3101), .Z(n5744) );
  NAND2_X2 U7133 ( .A1(n5745), .A2(n3062), .ZN(n5754) );
  MUX2_X2 U7134 ( .A(mem_18__22_), .B(mem_19__22_), .S(n3101), .Z(n5747) );
  NAND2_X2 U7135 ( .A1(n5748), .A2(n3064), .ZN(n5753) );
  MUX2_X2 U7136 ( .A(mem_14__22_), .B(mem_15__22_), .S(n3101), .Z(n5750) );
  NAND2_X2 U7137 ( .A1(n5751), .A2(n3062), .ZN(n5752) );
  NAND3_X2 U7138 ( .A1(n5754), .A2(n5753), .A3(n5752), .ZN(n5793) );
  MUX2_X2 U7139 ( .A(mem_30__22_), .B(mem_31__22_), .S(n3102), .Z(n5755) );
  NAND3_X2 U7140 ( .A1(n3063), .A2(n5755), .A3(n5798), .ZN(n5760) );
  MUX2_X2 U7141 ( .A(mem_28__22_), .B(mem_29__22_), .S(n3098), .Z(n5757) );
  NAND3_X2 U7142 ( .A1(n3063), .A2(n5757), .A3(n5756), .ZN(n5759) );
  NAND3_X2 U7143 ( .A1(n5760), .A2(n5759), .A3(n5758), .ZN(n5779) );
  MUX2_X2 U7144 ( .A(mem_22__22_), .B(mem_23__22_), .S(n3099), .Z(n5761) );
  NAND3_X2 U7145 ( .A1(n3059), .A2(n5761), .A3(n2382), .ZN(n5770) );
  MUX2_X2 U7146 ( .A(mem_24__22_), .B(mem_25__22_), .S(n3098), .Z(n5762) );
  NAND3_X2 U7147 ( .A1(n3063), .A2(n5762), .A3(n2861), .ZN(n5769) );
  MUX2_X2 U7148 ( .A(mem_26__22_), .B(mem_27__22_), .S(n3098), .Z(n5764) );
  NAND3_X2 U7149 ( .A1(n3063), .A2(n5764), .A3(n5763), .ZN(n5768) );
  MUX2_X2 U7150 ( .A(mem_20__22_), .B(mem_21__22_), .S(n3098), .Z(n5766) );
  NAND3_X2 U7151 ( .A1(n3061), .A2(n5766), .A3(n5765), .ZN(n5767) );
  NAND4_X2 U7152 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n5778)
         );
  OAI221_X2 U7153 ( .B1(mem_11__22_), .B2(n3105), .C1(n3103), .C2(mem_10__22_), 
        .A(n3081), .ZN(n5773) );
  NAND4_X2 U7154 ( .A1(n2367), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n5777)
         );
  MUX2_X2 U7155 ( .A(mem_16__22_), .B(mem_17__22_), .S(n3101), .Z(n5774) );
  NAND2_X2 U7156 ( .A1(n5775), .A2(n3064), .ZN(n5776) );
  OAI211_X2 U7157 ( .C1(n5779), .C2(n5778), .A(n5777), .B(n5776), .ZN(n5792)
         );
  OAI211_X2 U7158 ( .C1(n5783), .C2(n5782), .A(n5781), .B(n5780), .ZN(n5789)
         );
  OAI211_X2 U7159 ( .C1(n5787), .C2(n5786), .A(n5785), .B(n5784), .ZN(n5788)
         );
  MUX2_X2 U7160 ( .A(n5789), .B(n5788), .S(n3067), .Z(n5790) );
  NAND3_X2 U7161 ( .A1(n5790), .A2(n3064), .A3(n3062), .ZN(n5791) );
  MUX2_X2 U7162 ( .A(n5794), .B(wData[22]), .S(n2347), .Z(n7204) );
  NAND2_X2 U7163 ( .A1(n5798), .A2(n3104), .ZN(n6145) );
  AOI211_X4 U7164 ( .C1(n5803), .C2(n5802), .A(n2383), .B(n2543), .ZN(n5813)
         );
  NOR3_X4 U7165 ( .A1(n5809), .A2(n5808), .A3(n5807), .ZN(n5810) );
  MUX2_X2 U7166 ( .A(n5813), .B(n5812), .S(n3063), .Z(n5833) );
  NOR2_X4 U7167 ( .A1(mem_29__23_), .A2(n2869), .ZN(n5826) );
  MUX2_X2 U7168 ( .A(n5831), .B(n5830), .S(n3063), .Z(n5832) );
  MUX2_X2 U7169 ( .A(n5833), .B(n5832), .S(n3059), .Z(n5834) );
  INV_X4 U7170 ( .A(n5834), .ZN(n5835) );
  MUX2_X2 U7171 ( .A(n5835), .B(wData[23]), .S(n2347), .Z(n7203) );
  NOR3_X4 U7172 ( .A1(n5841), .A2(n5840), .A3(n5839), .ZN(n5842) );
  AOI211_X4 U7173 ( .C1(n5843), .C2(n5842), .A(n2386), .B(n2544), .ZN(n5853)
         );
  NOR3_X4 U7174 ( .A1(n5849), .A2(n5848), .A3(n5847), .ZN(n5850) );
  MUX2_X2 U7175 ( .A(n5853), .B(n5852), .S(n3063), .Z(n5873) );
  NOR3_X4 U7176 ( .A1(n5859), .A2(n5858), .A3(n5857), .ZN(n5860) );
  NOR3_X4 U7177 ( .A1(n5867), .A2(n5866), .A3(n5865), .ZN(n5868) );
  MUX2_X2 U7178 ( .A(n5873), .B(n5872), .S(n3059), .Z(n5874) );
  INV_X4 U7179 ( .A(n5874), .ZN(n5875) );
  MUX2_X2 U7180 ( .A(n5875), .B(wData[24]), .S(n2347), .Z(n7202) );
  NOR3_X4 U7181 ( .A1(n5889), .A2(n5888), .A3(n5887), .ZN(n5890) );
  MUX2_X2 U7182 ( .A(n5893), .B(n5892), .S(n3063), .Z(n5913) );
  NOR3_X4 U7183 ( .A1(n5899), .A2(n5898), .A3(n5897), .ZN(n5900) );
  NOR3_X4 U7184 ( .A1(n5907), .A2(n5906), .A3(n5905), .ZN(n5908) );
  MUX2_X2 U7185 ( .A(n5911), .B(n5910), .S(n3063), .Z(n5912) );
  MUX2_X2 U7186 ( .A(n5913), .B(n5912), .S(n3059), .Z(n5914) );
  INV_X4 U7187 ( .A(n5914), .ZN(n5915) );
  MUX2_X2 U7188 ( .A(n5915), .B(wData[25]), .S(n2347), .Z(n7201) );
  MUX2_X2 U7189 ( .A(n5933), .B(n5932), .S(n3063), .Z(n5953) );
  NOR3_X4 U7190 ( .A1(n5939), .A2(n5938), .A3(n5937), .ZN(n5940) );
  NOR3_X4 U7191 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n5948) );
  MUX2_X2 U7192 ( .A(n5953), .B(n5952), .S(n3059), .Z(n5954) );
  INV_X4 U7193 ( .A(n5954), .ZN(n5955) );
  MUX2_X2 U7194 ( .A(n5955), .B(wData[26]), .S(n2347), .Z(n7200) );
  NOR3_X4 U7195 ( .A1(n5961), .A2(n5960), .A3(n5959), .ZN(n5962) );
  AOI211_X4 U7196 ( .C1(n5963), .C2(n5962), .A(n2398), .B(n2547), .ZN(n5973)
         );
  NOR3_X4 U7197 ( .A1(n5969), .A2(n5968), .A3(n5967), .ZN(n5970) );
  MUX2_X2 U7198 ( .A(n5973), .B(n5972), .S(n3063), .Z(n5993) );
  NOR3_X4 U7199 ( .A1(n5979), .A2(n5978), .A3(n5977), .ZN(n5980) );
  NOR3_X4 U7200 ( .A1(n5987), .A2(n5986), .A3(n5985), .ZN(n5988) );
  MUX2_X2 U7201 ( .A(n5991), .B(n5990), .S(n3063), .Z(n5992) );
  MUX2_X2 U7202 ( .A(n5993), .B(n5992), .S(n3059), .Z(n5994) );
  INV_X4 U7203 ( .A(n5994), .ZN(n5995) );
  MUX2_X2 U7204 ( .A(n5995), .B(wData[27]), .S(n2347), .Z(n7199) );
  MUX2_X2 U7205 ( .A(n6013), .B(n6012), .S(n3063), .Z(n6033) );
  NOR3_X4 U7206 ( .A1(n6019), .A2(n6018), .A3(n6017), .ZN(n6020) );
  NOR3_X4 U7207 ( .A1(n6027), .A2(n6026), .A3(n6025), .ZN(n6028) );
  MUX2_X2 U7208 ( .A(n6031), .B(n6030), .S(n3063), .Z(n6032) );
  MUX2_X2 U7209 ( .A(n6033), .B(n6032), .S(n3059), .Z(n6034) );
  INV_X4 U7210 ( .A(n6034), .ZN(n6035) );
  MUX2_X2 U7211 ( .A(n6035), .B(wData[28]), .S(n2347), .Z(n7198) );
  NOR3_X4 U7212 ( .A1(n6049), .A2(n6048), .A3(n6047), .ZN(n6050) );
  MUX2_X2 U7213 ( .A(n6053), .B(n6052), .S(n3063), .Z(n6073) );
  NOR3_X4 U7214 ( .A1(n6067), .A2(n6066), .A3(n6065), .ZN(n6068) );
  MUX2_X2 U7215 ( .A(n6071), .B(n6070), .S(n3063), .Z(n6072) );
  MUX2_X2 U7216 ( .A(n6073), .B(n6072), .S(n3059), .Z(n6074) );
  INV_X4 U7217 ( .A(n6074), .ZN(n6075) );
  MUX2_X2 U7218 ( .A(n6075), .B(wData[29]), .S(n2347), .Z(n7197) );
  NOR3_X4 U7219 ( .A1(n6089), .A2(n6088), .A3(n6087), .ZN(n6090) );
  MUX2_X2 U7220 ( .A(n6093), .B(n6092), .S(n3063), .Z(n6113) );
  NOR3_X4 U7221 ( .A1(n6107), .A2(n6106), .A3(n6105), .ZN(n6108) );
  MUX2_X2 U7222 ( .A(n6111), .B(n6110), .S(n3063), .Z(n6112) );
  MUX2_X2 U7223 ( .A(n6113), .B(n6112), .S(n3059), .Z(n6114) );
  INV_X4 U7224 ( .A(n6114), .ZN(n6115) );
  MUX2_X2 U7225 ( .A(n6115), .B(wData[30]), .S(n2347), .Z(n7196) );
  NOR3_X4 U7226 ( .A1(n6129), .A2(n6128), .A3(n6127), .ZN(n6130) );
  MUX2_X2 U7227 ( .A(n6133), .B(n6132), .S(n3063), .Z(n6155) );
  NOR3_X4 U7228 ( .A1(n6139), .A2(n6138), .A3(n6137), .ZN(n6140) );
  NOR2_X4 U7229 ( .A1(mem_29__31_), .A2(n2871), .ZN(n6148) );
  NOR3_X4 U7230 ( .A1(n6149), .A2(n6148), .A3(n6147), .ZN(n6150) );
  MUX2_X2 U7231 ( .A(n6153), .B(n6152), .S(n3063), .Z(n6154) );
  MUX2_X2 U7232 ( .A(n6155), .B(n6154), .S(n3059), .Z(n6156) );
  INV_X4 U7233 ( .A(n6156), .ZN(n6157) );
  MUX2_X2 U7234 ( .A(n6157), .B(wData[31]), .S(n2347), .Z(n7195) );
  NOR2_X1 U7235 ( .A1(n3164), .A2(rd[0]), .ZN(n6158) );
  OAI22_X1 U7236 ( .A1(n6158), .A2(n6165), .B1(rs2[1]), .B2(n6158), .ZN(n6162)
         );
  AND2_X1 U7237 ( .A1(rd[0]), .A2(n3164), .ZN(n6159) );
  OAI22_X1 U7238 ( .A1(rd[1]), .A2(n6159), .B1(n6159), .B2(n3155), .ZN(n6161)
         );
  XNOR2_X1 U7239 ( .A(n3134), .B(rd[2]), .ZN(n6160) );
  XOR2_X1 U7240 ( .A(n3114), .B(rd[3]), .Z(n6164) );
  XOR2_X1 U7241 ( .A(rs2[4]), .B(rd[4]), .Z(n6163) );
  INV_X4 U7242 ( .A(rd[1]), .ZN(n6165) );
  NOR2_X1 U7243 ( .A1(n3110), .A2(rd[0]), .ZN(n6166) );
  OAI22_X1 U7244 ( .A1(n6166), .A2(n6165), .B1(n3082), .B2(n6166), .ZN(n6170)
         );
  AND2_X1 U7245 ( .A1(rd[0]), .A2(n3107), .ZN(n6167) );
  OAI22_X1 U7246 ( .A1(rd[1]), .A2(n6167), .B1(n6167), .B2(n3085), .ZN(n6169)
         );
  XNOR2_X1 U7247 ( .A(n3067), .B(rd[2]), .ZN(n6168) );
  NAND3_X1 U7248 ( .A1(n6170), .A2(n6169), .A3(n6168), .ZN(n6171) );
  INV_X4 U7249 ( .A(rd[4]), .ZN(n7227) );
  INV_X4 U7250 ( .A(rd[3]), .ZN(n7228) );
  INV_X4 U7251 ( .A(rd[2]), .ZN(n7229) );
  INV_X4 U7252 ( .A(rd[0]), .ZN(n7230) );
  SDFF_X1 rData2_reg_23_ ( .D(n4170), .SI(wData[23]), .SE(n2350), .CK(n2238), 
        .Q(rData2[23]) );
  SDFF_X1 rData2_reg_26_ ( .D(n4359), .SI(wData[26]), .SE(n2349), .CK(n2238), 
        .Q(rData2[26]) );
endmodule

