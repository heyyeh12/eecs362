
module alu ( a, b, alu_ctrl, inverse_set, res, zf, of, cf );
  input [31:0] a;
  input [31:0] b;
  input [3:0] alu_ctrl;
  output [31:0] res;
  input inverse_set;
  output zf, of, cf;
  wire   n76, n90, n91, n92, n93, n97, n98, n100, n109, n111, n112, n115, n246,
         n248, n558, n559, n560, n564, n570, n573, n577, n580, n582, n585,
         n586, n587, n588, n589, n592, n593, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1882, n1883;

  NOR4_X2 U421 ( .A1(n592), .A2(b[23]), .A3(b[25]), .A4(b[24]), .ZN(n589) );
  NOR4_X2 U423 ( .A1(n593), .A2(b[16]), .A3(b[18]), .A4(b[17]), .ZN(n588) );
  NAND4_X2 U424 ( .A1(n100), .A2(n1288), .A3(n98), .A4(n97), .ZN(n593) );
  INV_X4 U598 ( .A(a[5]), .ZN(n76) );
  INV_X4 U631 ( .A(b[8]), .ZN(n109) );
  INV_X4 U633 ( .A(b[6]), .ZN(n111) );
  INV_X4 U634 ( .A(b[5]), .ZN(n112) );
  INV_X4 U637 ( .A(b[4]), .ZN(n115) );
  AOI22_X1 U660 ( .A1(n1716), .A2(n1640), .B1(n1720), .B2(n1778), .ZN(n1173)
         );
  INV_X8 U661 ( .A(n1727), .ZN(n1721) );
  NAND4_X2 U662 ( .A1(n1581), .A2(n1574), .A3(n1577), .A4(n1573), .ZN(n630) );
  NAND4_X2 U663 ( .A1(n1581), .A2(n1574), .A3(n1577), .A4(n1573), .ZN(n1522)
         );
  AND2_X2 U664 ( .A1(n630), .A2(n1388), .ZN(n655) );
  XOR2_X1 U665 ( .A(n1757), .B(n685), .Z(n642) );
  XNOR2_X2 U666 ( .A(n1426), .B(n671), .ZN(n1750) );
  NAND2_X2 U667 ( .A1(n1375), .A2(n1396), .ZN(n1426) );
  OAI221_X4 U668 ( .B1(n1486), .B2(n1452), .C1(n1494), .C2(n1449), .A(n776), 
        .ZN(n1317) );
  INV_X4 U669 ( .A(n683), .ZN(n631) );
  INV_X4 U670 ( .A(n683), .ZN(n632) );
  INV_X8 U671 ( .A(n1882), .ZN(n682) );
  NOR2_X4 U672 ( .A1(n838), .A2(n1840), .ZN(n1882) );
  INV_X8 U673 ( .A(n682), .ZN(n683) );
  OAI21_X2 U674 ( .B1(n1281), .B2(n1309), .A(n1194), .ZN(n1079) );
  OAI21_X2 U675 ( .B1(n1221), .B2(n1309), .A(n1194), .ZN(n1154) );
  NAND2_X2 U676 ( .A1(b[1]), .A2(n1883), .ZN(n246) );
  INV_X4 U677 ( .A(n1406), .ZN(n1432) );
  NOR3_X2 U678 ( .A1(n1760), .A2(n1759), .A3(n1758), .ZN(n1761) );
  NOR2_X2 U679 ( .A1(n775), .A2(n774), .ZN(n1453) );
  NAND2_X2 U680 ( .A1(n1499), .A2(n1454), .ZN(n1449) );
  NAND2_X2 U681 ( .A1(a[2]), .A2(n801), .ZN(n1693) );
  NOR2_X2 U682 ( .A1(alu_ctrl[2]), .A2(alu_ctrl[0]), .ZN(n945) );
  INV_X4 U683 ( .A(n653), .ZN(n671) );
  OAI21_X2 U684 ( .B1(n1210), .B2(n1309), .A(n1194), .ZN(n1195) );
  OAI21_X2 U685 ( .B1(n1269), .B2(n1309), .A(n1194), .ZN(n1105) );
  NOR3_X2 U686 ( .A1(n1123), .A2(n1066), .A3(n1124), .ZN(n1067) );
  OAI21_X2 U687 ( .B1(n1211), .B2(n687), .A(n1140), .ZN(n1117) );
  INV_X4 U688 ( .A(n694), .ZN(n692) );
  NOR2_X2 U689 ( .A1(n1682), .A2(n637), .ZN(n1686) );
  NAND3_X2 U690 ( .A1(n1094), .A2(n1093), .A3(n1092), .ZN(n1657) );
  AOI21_X2 U691 ( .B1(n1223), .B2(n1427), .A(n1091), .ZN(n1092) );
  AOI222_X1 U692 ( .A1(n1722), .A2(n1587), .B1(n1844), .B2(n1559), .C1(n1719), 
        .C2(n1558), .ZN(n1560) );
  NOR2_X2 U693 ( .A1(n633), .A2(n1783), .ZN(n1548) );
  AOI222_X1 U694 ( .A1(n1587), .A2(n1844), .B1(n1722), .B2(n1559), .C1(n1659), 
        .C2(n1558), .ZN(n1275) );
  NAND4_X2 U695 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(n592) );
  NOR2_X2 U696 ( .A1(b[5]), .A2(b[6]), .ZN(n701) );
  INV_X4 U697 ( .A(b[10]), .ZN(n674) );
  NAND2_X2 U698 ( .A1(n759), .A2(n760), .ZN(n757) );
  NOR3_X2 U699 ( .A1(n1318), .A2(n1334), .A3(n780), .ZN(n823) );
  NAND3_X2 U700 ( .A1(n1459), .A2(n1454), .A3(n1499), .ZN(n780) );
  NAND3_X2 U701 ( .A1(n1335), .A2(n1376), .A3(n652), .ZN(n745) );
  AOI21_X2 U702 ( .B1(b[3]), .B2(n984), .A(n1882), .ZN(n871) );
  INV_X8 U703 ( .A(n560), .ZN(n688) );
  NOR2_X2 U704 ( .A1(n586), .A2(alu_ctrl[1]), .ZN(n560) );
  AOI21_X2 U705 ( .B1(n651), .B2(n1824), .A(n1823), .ZN(n1825) );
  INV_X4 U706 ( .A(n683), .ZN(n924) );
  AOI21_X2 U707 ( .B1(n1482), .B2(n1454), .A(n1453), .ZN(n1455) );
  AOI21_X2 U708 ( .B1(n1025), .B2(n1029), .A(n651), .ZN(n830) );
  NOR2_X2 U709 ( .A1(n641), .A2(n921), .ZN(n859) );
  NAND3_X2 U710 ( .A1(n1851), .A2(n1850), .A3(n1849), .ZN(n1856) );
  NOR3_X2 U711 ( .A1(res[22]), .A2(res[23]), .A3(res[24]), .ZN(n1865) );
  NOR2_X2 U712 ( .A1(res[25]), .A2(res[26]), .ZN(n1866) );
  NOR3_X2 U713 ( .A1(res[15]), .A2(res[16]), .A3(res[17]), .ZN(n1861) );
  NOR2_X2 U714 ( .A1(res[20]), .A2(res[21]), .ZN(n1862) );
  NOR2_X2 U715 ( .A1(n1840), .A2(n649), .ZN(n1842) );
  AOI21_X2 U716 ( .B1(n1671), .B2(n1670), .A(n1669), .ZN(n1674) );
  NOR2_X2 U717 ( .A1(n1667), .A2(n1695), .ZN(n1671) );
  NOR2_X2 U718 ( .A1(a[8]), .A2(n696), .ZN(n1601) );
  OAI21_X2 U719 ( .B1(a[12]), .B2(n697), .A(n693), .ZN(n1515) );
  NOR2_X2 U720 ( .A1(a[13]), .A2(n696), .ZN(n1502) );
  AOI21_X2 U721 ( .B1(n1484), .B2(n1483), .A(n1482), .ZN(n1485) );
  NOR2_X2 U722 ( .A1(n1357), .A2(n1356), .ZN(n1506) );
  NOR2_X2 U723 ( .A1(n248), .A2(n1407), .ZN(n1265) );
  NOR2_X2 U724 ( .A1(n1403), .A2(n1365), .ZN(n1264) );
  NAND3_X2 U725 ( .A1(n1274), .A2(n1273), .A3(n1272), .ZN(n1559) );
  NOR2_X2 U726 ( .A1(a[23]), .A2(n696), .ZN(n1204) );
  NAND2_X2 U727 ( .A1(n1189), .A2(n1169), .ZN(n1172) );
  NAND2_X2 U728 ( .A1(n1131), .A2(n1071), .ZN(n1073) );
  AOI222_X2 U729 ( .A1(n982), .A2(n981), .B1(n1102), .B2(n690), .C1(n1053), 
        .C2(n1427), .ZN(n1714) );
  OAI21_X2 U730 ( .B1(n1222), .B2(n687), .A(n1140), .ZN(n1141) );
  INV_X4 U731 ( .A(n694), .ZN(n693) );
  NOR2_X2 U732 ( .A1(n651), .A2(n935), .ZN(n942) );
  NOR2_X2 U733 ( .A1(res[30]), .A2(n1878), .ZN(n1875) );
  NOR2_X2 U734 ( .A1(n1728), .A2(n649), .ZN(n1729) );
  OAI21_X2 U735 ( .B1(n1738), .B2(n1737), .A(n1736), .ZN(n1743) );
  NOR2_X2 U736 ( .A1(n691), .A2(n1733), .ZN(n1738) );
  OAI21_X2 U737 ( .B1(n691), .B2(n1735), .A(b[1]), .ZN(n1736) );
  NOR2_X2 U738 ( .A1(n656), .A2(n633), .ZN(n1742) );
  OAI21_X2 U739 ( .B1(a[2]), .B2(n696), .A(n693), .ZN(n1712) );
  NOR2_X2 U740 ( .A1(n1699), .A2(n1698), .ZN(n1700) );
  OAI21_X2 U741 ( .B1(a[3]), .B2(n696), .A(n692), .ZN(n1697) );
  NOR2_X2 U742 ( .A1(n654), .A2(n633), .ZN(n1701) );
  NOR2_X2 U743 ( .A1(n1706), .A2(n1705), .ZN(n1707) );
  NOR2_X2 U744 ( .A1(n1704), .A2(n637), .ZN(n1705) );
  NOR2_X2 U745 ( .A1(n1714), .A2(n636), .ZN(n1706) );
  NOR2_X2 U746 ( .A1(n1676), .A2(n115), .ZN(n1677) );
  OAI21_X2 U747 ( .B1(a[4]), .B2(n696), .A(n692), .ZN(n1675) );
  NOR2_X2 U748 ( .A1(n1755), .A2(n633), .ZN(n1678) );
  AOI21_X2 U749 ( .B1(n1652), .B2(n1651), .A(n112), .ZN(n1655) );
  AOI21_X2 U750 ( .B1(n76), .B2(n698), .A(n691), .ZN(n1652) );
  NOR2_X2 U751 ( .A1(n1653), .A2(n76), .ZN(n1654) );
  AOI21_X2 U752 ( .B1(n112), .B2(n698), .A(n691), .ZN(n1653) );
  NOR2_X2 U753 ( .A1(n633), .A2(n1762), .ZN(n1656) );
  NOR2_X2 U754 ( .A1(n1635), .A2(n111), .ZN(n1636) );
  OAI21_X2 U755 ( .B1(a[6]), .B2(n697), .A(n692), .ZN(n1634) );
  AOI21_X2 U756 ( .B1(n1633), .B2(n692), .A(n1632), .ZN(n1637) );
  NOR2_X2 U757 ( .A1(n1617), .A2(n1616), .ZN(n1618) );
  OAI21_X2 U758 ( .B1(a[7]), .B2(n697), .A(n692), .ZN(n1615) );
  NOR2_X2 U759 ( .A1(n1614), .A2(n634), .ZN(n1619) );
  NOR2_X2 U760 ( .A1(n1579), .A2(n1578), .ZN(n1580) );
  OAI21_X2 U761 ( .B1(n1568), .B2(n1567), .A(n1566), .ZN(n1571) );
  NOR2_X2 U762 ( .A1(n691), .A2(n1564), .ZN(n1568) );
  OAI21_X2 U763 ( .B1(n691), .B2(n1565), .A(b[9]), .ZN(n1566) );
  NOR2_X2 U764 ( .A1(n1569), .A2(n634), .ZN(n1570) );
  NOR2_X2 U765 ( .A1(n1609), .A2(n649), .ZN(n1585) );
  OAI21_X2 U766 ( .B1(a[10]), .B2(n697), .A(n693), .ZN(n1553) );
  OAI21_X2 U767 ( .B1(a[11]), .B2(n696), .A(n693), .ZN(n1534) );
  NOR2_X2 U768 ( .A1(n1506), .A2(n649), .ZN(n1478) );
  NOR2_X2 U769 ( .A1(n1476), .A2(n1475), .ZN(n1477) );
  OAI21_X2 U770 ( .B1(a[14]), .B2(n697), .A(n692), .ZN(n1474) );
  NOR2_X2 U771 ( .A1(n1409), .A2(n1408), .ZN(n1413) );
  NOR2_X2 U772 ( .A1(n1407), .A2(n1406), .ZN(n1408) );
  NOR2_X2 U773 ( .A1(n1424), .A2(n637), .ZN(n1425) );
  NOR2_X2 U774 ( .A1(n1506), .A2(n637), .ZN(n1420) );
  OAI21_X2 U775 ( .B1(n1419), .B2(n1418), .A(n1417), .ZN(n1421) );
  OAI21_X2 U776 ( .B1(n694), .B2(n1416), .A(b[17]), .ZN(n1417) );
  NOR2_X2 U777 ( .A1(n694), .A2(n1415), .ZN(n1419) );
  OAI221_X2 U778 ( .B1(n248), .B2(n1404), .C1(n1403), .C2(n1406), .A(n1402), 
        .ZN(n1488) );
  NOR2_X2 U779 ( .A1(n1506), .A2(n636), .ZN(n1362) );
  NOR2_X2 U780 ( .A1(n1360), .A2(n1359), .ZN(n1361) );
  OAI21_X2 U781 ( .B1(a[18]), .B2(n697), .A(n692), .ZN(n1358) );
  NOR2_X2 U782 ( .A1(n1368), .A2(n1367), .ZN(n1369) );
  NOR2_X2 U783 ( .A1(n1366), .A2(n1365), .ZN(n1367) );
  NOR2_X2 U784 ( .A1(n248), .A2(n1364), .ZN(n1368) );
  NOR2_X2 U785 ( .A1(n1514), .A2(n636), .ZN(n1345) );
  OAI21_X2 U786 ( .B1(n1341), .B2(n1340), .A(n1339), .ZN(n1346) );
  OAI21_X2 U787 ( .B1(n694), .B2(n1338), .A(b[19]), .ZN(n1339) );
  NOR2_X2 U788 ( .A1(n694), .A2(n1337), .ZN(n1341) );
  NOR2_X2 U789 ( .A1(a[19]), .A2(n696), .ZN(n1338) );
  NOR2_X2 U790 ( .A1(n1327), .A2(n633), .ZN(n1348) );
  NOR2_X2 U791 ( .A1(n1330), .A2(n1329), .ZN(n1331) );
  NOR2_X2 U792 ( .A1(n1312), .A2(n1311), .ZN(n1313) );
  NOR2_X2 U793 ( .A1(n1407), .A2(n1365), .ZN(n1311) );
  NOR2_X2 U794 ( .A1(n248), .A2(n1405), .ZN(n1312) );
  NOR2_X2 U795 ( .A1(n1315), .A2(n637), .ZN(n1316) );
  NOR2_X2 U796 ( .A1(n1315), .A2(n636), .ZN(n1291) );
  NOR2_X2 U797 ( .A1(n1289), .A2(n1288), .ZN(n1290) );
  OAI21_X2 U798 ( .B1(a[20]), .B2(n697), .A(n692), .ZN(n1287) );
  NOR2_X2 U799 ( .A1(n1298), .A2(n1297), .ZN(n1299) );
  NOR2_X2 U800 ( .A1(n1371), .A2(n1365), .ZN(n1297) );
  NOR2_X2 U801 ( .A1(n248), .A2(n1366), .ZN(n1298) );
  NOR2_X2 U802 ( .A1(n1302), .A2(n1301), .ZN(n1303) );
  NOR2_X2 U803 ( .A1(n1545), .A2(n637), .ZN(n1301) );
  NOR2_X2 U804 ( .A1(n1555), .A2(n634), .ZN(n1302) );
  NOR2_X2 U805 ( .A1(n1555), .A2(n649), .ZN(n1267) );
  OAI21_X2 U806 ( .B1(a[21]), .B2(n697), .A(n692), .ZN(n1252) );
  NOR2_X2 U807 ( .A1(n1569), .A2(n636), .ZN(n1230) );
  NOR2_X2 U808 ( .A1(n1228), .A2(n97), .ZN(n1229) );
  OAI21_X2 U809 ( .B1(a[22]), .B2(n697), .A(n692), .ZN(n1227) );
  NOR2_X2 U810 ( .A1(n1242), .A2(n1241), .ZN(n1246) );
  NOR2_X2 U811 ( .A1(n1244), .A2(n1243), .ZN(n1245) );
  NOR2_X2 U812 ( .A1(n1370), .A2(n1365), .ZN(n1241) );
  NOR2_X2 U813 ( .A1(n1197), .A2(n1196), .ZN(n1202) );
  NOR2_X2 U814 ( .A1(n1200), .A2(n1199), .ZN(n1201) );
  NOR2_X2 U815 ( .A1(n1314), .A2(n1365), .ZN(n1196) );
  NOR2_X2 U816 ( .A1(n1148), .A2(n1147), .ZN(n1149) );
  OAI21_X2 U817 ( .B1(a[24]), .B2(n696), .A(n692), .ZN(n1146) );
  NOR2_X2 U818 ( .A1(n1614), .A2(n636), .ZN(n1150) );
  NOR2_X2 U819 ( .A1(n1159), .A2(n1158), .ZN(n1160) );
  NOR2_X2 U820 ( .A1(n1156), .A2(n1155), .ZN(n1161) );
  NOR2_X2 U821 ( .A1(n246), .A2(n638), .ZN(n1159) );
  AOI21_X2 U822 ( .B1(n1127), .B2(n1126), .A(n1125), .ZN(n1133) );
  NAND3_X2 U823 ( .A1(n1110), .A2(n1109), .A3(n1108), .ZN(n1641) );
  NOR2_X2 U824 ( .A1(n1107), .A2(n1106), .ZN(n1108) );
  OAI21_X2 U825 ( .B1(n1115), .B2(n1114), .A(n1113), .ZN(n1122) );
  NOR2_X2 U826 ( .A1(n691), .A2(n1111), .ZN(n1115) );
  OAI21_X2 U827 ( .B1(n691), .B2(n1112), .A(b[25]), .ZN(n1113) );
  NOR2_X2 U828 ( .A1(n1120), .A2(n636), .ZN(n1121) );
  OAI21_X2 U829 ( .B1(n1089), .B2(n1088), .A(n1087), .ZN(n1097) );
  NOR2_X2 U830 ( .A1(n694), .A2(n1085), .ZN(n1089) );
  OAI21_X2 U831 ( .B1(n691), .B2(n1086), .A(b[26]), .ZN(n1087) );
  NAND3_X2 U832 ( .A1(n1084), .A2(n1083), .A3(n1082), .ZN(n1658) );
  NOR2_X2 U833 ( .A1(n1081), .A2(n1080), .ZN(n1082) );
  NOR2_X2 U834 ( .A1(n1095), .A2(n636), .ZN(n1096) );
  NAND3_X2 U835 ( .A1(n1042), .A2(n1041), .A3(n1040), .ZN(n1660) );
  AOI21_X2 U836 ( .B1(n1430), .B2(n1117), .A(n1091), .ZN(n1040) );
  NAND3_X2 U837 ( .A1(n1061), .A2(n1060), .A3(n1059), .ZN(n1681) );
  NOR2_X2 U838 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  INV_X4 U839 ( .A(n649), .ZN(n1719) );
  NOR2_X2 U840 ( .A1(n1044), .A2(n92), .ZN(n1045) );
  OAI21_X2 U841 ( .B1(a[27]), .B2(n697), .A(n692), .ZN(n1043) );
  NOR2_X2 U842 ( .A1(n1683), .A2(n636), .ZN(n1046) );
  NAND3_X2 U843 ( .A1(n991), .A2(n990), .A3(n989), .ZN(n1680) );
  NOR2_X2 U844 ( .A1(n988), .A2(n987), .ZN(n989) );
  OAI21_X2 U845 ( .B1(n1009), .B2(n1008), .A(n1007), .ZN(n1014) );
  NOR2_X2 U846 ( .A1(n691), .A2(n1005), .ZN(n1009) );
  OAI21_X2 U847 ( .B1(n691), .B2(n1006), .A(b[28]), .ZN(n1007) );
  NOR2_X2 U848 ( .A1(n1714), .A2(n634), .ZN(n993) );
  NOR2_X2 U849 ( .A1(n1704), .A2(n649), .ZN(n992) );
  NOR2_X2 U850 ( .A1(n1021), .A2(n90), .ZN(n1022) );
  OAI21_X2 U851 ( .B1(a[29]), .B2(n697), .A(n692), .ZN(n1020) );
  NOR2_X2 U852 ( .A1(n1019), .A2(n636), .ZN(n1023) );
  NOR2_X2 U853 ( .A1(n969), .A2(n634), .ZN(n974) );
  NOR2_X2 U854 ( .A1(n1728), .A2(n637), .ZN(n973) );
  OAI21_X2 U855 ( .B1(a[30]), .B2(n697), .A(n692), .ZN(n959) );
  AOI21_X2 U856 ( .B1(n1430), .B2(n983), .A(n863), .ZN(n885) );
  INV_X4 U857 ( .A(n637), .ZN(n1659) );
  NOR2_X2 U858 ( .A1(n1822), .A2(n696), .ZN(n946) );
  OAI21_X2 U859 ( .B1(n953), .B2(n692), .A(n952), .ZN(n955) );
  NOR3_X2 U860 ( .A1(n1765), .A2(n1764), .A3(n1763), .ZN(n1770) );
  NOR3_X2 U861 ( .A1(b[30]), .A2(b[9]), .A3(b[7]), .ZN(n700) );
  NAND2_X2 U862 ( .A1(n1797), .A2(n1796), .ZN(n1806) );
  NAND2_X2 U863 ( .A1(a[6]), .A2(n795), .ZN(n1593) );
  NOR2_X2 U864 ( .A1(n1840), .A2(n115), .ZN(n1209) );
  NAND2_X2 U865 ( .A1(n115), .A2(n922), .ZN(n845) );
  NOR2_X2 U866 ( .A1(n748), .A2(n1162), .ZN(n824) );
  NAND3_X2 U867 ( .A1(n1169), .A2(n1129), .A3(n1071), .ZN(n748) );
  OAI21_X2 U868 ( .B1(n660), .B2(n828), .A(n827), .ZN(n1025) );
  NOR2_X2 U869 ( .A1(n1808), .A2(n663), .ZN(n1800) );
  AOI21_X2 U870 ( .B1(n650), .B2(a[28]), .A(n1882), .ZN(n895) );
  OAI21_X2 U871 ( .B1(n806), .B2(b[0]), .A(a[0]), .ZN(n1739) );
  NAND2_X2 U872 ( .A1(n1591), .A2(n1646), .ZN(n1649) );
  NAND2_X2 U873 ( .A1(a[7]), .A2(n785), .ZN(n1596) );
  NAND2_X2 U874 ( .A1(n1695), .A2(n1668), .ZN(n815) );
  NAND2_X2 U875 ( .A1(n777), .A2(n822), .ZN(n743) );
  NAND3_X2 U876 ( .A1(n1322), .A2(n1321), .A3(n1320), .ZN(n1375) );
  NOR2_X2 U877 ( .A1(n1390), .A2(n1449), .ZN(n1322) );
  INV_X4 U878 ( .A(n681), .ZN(n1179) );
  NAND3_X2 U879 ( .A1(n873), .A2(n872), .A3(n871), .ZN(n883) );
  NOR2_X2 U880 ( .A1(n1820), .A2(n1819), .ZN(n1830) );
  AOI21_X2 U881 ( .B1(n915), .B2(a[1]), .A(n662), .ZN(n912) );
  NOR2_X2 U882 ( .A1(a[1]), .A2(n696), .ZN(n1735) );
  NOR2_X2 U883 ( .A1(a[9]), .A2(n696), .ZN(n1565) );
  OAI21_X2 U884 ( .B1(n1541), .B2(n1556), .A(n1540), .ZN(n1543) );
  NOR2_X2 U885 ( .A1(n1539), .A2(n1538), .ZN(n1540) );
  OAI21_X2 U886 ( .B1(n1296), .B2(n687), .A(n1140), .ZN(n1280) );
  OAI21_X2 U887 ( .B1(n1240), .B2(n687), .A(n1140), .ZN(n1353) );
  OAI21_X2 U888 ( .B1(n1263), .B2(n687), .A(n1140), .ZN(n1342) );
  NOR2_X2 U889 ( .A1(n246), .A2(n1405), .ZN(n1409) );
  OAI21_X2 U890 ( .B1(n1459), .B2(n1458), .A(n1457), .ZN(n1752) );
  NOR2_X2 U891 ( .A1(a[17]), .A2(n696), .ZN(n1416) );
  NAND2_X2 U892 ( .A1(n736), .A2(n1376), .ZN(n1378) );
  NOR2_X2 U893 ( .A1(n638), .A2(n1406), .ZN(n1243) );
  NOR2_X2 U894 ( .A1(n246), .A2(n1300), .ZN(n1244) );
  NOR2_X2 U895 ( .A1(n248), .A2(n1371), .ZN(n1242) );
  NOR2_X2 U896 ( .A1(n1198), .A2(n1406), .ZN(n1199) );
  NOR2_X2 U897 ( .A1(n246), .A2(n639), .ZN(n1200) );
  NOR2_X2 U898 ( .A1(n248), .A2(n1403), .ZN(n1197) );
  NOR2_X2 U899 ( .A1(n1300), .A2(n1365), .ZN(n1155) );
  NOR2_X2 U900 ( .A1(n248), .A2(n1370), .ZN(n1156) );
  NOR2_X2 U901 ( .A1(n1157), .A2(n1406), .ZN(n1158) );
  NOR2_X2 U902 ( .A1(n248), .A2(n1314), .ZN(n1107) );
  NOR2_X2 U903 ( .A1(n639), .A2(n1365), .ZN(n1106) );
  NOR2_X2 U904 ( .A1(a[25]), .A2(n696), .ZN(n1112) );
  NOR2_X2 U905 ( .A1(a[26]), .A2(n696), .ZN(n1086) );
  NOR2_X2 U906 ( .A1(n248), .A2(n1300), .ZN(n1081) );
  NOR2_X2 U907 ( .A1(n638), .A2(n1365), .ZN(n1080) );
  NOR2_X2 U908 ( .A1(n248), .A2(n1840), .ZN(n1091) );
  OAI21_X2 U909 ( .B1(n1310), .B2(n687), .A(n1140), .ZN(n1271) );
  OAI21_X2 U910 ( .B1(n1270), .B2(n687), .A(n1140), .ZN(n1212) );
  NOR2_X2 U911 ( .A1(n1198), .A2(n1365), .ZN(n1057) );
  NOR2_X2 U912 ( .A1(n248), .A2(n639), .ZN(n1058) );
  NAND3_X2 U913 ( .A1(n904), .A2(n903), .A3(n902), .ZN(n1101) );
  AOI21_X2 U914 ( .B1(b[3]), .B2(n1192), .A(n1882), .ZN(n902) );
  AOI21_X2 U915 ( .B1(n650), .B2(a[26]), .A(n1882), .ZN(n929) );
  NOR2_X2 U916 ( .A1(n1157), .A2(n1365), .ZN(n987) );
  NOR2_X2 U917 ( .A1(n248), .A2(n638), .ZN(n988) );
  NOR2_X2 U918 ( .A1(a[28]), .A2(n696), .ZN(n1006) );
  OAI21_X2 U919 ( .B1(n1282), .B2(n687), .A(n1140), .ZN(n1223) );
  INV_X4 U920 ( .A(n246), .ZN(n1427) );
  NOR2_X2 U921 ( .A1(n856), .A2(n855), .ZN(n860) );
  INV_X4 U922 ( .A(n1365), .ZN(n1430) );
  NAND3_X2 U923 ( .A1(n850), .A2(n849), .A3(n848), .ZN(n983) );
  AOI21_X2 U924 ( .B1(b[3]), .B2(n1077), .A(n1882), .ZN(n848) );
  OAI21_X2 U925 ( .B1(n837), .B2(n659), .A(n1720), .ZN(n958) );
  AOI21_X2 U926 ( .B1(n835), .B2(n1821), .A(n834), .ZN(n837) );
  AOI21_X2 U927 ( .B1(n691), .B2(n664), .A(n1839), .ZN(n1846) );
  NOR2_X2 U928 ( .A1(n642), .A2(n633), .ZN(n1841) );
  OAI21_X2 U929 ( .B1(n1604), .B2(n1603), .A(n1602), .ZN(n1605) );
  NOR2_X2 U930 ( .A1(n691), .A2(n1600), .ZN(n1604) );
  OAI21_X2 U931 ( .B1(n691), .B2(n1601), .A(b[8]), .ZN(n1602) );
  AOI211_X2 U932 ( .C1(a[12]), .C2(n1520), .A(n1519), .B(n1518), .ZN(n1533) );
  NOR2_X2 U933 ( .A1(n1514), .A2(n634), .ZN(n1519) );
  NOR2_X2 U934 ( .A1(n1517), .A2(n1516), .ZN(n1518) );
  OAI21_X2 U935 ( .B1(n1505), .B2(n1504), .A(n1503), .ZN(n1508) );
  NOR2_X2 U936 ( .A1(n691), .A2(n1501), .ZN(n1505) );
  OAI21_X2 U937 ( .B1(n691), .B2(n1502), .A(b[13]), .ZN(n1503) );
  NOR2_X2 U938 ( .A1(n1506), .A2(n634), .ZN(n1507) );
  OAI21_X2 U939 ( .B1(n1495), .B2(n680), .A(n1494), .ZN(n1498) );
  NAND2_X2 U940 ( .A1(n1389), .A2(n655), .ZN(n680) );
  AOI211_X2 U941 ( .C1(n1468), .C2(n1467), .A(n1466), .B(n1465), .ZN(n1469) );
  OAI21_X2 U942 ( .B1(n1207), .B2(n1206), .A(n1205), .ZN(n1208) );
  NOR2_X2 U943 ( .A1(n691), .A2(n1203), .ZN(n1207) );
  OAI21_X2 U944 ( .B1(n691), .B2(n1204), .A(b[23]), .ZN(n1205) );
  NOR2_X2 U945 ( .A1(n1730), .A2(n1729), .ZN(n1747) );
  OAI21_X2 U946 ( .B1(n691), .B2(n1713), .A(a[2]), .ZN(n1725) );
  AOI211_X2 U947 ( .C1(a[3]), .C2(n1702), .A(n1701), .B(n1700), .ZN(n1710) );
  NAND3_X2 U948 ( .A1(n1689), .A2(n1688), .A3(n1687), .ZN(res[4]) );
  NOR2_X2 U949 ( .A1(n1686), .A2(n1685), .ZN(n1687) );
  AOI211_X2 U950 ( .C1(a[4]), .C2(n1679), .A(n1678), .B(n1677), .ZN(n1689) );
  NOR3_X2 U951 ( .A1(n1656), .A2(n1655), .A3(n1654), .ZN(n1664) );
  NOR2_X2 U952 ( .A1(n1637), .A2(n1636), .ZN(n1645) );
  AOI211_X2 U953 ( .C1(a[7]), .C2(n1620), .A(n1619), .B(n1618), .ZN(n1631) );
  NOR2_X2 U954 ( .A1(n633), .A2(n1754), .ZN(n1586) );
  OAI21_X2 U955 ( .B1(n691), .B2(n1554), .A(a[10]), .ZN(n1562) );
  OAI21_X2 U956 ( .B1(n694), .B2(n1535), .A(a[11]), .ZN(n1551) );
  AOI211_X2 U957 ( .C1(a[14]), .C2(n1479), .A(n1478), .B(n1477), .ZN(n1493) );
  AOI21_X2 U958 ( .B1(n1844), .B2(n1488), .A(n1425), .ZN(n1447) );
  AOI211_X2 U959 ( .C1(n1444), .C2(n1467), .A(n1443), .B(n1442), .ZN(n1445) );
  AOI21_X2 U960 ( .B1(n1719), .B2(n1488), .A(n1414), .ZN(n1423) );
  NOR2_X2 U961 ( .A1(n1424), .A2(n636), .ZN(n1414) );
  AOI211_X2 U962 ( .C1(a[18]), .C2(n1363), .A(n1362), .B(n1361), .ZN(n1384) );
  AOI211_X2 U963 ( .C1(n1348), .C2(n1347), .A(n1346), .B(n1345), .ZN(n1349) );
  AOI211_X2 U964 ( .C1(a[20]), .C2(n1292), .A(n1291), .B(n1290), .ZN(n1306) );
  OAI21_X2 U965 ( .B1(n691), .B2(n1253), .A(a[21]), .ZN(n1277) );
  NOR2_X2 U966 ( .A1(n1268), .A2(n1267), .ZN(n1276) );
  AOI211_X2 U967 ( .C1(a[22]), .C2(n1231), .A(n1230), .B(n1229), .ZN(n1251) );
  AOI211_X2 U968 ( .C1(a[24]), .C2(n1151), .A(n1150), .B(n1149), .ZN(n1176) );
  AOI21_X2 U969 ( .B1(n1844), .B2(n1658), .A(n1135), .ZN(n1136) );
  AOI211_X2 U970 ( .C1(n1719), .C2(n1641), .A(n1122), .B(n1121), .ZN(n1137) );
  OAI21_X2 U971 ( .B1(n633), .B2(n1748), .A(n1134), .ZN(n1135) );
  AOI211_X2 U972 ( .C1(n1719), .C2(n1658), .A(n1097), .B(n1096), .ZN(n1098) );
  AOI211_X2 U973 ( .C1(a[27]), .C2(n1047), .A(n1046), .B(n1045), .ZN(n1065) );
  NOR2_X2 U974 ( .A1(n993), .A2(n992), .ZN(n1017) );
  AOI211_X2 U975 ( .C1(a[29]), .C2(n1024), .A(n1023), .B(n1022), .ZN(n1037) );
  OAI21_X2 U976 ( .B1(n691), .B2(n960), .A(a[30]), .ZN(n977) );
  NOR3_X2 U977 ( .A1(n974), .A2(n973), .A3(n972), .ZN(n975) );
  AOI21_X2 U978 ( .B1(n1720), .B2(n947), .A(n946), .ZN(n957) );
  INV_X4 U979 ( .A(n634), .ZN(n1844) );
  NAND2_X2 U980 ( .A1(alu_ctrl[2]), .A2(n699), .ZN(n633) );
  INV_X4 U981 ( .A(n1734), .ZN(n695) );
  NAND2_X2 U982 ( .A1(n968), .A2(n967), .ZN(n634) );
  NAND2_X2 U983 ( .A1(b[1]), .A2(b[2]), .ZN(n248) );
  AND2_X4 U984 ( .A1(n115), .A2(n1698), .ZN(n635) );
  INV_X4 U985 ( .A(n698), .ZN(n696) );
  NAND2_X2 U986 ( .A1(n954), .A2(n967), .ZN(n636) );
  NAND2_X2 U987 ( .A1(n954), .A2(b[0]), .ZN(n637) );
  AND3_X4 U988 ( .A1(n986), .A2(n1194), .A3(n668), .ZN(n638) );
  AND3_X4 U989 ( .A1(n1056), .A2(n1194), .A3(n669), .ZN(n639) );
  AND2_X4 U990 ( .A1(n699), .A2(n1817), .ZN(n640) );
  AND3_X4 U991 ( .A1(n858), .A2(n632), .A3(n857), .ZN(n641) );
  AND2_X4 U992 ( .A1(n1236), .A2(n1184), .ZN(n643) );
  INV_X4 U993 ( .A(n635), .ZN(n687) );
  AND3_X4 U994 ( .A1(n911), .A2(n924), .A3(n910), .ZN(n644) );
  INV_X4 U995 ( .A(n1711), .ZN(n694) );
  AND2_X2 U996 ( .A1(n1152), .A2(n1698), .ZN(n645) );
  AND2_X4 U997 ( .A1(n1077), .A2(n1698), .ZN(n646) );
  AND2_X4 U998 ( .A1(n1192), .A2(n1698), .ZN(n647) );
  AND2_X4 U999 ( .A1(n1103), .A2(n1698), .ZN(n648) );
  INV_X16 U1000 ( .A(alu_ctrl[3]), .ZN(n699) );
  NAND3_X2 U1001 ( .A1(b[0]), .A2(alu_ctrl[1]), .A3(n640), .ZN(n649) );
  INV_X4 U1002 ( .A(n1734), .ZN(n698) );
  AND2_X4 U1003 ( .A1(n635), .A2(n922), .ZN(n650) );
  AND2_X4 U1004 ( .A1(a[29]), .A2(n829), .ZN(n651) );
  AND2_X4 U1005 ( .A1(n1372), .A2(n1395), .ZN(n652) );
  XOR2_X2 U1006 ( .A(n740), .B(n1439), .Z(n653) );
  XOR2_X2 U1007 ( .A(n1696), .B(n1695), .Z(n654) );
  NAND2_X2 U1008 ( .A1(b[3]), .A2(n115), .ZN(n1309) );
  NAND2_X2 U1009 ( .A1(b[2]), .A2(n981), .ZN(n1365) );
  NAND2_X2 U1010 ( .A1(n1883), .A2(n981), .ZN(n1406) );
  XOR2_X2 U1011 ( .A(n1741), .B(n1740), .Z(n656) );
  INV_X4 U1012 ( .A(b[11]), .ZN(n675) );
  NOR3_X2 U1013 ( .A1(n1266), .A2(n1265), .A3(n1264), .ZN(n1555) );
  AND2_X4 U1014 ( .A1(n938), .A2(n1029), .ZN(n657) );
  AND2_X4 U1015 ( .A1(n1178), .A2(n1259), .ZN(n658) );
  AND2_X4 U1016 ( .A1(n836), .A2(a[31]), .ZN(n659) );
  AND2_X4 U1017 ( .A1(n999), .A2(n998), .ZN(n660) );
  OR2_X4 U1018 ( .A1(n644), .A2(n921), .ZN(n661) );
  AND2_X4 U1019 ( .A1(n650), .A2(a[30]), .ZN(n662) );
  NAND2_X2 U1020 ( .A1(n1578), .A2(n1386), .ZN(n1387) );
  INV_X4 U1021 ( .A(n1387), .ZN(n679) );
  OR2_X4 U1022 ( .A1(n1820), .A2(n1799), .ZN(n663) );
  NAND2_X2 U1023 ( .A1(n1717), .A2(n1693), .ZN(n1666) );
  OR2_X4 U1024 ( .A1(a[0]), .A2(b[0]), .ZN(n664) );
  INV_X4 U1025 ( .A(n248), .ZN(n690) );
  AND2_X4 U1026 ( .A1(n1659), .A2(n995), .ZN(n665) );
  AND2_X4 U1027 ( .A1(n1659), .A2(n1715), .ZN(n666) );
  INV_X4 U1028 ( .A(n633), .ZN(n1720) );
  OR2_X4 U1029 ( .A1(n644), .A2(n1309), .ZN(n667) );
  OR2_X4 U1030 ( .A1(n1295), .A2(n1309), .ZN(n668) );
  OR2_X4 U1031 ( .A1(n1308), .A2(n1309), .ZN(n669) );
  OR2_X4 U1032 ( .A1(n641), .A2(n1309), .ZN(n670) );
  INV_X4 U1033 ( .A(n1711), .ZN(n691) );
  INV_X4 U1034 ( .A(n695), .ZN(n697) );
  NOR2_X1 U1035 ( .A1(n1838), .A2(n1837), .ZN(n1839) );
  INV_X4 U1036 ( .A(n1838), .ZN(n1732) );
  AND2_X4 U1037 ( .A1(n689), .A2(n115), .ZN(n559) );
  INV_X16 U1038 ( .A(n688), .ZN(n689) );
  INV_X2 U1039 ( .A(n1775), .ZN(n1239) );
  NAND2_X2 U1040 ( .A1(n1459), .A2(n1317), .ZN(n1373) );
  INV_X2 U1041 ( .A(n740), .ZN(n739) );
  OAI211_X2 U1042 ( .C1(n1377), .C2(n671), .A(n1395), .B(n1376), .ZN(n1379) );
  INV_X1 U1043 ( .A(n1328), .ZN(n1329) );
  NAND3_X4 U1044 ( .A1(n1395), .A2(n1376), .A3(n671), .ZN(n1328) );
  AOI22_X2 U1045 ( .A1(n1496), .A2(n1497), .B1(n1498), .B2(n1499), .ZN(n672)
         );
  INV_X4 U1046 ( .A(n672), .ZN(n1753) );
  INV_X4 U1047 ( .A(n1496), .ZN(n1499) );
  XNOR2_X2 U1048 ( .A(n673), .B(n1330), .ZN(n1790) );
  AND2_X2 U1049 ( .A1(n1379), .A2(n1378), .ZN(n673) );
  NAND2_X4 U1050 ( .A1(alu_ctrl[1]), .A2(n699), .ZN(n760) );
  NAND2_X2 U1051 ( .A1(n1262), .A2(n677), .ZN(n1777) );
  INV_X1 U1052 ( .A(n1254), .ZN(n1255) );
  INV_X16 U1053 ( .A(alu_ctrl[1]), .ZN(n949) );
  NAND2_X4 U1054 ( .A1(a[11]), .A2(n762), .ZN(n1527) );
  AND4_X2 U1055 ( .A1(n676), .A2(n674), .A3(n1516), .A4(n675), .ZN(n587) );
  NOR3_X2 U1056 ( .A1(b[14]), .A2(b[15]), .A3(b[13]), .ZN(n676) );
  OAI21_X2 U1057 ( .B1(n1133), .B2(n1132), .A(n1131), .ZN(n1748) );
  NOR2_X2 U1058 ( .A1(alu_ctrl[0]), .A2(n1833), .ZN(n1834) );
  NAND2_X1 U1059 ( .A1(n1234), .A2(n1235), .ZN(n677) );
  NAND2_X4 U1060 ( .A1(n1575), .A2(n797), .ZN(n1577) );
  XNOR2_X2 U1061 ( .A(n1004), .B(n1003), .ZN(n678) );
  INV_X1 U1062 ( .A(n1776), .ZN(n1074) );
  NAND2_X4 U1063 ( .A1(n733), .A2(n699), .ZN(n802) );
  INV_X1 U1064 ( .A(n1797), .ZN(n1052) );
  NAND2_X1 U1065 ( .A1(b[1]), .A2(n963), .ZN(n884) );
  NAND2_X1 U1066 ( .A1(n1432), .A2(n1075), .ZN(n1084) );
  NAND2_X1 U1067 ( .A1(n1075), .A2(n1427), .ZN(n991) );
  NAND2_X4 U1068 ( .A1(n681), .A2(n1177), .ZN(n1167) );
  NAND2_X4 U1069 ( .A1(n1261), .A2(n1236), .ZN(n1238) );
  OAI22_X4 U1070 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n800) );
  OAI21_X2 U1071 ( .B1(n1030), .B2(n1029), .A(n1826), .ZN(n1796) );
  AOI21_X2 U1072 ( .B1(n1233), .B2(n1183), .A(n1182), .ZN(n1187) );
  NAND2_X4 U1073 ( .A1(n1190), .A2(n1189), .ZN(n1191) );
  NOR2_X2 U1074 ( .A1(n633), .A2(n1777), .ZN(n1268) );
  NAND2_X2 U1075 ( .A1(n1373), .A2(n1375), .ZN(n1333) );
  XNOR2_X2 U1076 ( .A(n799), .B(n800), .ZN(n1717) );
  NOR2_X1 U1077 ( .A1(n678), .A2(n1806), .ZN(n1801) );
  XNOR2_X1 U1078 ( .A(n1639), .B(n1638), .ZN(n1765) );
  NAND2_X2 U1079 ( .A1(n1649), .A2(n1592), .ZN(n1639) );
  NAND2_X2 U1080 ( .A1(n1163), .A2(n1256), .ZN(n1168) );
  INV_X4 U1081 ( .A(n684), .ZN(n685) );
  INV_X8 U1082 ( .A(n684), .ZN(n686) );
  INV_X8 U1083 ( .A(n1756), .ZN(n684) );
  INV_X2 U1084 ( .A(n1668), .ZN(n1669) );
  NAND2_X2 U1085 ( .A1(n1668), .A2(n1667), .ZN(n817) );
  NAND2_X4 U1086 ( .A1(n1234), .A2(n1235), .ZN(n1261) );
  OAI21_X2 U1087 ( .B1(n1594), .B2(n1638), .A(n1593), .ZN(n1621) );
  NAND2_X4 U1088 ( .A1(a[5]), .A2(n791), .ZN(n1592) );
  OAI22_X4 U1089 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n790) );
  NAND3_X2 U1090 ( .A1(n882), .A2(n881), .A3(n880), .ZN(n1075) );
  AOI21_X2 U1091 ( .B1(b[3]), .B2(n1152), .A(n683), .ZN(n880) );
  INV_X1 U1092 ( .A(n1167), .ZN(n1126) );
  NAND3_X4 U1093 ( .A1(n821), .A2(n822), .A3(n823), .ZN(n681) );
  NAND3_X2 U1094 ( .A1(n823), .A2(n822), .A3(n821), .ZN(n1257) );
  NAND4_X4 U1095 ( .A1(n1257), .A2(n1177), .A3(n1256), .A4(n824), .ZN(n937) );
  NAND3_X2 U1096 ( .A1(n1256), .A2(n681), .A3(n1255), .ZN(n1294) );
  NOR3_X4 U1097 ( .A1(n1871), .A2(n1870), .A3(n1869), .ZN(n1873) );
  NAND2_X4 U1098 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X4 U1099 ( .A1(n1799), .A2(n699), .ZN(n783) );
  AOI22_X1 U1100 ( .A1(n1716), .A2(n1500), .B1(n1720), .B2(n1790), .ZN(n1381)
         );
  NOR2_X4 U1101 ( .A1(n1790), .A2(n1789), .ZN(n1791) );
  NAND2_X1 U1102 ( .A1(n1692), .A2(n1691), .ZN(n1718) );
  INV_X1 U1103 ( .A(n1794), .ZN(n947) );
  INV_X1 U1104 ( .A(n1796), .ZN(n1031) );
  NAND3_X1 U1105 ( .A1(n1812), .A2(n1811), .A3(alu_ctrl[0]), .ZN(n1813) );
  NAND2_X4 U1106 ( .A1(n742), .A2(n1335), .ZN(n822) );
  OAI22_X4 U1107 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n738) );
  NAND4_X4 U1108 ( .A1(n1693), .A2(n1691), .A3(n1668), .A4(n1692), .ZN(n816)
         );
  NOR2_X1 U1109 ( .A1(n1727), .A2(n637), .ZN(n1730) );
  OAI211_X2 U1110 ( .C1(n1396), .C2(n671), .A(n1395), .B(n1394), .ZN(n1397) );
  NOR2_X2 U1111 ( .A1(n1877), .A2(n1876), .ZN(zf) );
  NOR2_X2 U1112 ( .A1(n1818), .A2(n1817), .ZN(n1835) );
  INV_X8 U1113 ( .A(n1811), .ZN(n1808) );
  NAND2_X4 U1114 ( .A1(alu_ctrl[0]), .A2(n949), .ZN(n733) );
  INV_X4 U1115 ( .A(n1480), .ZN(n1484) );
  NAND3_X2 U1116 ( .A1(n630), .A2(n1448), .A3(n679), .ZN(n1480) );
  AOI211_X1 U1117 ( .C1(n1720), .C2(n678), .A(n1014), .B(n666), .ZN(n1015) );
  OAI22_X2 U1118 ( .A1(n1051), .A2(n1050), .B1(n1049), .B2(n1048), .ZN(n1797)
         );
  INV_X2 U1119 ( .A(n1050), .ZN(n1048) );
  NAND2_X4 U1120 ( .A1(alu_ctrl[1]), .A2(n699), .ZN(n784) );
  NAND3_X1 U1121 ( .A1(alu_ctrl[3]), .A2(alu_ctrl[1]), .A3(n945), .ZN(n1734)
         );
  NAND3_X1 U1122 ( .A1(alu_ctrl[3]), .A2(n1817), .A3(n949), .ZN(n1838) );
  OAI22_X1 U1123 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n714) );
  OAI22_X1 U1124 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n731) );
  OAI22_X1 U1125 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n805) );
  INV_X1 U1126 ( .A(n1481), .ZN(n1450) );
  INV_X2 U1127 ( .A(n1768), .ZN(n1487) );
  INV_X2 U1128 ( .A(n1577), .ZN(n1579) );
  NOR2_X2 U1129 ( .A1(n1556), .A2(n1385), .ZN(n779) );
  INV_X2 U1130 ( .A(n1556), .ZN(n1448) );
  NAND2_X1 U1131 ( .A1(n1844), .A2(n1544), .ZN(n1350) );
  NAND2_X1 U1132 ( .A1(n1719), .A2(n1544), .ZN(n1304) );
  NAND2_X1 U1133 ( .A1(n1722), .A2(n1544), .ZN(n1531) );
  NOR2_X2 U1134 ( .A1(n1548), .A2(n1547), .ZN(n1549) );
  AOI21_X1 U1135 ( .B1(n559), .B2(a[9]), .A(n1882), .ZN(n582) );
  AOI21_X1 U1136 ( .B1(n559), .B2(a[8]), .A(n683), .ZN(n564) );
  AOI21_X1 U1137 ( .B1(n559), .B2(a[13]), .A(n683), .ZN(n585) );
  AOI21_X1 U1138 ( .B1(n559), .B2(a[12]), .A(n683), .ZN(n558) );
  AOI21_X1 U1139 ( .B1(n559), .B2(a[11]), .A(n683), .ZN(n577) );
  AOI21_X1 U1140 ( .B1(n559), .B2(a[15]), .A(n1882), .ZN(n580) );
  AOI21_X1 U1141 ( .B1(n559), .B2(a[10]), .A(n1882), .ZN(n570) );
  AOI21_X1 U1142 ( .B1(n559), .B2(a[14]), .A(n1882), .ZN(n573) );
  NAND2_X4 U1143 ( .A1(n1574), .A2(n1573), .ZN(n1646) );
  NAND3_X1 U1144 ( .A1(n1576), .A2(n1646), .A3(n1575), .ZN(n1582) );
  INV_X1 U1145 ( .A(n1646), .ZN(n1648) );
  XNOR2_X2 U1146 ( .A(n1598), .B(n1597), .ZN(n1749) );
  NAND2_X4 U1147 ( .A1(n1814), .A2(n1813), .ZN(n1815) );
  OAI21_X2 U1148 ( .B1(n1480), .B2(n1456), .A(n1455), .ZN(n1458) );
  NAND2_X4 U1149 ( .A1(n1030), .A2(n1029), .ZN(n1826) );
  NAND4_X4 U1150 ( .A1(n817), .A2(n816), .A3(n1672), .A4(n815), .ZN(n1573) );
  NAND2_X4 U1151 ( .A1(n1794), .A2(n1822), .ZN(n1811) );
  OAI21_X1 U1152 ( .B1(n807), .B2(n1757), .A(n1739), .ZN(n1741) );
  NAND2_X4 U1153 ( .A1(n1757), .A2(n1739), .ZN(n809) );
  NAND2_X4 U1154 ( .A1(n1178), .A2(n1177), .ZN(n1254) );
  NAND2_X4 U1155 ( .A1(n1326), .A2(n745), .ZN(n1177) );
  INV_X2 U1156 ( .A(n1524), .ZN(n1539) );
  NOR2_X1 U1157 ( .A1(n1481), .A2(n1496), .ZN(n1483) );
  NAND2_X4 U1158 ( .A1(n1389), .A2(n1388), .ZN(n1481) );
  NAND2_X4 U1159 ( .A1(n1524), .A2(n1527), .ZN(n1388) );
  OAI21_X1 U1160 ( .B1(n1494), .B2(n1496), .A(n1452), .ZN(n1482) );
  INV_X2 U1161 ( .A(n1294), .ZN(n1260) );
  NOR2_X1 U1162 ( .A1(n1803), .A2(n633), .ZN(n972) );
  NAND2_X1 U1163 ( .A1(n1808), .A2(n1803), .ZN(n1795) );
  OAI21_X2 U1164 ( .B1(n831), .B2(n1000), .A(n830), .ZN(n970) );
  NAND2_X1 U1165 ( .A1(n1067), .A2(n1256), .ZN(n1070) );
  INV_X8 U1166 ( .A(n1256), .ZN(n1181) );
  NAND3_X2 U1167 ( .A1(n1753), .A2(n1752), .A3(n1751), .ZN(n1772) );
  NOR4_X4 U1168 ( .A1(n1774), .A2(n1773), .A3(n1772), .A4(n1771), .ZN(n1793)
         );
  NAND3_X1 U1169 ( .A1(n1693), .A2(n1691), .A3(n1692), .ZN(n1670) );
  OAI21_X1 U1170 ( .B1(n1694), .B2(n1717), .A(n1693), .ZN(n1696) );
  NAND2_X4 U1171 ( .A1(n1000), .A2(n999), .ZN(n1050) );
  NAND2_X1 U1172 ( .A1(n1880), .A2(n1879), .ZN(res[0]) );
  NOR2_X2 U1173 ( .A1(n1807), .A2(n1795), .ZN(n1802) );
  INV_X8 U1174 ( .A(n1807), .ZN(n1809) );
  NOR3_X1 U1175 ( .A1(n1391), .A2(n1390), .A3(n671), .ZN(n1392) );
  NAND3_X2 U1176 ( .A1(n936), .A2(n937), .A3(n1072), .ZN(n1000) );
  NAND2_X4 U1177 ( .A1(n937), .A2(n936), .ZN(n1027) );
  INV_X2 U1178 ( .A(n1319), .ZN(n1320) );
  NAND2_X1 U1179 ( .A1(n679), .A2(n630), .ZN(n1583) );
  AOI22_X4 U1180 ( .A1(n772), .A2(n771), .B1(a[12]), .B2(n770), .ZN(n1494) );
  NAND4_X4 U1181 ( .A1(n777), .A2(n1459), .A3(n822), .A4(n1317), .ZN(n1256) );
  NAND2_X4 U1182 ( .A1(n733), .A2(n699), .ZN(n1756) );
  INV_X8 U1183 ( .A(n839), .ZN(n922) );
  INV_X4 U1184 ( .A(b[19]), .ZN(n100) );
  INV_X4 U1185 ( .A(b[21]), .ZN(n98) );
  INV_X4 U1186 ( .A(b[22]), .ZN(n97) );
  INV_X4 U1187 ( .A(b[26]), .ZN(n93) );
  INV_X4 U1188 ( .A(b[27]), .ZN(n92) );
  INV_X4 U1189 ( .A(b[28]), .ZN(n91) );
  INV_X4 U1190 ( .A(b[29]), .ZN(n90) );
  INV_X4 U1191 ( .A(b[31]), .ZN(n953) );
  NAND3_X2 U1192 ( .A1(n587), .A2(n953), .A3(n700), .ZN(n703) );
  NAND4_X2 U1193 ( .A1(n588), .A2(n589), .A3(n109), .A4(n701), .ZN(n702) );
  OR2_X2 U1194 ( .A1(n703), .A2(n702), .ZN(n586) );
  INV_X4 U1195 ( .A(n586), .ZN(n838) );
  NAND2_X2 U1196 ( .A1(a[31]), .A2(alu_ctrl[0]), .ZN(n1840) );
  INV_X4 U1197 ( .A(b[2]), .ZN(n1883) );
  INV_X4 U1198 ( .A(b[30]), .ZN(n704) );
  XNOR2_X2 U1199 ( .A(n686), .B(n704), .ZN(n832) );
  INV_X4 U1200 ( .A(a[30]), .ZN(n705) );
  XNOR2_X2 U1201 ( .A(n832), .B(n705), .ZN(n1824) );
  XNOR2_X2 U1202 ( .A(n686), .B(n92), .ZN(n707) );
  INV_X4 U1203 ( .A(a[27]), .ZN(n706) );
  XNOR2_X2 U1204 ( .A(n707), .B(n706), .ZN(n1051) );
  INV_X4 U1205 ( .A(n1051), .ZN(n1049) );
  NAND2_X2 U1206 ( .A1(a[27]), .A2(n707), .ZN(n998) );
  NAND2_X2 U1207 ( .A1(n1049), .A2(n998), .ZN(n1001) );
  XNOR2_X2 U1208 ( .A(n685), .B(n91), .ZN(n826) );
  INV_X4 U1209 ( .A(a[28]), .ZN(n1008) );
  XNOR2_X2 U1210 ( .A(n826), .B(n1008), .ZN(n1003) );
  NAND2_X2 U1211 ( .A1(n1001), .A2(n1003), .ZN(n828) );
  INV_X4 U1212 ( .A(n828), .ZN(n709) );
  XNOR2_X2 U1213 ( .A(n686), .B(n90), .ZN(n829) );
  INV_X4 U1214 ( .A(a[29]), .ZN(n708) );
  XNOR2_X2 U1215 ( .A(n829), .B(n708), .ZN(n1029) );
  NAND2_X2 U1216 ( .A1(n709), .A2(n1029), .ZN(n831) );
  XNOR2_X2 U1217 ( .A(n686), .B(n1147), .ZN(n725) );
  NAND2_X2 U1218 ( .A1(a[24]), .A2(n725), .ZN(n1129) );
  INV_X4 U1219 ( .A(n1129), .ZN(n1066) );
  XOR2_X2 U1220 ( .A(n686), .B(b[23]), .Z(n710) );
  NAND2_X2 U1221 ( .A1(a[23]), .A2(n710), .ZN(n1169) );
  INV_X4 U1222 ( .A(n1169), .ZN(n727) );
  XNOR2_X2 U1223 ( .A(n686), .B(n98), .ZN(n711) );
  NAND2_X2 U1224 ( .A1(a[21]), .A2(n711), .ZN(n1236) );
  XNOR2_X2 U1225 ( .A(n685), .B(n97), .ZN(n712) );
  NAND2_X2 U1226 ( .A1(a[22]), .A2(n712), .ZN(n1184) );
  XNOR2_X2 U1227 ( .A(b[20]), .B(n714), .ZN(n713) );
  NAND2_X2 U1228 ( .A1(a[20]), .A2(n713), .ZN(n1259) );
  INV_X4 U1229 ( .A(n1259), .ZN(n719) );
  XNOR2_X2 U1230 ( .A(a[20]), .B(b[20]), .ZN(n715) );
  XNOR2_X2 U1231 ( .A(n715), .B(n714), .ZN(n1293) );
  INV_X4 U1232 ( .A(n1293), .ZN(n718) );
  XNOR2_X2 U1233 ( .A(a[21]), .B(b[21]), .ZN(n716) );
  XNOR2_X2 U1234 ( .A(n731), .B(n716), .ZN(n1258) );
  INV_X4 U1235 ( .A(n1258), .ZN(n717) );
  OAI21_X4 U1236 ( .B1(n719), .B2(n718), .A(n717), .ZN(n1232) );
  INV_X4 U1237 ( .A(n1184), .ZN(n722) );
  XOR2_X2 U1238 ( .A(a[22]), .B(b[22]), .Z(n720) );
  XNOR2_X2 U1239 ( .A(n807), .B(n720), .ZN(n1237) );
  XOR2_X2 U1240 ( .A(a[23]), .B(b[23]), .Z(n721) );
  XNOR2_X2 U1241 ( .A(n807), .B(n721), .ZN(n1165) );
  OAI21_X4 U1242 ( .B1(n722), .B2(n1237), .A(n1165), .ZN(n723) );
  AOI21_X4 U1243 ( .B1(n643), .B2(n1232), .A(n723), .ZN(n726) );
  INV_X4 U1244 ( .A(a[24]), .ZN(n724) );
  XNOR2_X2 U1245 ( .A(n725), .B(n724), .ZN(n1170) );
  OAI21_X4 U1246 ( .B1(n727), .B2(n726), .A(n1170), .ZN(n1125) );
  INV_X4 U1247 ( .A(n1125), .ZN(n729) );
  INV_X4 U1248 ( .A(b[25]), .ZN(n728) );
  XNOR2_X2 U1249 ( .A(n686), .B(n728), .ZN(n730) );
  INV_X4 U1250 ( .A(a[25]), .ZN(n1114) );
  XNOR2_X2 U1251 ( .A(n730), .B(n1114), .ZN(n1128) );
  OAI21_X4 U1252 ( .B1(n1066), .B2(n729), .A(n1128), .ZN(n1068) );
  NAND2_X2 U1253 ( .A1(a[25]), .A2(n730), .ZN(n1071) );
  NAND2_X2 U1254 ( .A1(n1068), .A2(n1071), .ZN(n936) );
  XNOR2_X2 U1255 ( .A(n685), .B(n93), .ZN(n825) );
  INV_X4 U1256 ( .A(a[26]), .ZN(n1088) );
  XNOR2_X2 U1257 ( .A(n825), .B(n1088), .ZN(n1072) );
  XNOR2_X2 U1258 ( .A(n731), .B(n100), .ZN(n746) );
  INV_X4 U1259 ( .A(a[19]), .ZN(n1340) );
  XNOR2_X2 U1260 ( .A(n746), .B(n1340), .ZN(n1334) );
  INV_X4 U1261 ( .A(n1334), .ZN(n777) );
  XOR2_X2 U1262 ( .A(a[17]), .B(b[17]), .Z(n732) );
  XNOR2_X2 U1263 ( .A(n684), .B(n732), .ZN(n1398) );
  INV_X4 U1264 ( .A(n1398), .ZN(n736) );
  INV_X4 U1265 ( .A(b[17]), .ZN(n734) );
  XNOR2_X2 U1266 ( .A(n1756), .B(n734), .ZN(n735) );
  NAND2_X2 U1267 ( .A1(a[17]), .A2(n735), .ZN(n1376) );
  XOR2_X2 U1268 ( .A(a[18]), .B(b[18]), .Z(n737) );
  XNOR2_X2 U1269 ( .A(n807), .B(n737), .ZN(n1380) );
  INV_X4 U1270 ( .A(b[16]), .ZN(n1440) );
  XNOR2_X2 U1271 ( .A(n738), .B(n1440), .ZN(n740) );
  NAND2_X2 U1272 ( .A1(a[16]), .A2(n739), .ZN(n1395) );
  INV_X4 U1273 ( .A(a[16]), .ZN(n1439) );
  NAND3_X4 U1274 ( .A1(n1378), .A2(n1380), .A3(n1328), .ZN(n742) );
  XNOR2_X2 U1275 ( .A(n686), .B(n1359), .ZN(n741) );
  NAND2_X2 U1276 ( .A1(a[18]), .A2(n741), .ZN(n1335) );
  INV_X4 U1277 ( .A(n743), .ZN(n1326) );
  INV_X4 U1278 ( .A(b[15]), .ZN(n1463) );
  XNOR2_X2 U1279 ( .A(n686), .B(n1463), .ZN(n744) );
  NAND2_X2 U1280 ( .A1(a[15]), .A2(n744), .ZN(n1372) );
  INV_X4 U1281 ( .A(n746), .ZN(n747) );
  NAND2_X2 U1282 ( .A1(a[19]), .A2(n747), .ZN(n1178) );
  NAND2_X2 U1283 ( .A1(n658), .A2(n643), .ZN(n1162) );
  XOR2_X2 U1284 ( .A(b[15]), .B(a[15]), .Z(n749) );
  XNOR2_X2 U1285 ( .A(n684), .B(n749), .ZN(n1459) );
  XOR2_X2 U1286 ( .A(b[14]), .B(a[14]), .Z(n750) );
  XNOR2_X2 U1287 ( .A(n684), .B(n750), .ZN(n1454) );
  INV_X4 U1288 ( .A(n1454), .ZN(n1486) );
  OAI22_X2 U1289 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n752) );
  INV_X4 U1290 ( .A(b[13]), .ZN(n751) );
  XNOR2_X2 U1291 ( .A(n752), .B(n751), .ZN(n773) );
  INV_X4 U1292 ( .A(n773), .ZN(n753) );
  NAND2_X2 U1293 ( .A1(a[13]), .A2(n753), .ZN(n1452) );
  INV_X4 U1294 ( .A(alu_ctrl[0]), .ZN(n1799) );
  NAND2_X2 U1295 ( .A1(n784), .A2(n783), .ZN(n769) );
  XNOR2_X2 U1296 ( .A(b[12]), .B(a[12]), .ZN(n754) );
  XNOR2_X2 U1297 ( .A(n769), .B(n754), .ZN(n1528) );
  INV_X4 U1298 ( .A(n1528), .ZN(n1389) );
  NOR2_X4 U1299 ( .A1(alu_ctrl[3]), .A2(alu_ctrl[0]), .ZN(n755) );
  INV_X4 U1300 ( .A(n755), .ZN(n759) );
  INV_X4 U1301 ( .A(a[11]), .ZN(n756) );
  XNOR2_X2 U1302 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X2 U1303 ( .A(n758), .B(n675), .ZN(n1524) );
  NAND2_X2 U1304 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X4 U1305 ( .A(n761), .ZN(n814) );
  XNOR2_X2 U1306 ( .A(n814), .B(n675), .ZN(n762) );
  INV_X4 U1307 ( .A(n1481), .ZN(n772) );
  XNOR2_X2 U1308 ( .A(b[10]), .B(a[10]), .ZN(n763) );
  OAI22_X2 U1309 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n767) );
  XNOR2_X2 U1310 ( .A(n763), .B(n767), .ZN(n1556) );
  NAND2_X2 U1311 ( .A1(n784), .A2(n783), .ZN(n765) );
  INV_X4 U1312 ( .A(b[9]), .ZN(n764) );
  XNOR2_X2 U1313 ( .A(n765), .B(n764), .ZN(n778) );
  INV_X4 U1314 ( .A(n778), .ZN(n766) );
  NAND2_X2 U1315 ( .A1(a[9]), .A2(n766), .ZN(n1523) );
  XNOR2_X2 U1316 ( .A(b[10]), .B(n800), .ZN(n768) );
  NAND2_X2 U1317 ( .A1(a[10]), .A2(n768), .ZN(n1525) );
  OAI211_X2 U1318 ( .C1(n1556), .C2(n1523), .A(n1525), .B(n1527), .ZN(n771) );
  XNOR2_X2 U1319 ( .A(n769), .B(b[12]), .ZN(n770) );
  INV_X4 U1320 ( .A(a[13]), .ZN(n1504) );
  XNOR2_X2 U1321 ( .A(n773), .B(n1504), .ZN(n1496) );
  XNOR2_X2 U1322 ( .A(n685), .B(b[14]), .ZN(n775) );
  INV_X4 U1323 ( .A(a[14]), .ZN(n774) );
  INV_X4 U1324 ( .A(n1453), .ZN(n776) );
  INV_X4 U1325 ( .A(a[9]), .ZN(n1567) );
  XNOR2_X2 U1326 ( .A(n778), .B(n1567), .ZN(n1385) );
  NAND2_X2 U1327 ( .A1(n779), .A2(n1450), .ZN(n1318) );
  XNOR2_X2 U1328 ( .A(n686), .B(n109), .ZN(n781) );
  NAND2_X2 U1329 ( .A1(a[8]), .A2(n781), .ZN(n1581) );
  XNOR2_X2 U1330 ( .A(n686), .B(n115), .ZN(n782) );
  NAND2_X2 U1331 ( .A1(a[4]), .A2(n782), .ZN(n1574) );
  XNOR2_X2 U1332 ( .A(b[7]), .B(n787), .ZN(n785) );
  INV_X4 U1333 ( .A(n1596), .ZN(n789) );
  XNOR2_X2 U1334 ( .A(a[7]), .B(b[7]), .ZN(n786) );
  XNOR2_X2 U1335 ( .A(n787), .B(n786), .ZN(n1622) );
  INV_X4 U1336 ( .A(n1622), .ZN(n1595) );
  INV_X4 U1337 ( .A(a[8]), .ZN(n1603) );
  XNOR2_X2 U1338 ( .A(n802), .B(n1603), .ZN(n788) );
  XNOR2_X2 U1339 ( .A(n788), .B(n109), .ZN(n1597) );
  OAI21_X4 U1340 ( .B1(n789), .B2(n1595), .A(n1597), .ZN(n820) );
  INV_X4 U1341 ( .A(n820), .ZN(n1575) );
  XNOR2_X2 U1342 ( .A(n790), .B(n112), .ZN(n818) );
  INV_X4 U1343 ( .A(n818), .ZN(n791) );
  INV_X4 U1344 ( .A(n1592), .ZN(n794) );
  XNOR2_X2 U1345 ( .A(a[6]), .B(b[6]), .ZN(n793) );
  OAI22_X2 U1346 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n792) );
  XNOR2_X2 U1347 ( .A(n793), .B(n792), .ZN(n1638) );
  INV_X4 U1348 ( .A(n1638), .ZN(n819) );
  NAND2_X2 U1349 ( .A1(n794), .A2(n819), .ZN(n796) );
  XOR2_X2 U1350 ( .A(n1756), .B(b[6]), .Z(n795) );
  NAND3_X2 U1351 ( .A1(n796), .A2(n1596), .A3(n1593), .ZN(n797) );
  XNOR2_X2 U1352 ( .A(n814), .B(n1698), .ZN(n798) );
  NAND2_X2 U1353 ( .A1(a[3]), .A2(n798), .ZN(n1668) );
  XNOR2_X2 U1354 ( .A(a[2]), .B(b[2]), .ZN(n799) );
  XNOR2_X2 U1355 ( .A(b[2]), .B(n800), .ZN(n801) );
  INV_X4 U1356 ( .A(b[1]), .ZN(n981) );
  XNOR2_X2 U1357 ( .A(n1756), .B(n981), .ZN(n803) );
  NAND2_X2 U1358 ( .A1(a[1]), .A2(n803), .ZN(n1691) );
  XNOR2_X2 U1359 ( .A(a[1]), .B(b[1]), .ZN(n804) );
  XNOR2_X2 U1360 ( .A(n805), .B(n804), .ZN(n1740) );
  INV_X4 U1361 ( .A(n1740), .ZN(n811) );
  INV_X4 U1362 ( .A(n686), .ZN(n807) );
  INV_X4 U1363 ( .A(n767), .ZN(n806) );
  NAND2_X2 U1364 ( .A1(n684), .A2(n1739), .ZN(n810) );
  XNOR2_X2 U1365 ( .A(a[0]), .B(b[0]), .ZN(n1832) );
  OAI22_X2 U1366 ( .A1(alu_ctrl[3]), .A2(n949), .B1(alu_ctrl[3]), .B2(
        alu_ctrl[0]), .ZN(n808) );
  XNOR2_X2 U1367 ( .A(n1832), .B(n808), .ZN(n1757) );
  NAND3_X4 U1368 ( .A1(n811), .A2(n810), .A3(n809), .ZN(n1692) );
  XOR2_X2 U1369 ( .A(b[4]), .B(a[4]), .Z(n812) );
  XNOR2_X2 U1370 ( .A(n684), .B(n812), .ZN(n1672) );
  XOR2_X2 U1371 ( .A(a[3]), .B(b[3]), .Z(n813) );
  XNOR2_X2 U1372 ( .A(n814), .B(n813), .ZN(n1695) );
  XNOR2_X2 U1373 ( .A(n818), .B(n76), .ZN(n1647) );
  INV_X4 U1374 ( .A(n1647), .ZN(n1591) );
  NAND2_X2 U1375 ( .A1(n1591), .A2(n819), .ZN(n1572) );
  OAI211_X2 U1376 ( .C1(n820), .C2(n1572), .A(n1581), .B(n1577), .ZN(n1386) );
  NAND2_X2 U1377 ( .A1(n1522), .A2(n1386), .ZN(n1319) );
  INV_X4 U1378 ( .A(n1319), .ZN(n821) );
  NAND2_X2 U1379 ( .A1(a[26]), .A2(n825), .ZN(n999) );
  NAND2_X2 U1380 ( .A1(a[28]), .A2(n826), .ZN(n827) );
  NAND2_X2 U1381 ( .A1(n1824), .A2(n970), .ZN(n835) );
  NAND2_X2 U1382 ( .A1(a[30]), .A2(n832), .ZN(n1821) );
  XNOR2_X2 U1383 ( .A(n686), .B(n953), .ZN(n836) );
  INV_X4 U1384 ( .A(a[31]), .ZN(n833) );
  XNOR2_X2 U1385 ( .A(n836), .B(n833), .ZN(n1819) );
  INV_X4 U1386 ( .A(n1819), .ZN(n834) );
  INV_X4 U1387 ( .A(n958), .ZN(cf) );
  NAND2_X2 U1388 ( .A1(alu_ctrl[1]), .A2(n838), .ZN(n839) );
  NAND2_X2 U1389 ( .A1(n635), .A2(n689), .ZN(n855) );
  INV_X4 U1390 ( .A(n855), .ZN(n915) );
  AOI22_X2 U1391 ( .A1(n650), .A2(a[27]), .B1(n915), .B2(a[4]), .ZN(n850) );
  NAND2_X2 U1392 ( .A1(b[4]), .A2(n1698), .ZN(n921) );
  INV_X4 U1393 ( .A(n921), .ZN(n842) );
  NAND2_X2 U1394 ( .A1(n689), .A2(a[20]), .ZN(n841) );
  NAND2_X2 U1395 ( .A1(n922), .A2(a[11]), .ZN(n840) );
  NAND3_X2 U1396 ( .A1(n841), .A2(n924), .A3(n840), .ZN(n1078) );
  NAND2_X2 U1397 ( .A1(n842), .A2(n1078), .ZN(n849) );
  NAND2_X2 U1398 ( .A1(n689), .A2(a[28]), .ZN(n844) );
  NAND2_X2 U1399 ( .A1(n922), .A2(a[3]), .ZN(n843) );
  NAND3_X2 U1400 ( .A1(n844), .A2(n924), .A3(n843), .ZN(n994) );
  NAND2_X2 U1401 ( .A1(n994), .A2(b[4]), .ZN(n847) );
  INV_X4 U1402 ( .A(n845), .ZN(n918) );
  NAND2_X2 U1403 ( .A1(n918), .A2(a[19]), .ZN(n846) );
  NAND3_X2 U1404 ( .A1(n558), .A2(n847), .A3(n846), .ZN(n1077) );
  NAND2_X2 U1405 ( .A1(n689), .A2(a[24]), .ZN(n852) );
  NAND2_X2 U1406 ( .A1(n922), .A2(a[7]), .ZN(n851) );
  NAND3_X2 U1407 ( .A1(n852), .A2(n632), .A3(n851), .ZN(n1139) );
  NAND2_X2 U1408 ( .A1(n1139), .A2(b[4]), .ZN(n854) );
  NAND2_X2 U1409 ( .A1(n918), .A2(a[23]), .ZN(n853) );
  NAND3_X2 U1410 ( .A1(n564), .A2(n854), .A3(n853), .ZN(n961) );
  INV_X4 U1411 ( .A(a[0]), .ZN(n856) );
  NAND2_X2 U1412 ( .A1(n689), .A2(a[16]), .ZN(n858) );
  NAND2_X2 U1413 ( .A1(n922), .A2(a[15]), .ZN(n857) );
  AOI211_X2 U1414 ( .C1(b[3]), .C2(n961), .A(n860), .B(n859), .ZN(n862) );
  AOI22_X2 U1415 ( .A1(n650), .A2(a[31]), .B1(n1882), .B2(n635), .ZN(n861) );
  AOI21_X2 U1416 ( .B1(n862), .B2(n861), .A(n1406), .ZN(n863) );
  AOI22_X2 U1417 ( .A1(n650), .A2(a[29]), .B1(n915), .B2(a[2]), .ZN(n873) );
  INV_X4 U1418 ( .A(n921), .ZN(n866) );
  NAND2_X2 U1419 ( .A1(n689), .A2(a[18]), .ZN(n865) );
  NAND2_X2 U1420 ( .A1(n922), .A2(a[13]), .ZN(n864) );
  NAND3_X2 U1421 ( .A1(n865), .A2(n924), .A3(n864), .ZN(n985) );
  NAND2_X2 U1422 ( .A1(n866), .A2(n985), .ZN(n872) );
  NAND2_X2 U1423 ( .A1(n689), .A2(a[26]), .ZN(n868) );
  NAND2_X2 U1424 ( .A1(n922), .A2(a[5]), .ZN(n867) );
  NAND3_X2 U1425 ( .A1(n868), .A2(n682), .A3(n867), .ZN(n1090) );
  NAND2_X2 U1426 ( .A1(n1090), .A2(b[4]), .ZN(n870) );
  NAND2_X2 U1427 ( .A1(n918), .A2(a[21]), .ZN(n869) );
  NAND3_X2 U1428 ( .A1(n570), .A2(n870), .A3(n869), .ZN(n984) );
  AOI22_X2 U1429 ( .A1(n650), .A2(a[25]), .B1(n915), .B2(a[6]), .ZN(n882) );
  NAND2_X2 U1430 ( .A1(n689), .A2(a[22]), .ZN(n875) );
  NAND2_X2 U1431 ( .A1(n922), .A2(a[9]), .ZN(n874) );
  NAND3_X2 U1432 ( .A1(n875), .A2(n632), .A3(n874), .ZN(n1153) );
  NAND2_X2 U1433 ( .A1(n866), .A2(n1153), .ZN(n881) );
  NAND2_X2 U1434 ( .A1(n689), .A2(a[30]), .ZN(n877) );
  NAND2_X2 U1435 ( .A1(n922), .A2(a[1]), .ZN(n876) );
  NAND3_X2 U1436 ( .A1(n877), .A2(n682), .A3(n876), .ZN(n964) );
  NAND2_X2 U1437 ( .A1(n964), .A2(b[4]), .ZN(n879) );
  NAND2_X2 U1438 ( .A1(n918), .A2(a[17]), .ZN(n878) );
  NAND3_X2 U1439 ( .A1(n573), .A2(n879), .A3(n878), .ZN(n1152) );
  MUX2_X2 U1440 ( .A(n883), .B(n1075), .S(b[2]), .Z(n963) );
  NAND2_X2 U1441 ( .A1(n885), .A2(n884), .ZN(n933) );
  NAND2_X2 U1442 ( .A1(n915), .A2(a[3]), .ZN(n894) );
  NAND2_X2 U1443 ( .A1(n689), .A2(a[19]), .ZN(n887) );
  NAND2_X2 U1444 ( .A1(n922), .A2(a[12]), .ZN(n886) );
  NAND3_X2 U1445 ( .A1(n887), .A2(n924), .A3(n886), .ZN(n1055) );
  NAND2_X2 U1446 ( .A1(n842), .A2(n1055), .ZN(n893) );
  NAND2_X2 U1447 ( .A1(n689), .A2(a[27]), .ZN(n889) );
  NAND2_X2 U1448 ( .A1(n922), .A2(a[4]), .ZN(n888) );
  NAND3_X2 U1449 ( .A1(n889), .A2(n632), .A3(n888), .ZN(n1039) );
  NAND2_X2 U1450 ( .A1(n1039), .A2(b[4]), .ZN(n891) );
  NAND2_X2 U1451 ( .A1(n918), .A2(a[20]), .ZN(n890) );
  NAND3_X2 U1452 ( .A1(n577), .A2(n891), .A3(n890), .ZN(n1054) );
  NAND2_X2 U1453 ( .A1(b[3]), .A2(n1054), .ZN(n892) );
  NAND4_X2 U1454 ( .A1(n895), .A2(n894), .A3(n893), .A4(n892), .ZN(n905) );
  AOI22_X2 U1455 ( .A1(n650), .A2(a[24]), .B1(n915), .B2(a[7]), .ZN(n904) );
  NAND2_X2 U1456 ( .A1(n689), .A2(a[23]), .ZN(n897) );
  NAND2_X2 U1457 ( .A1(n922), .A2(a[8]), .ZN(n896) );
  NAND3_X2 U1458 ( .A1(n897), .A2(n632), .A3(n896), .ZN(n1193) );
  NAND2_X2 U1459 ( .A1(n842), .A2(n1193), .ZN(n903) );
  NAND2_X2 U1460 ( .A1(n689), .A2(a[31]), .ZN(n899) );
  NAND2_X2 U1461 ( .A1(n922), .A2(a[0]), .ZN(n898) );
  NAND3_X2 U1462 ( .A1(n899), .A2(n682), .A3(n898), .ZN(n948) );
  NAND2_X2 U1463 ( .A1(n948), .A2(b[4]), .ZN(n901) );
  NAND2_X2 U1464 ( .A1(n918), .A2(a[16]), .ZN(n900) );
  NAND3_X2 U1465 ( .A1(n580), .A2(n901), .A3(n900), .ZN(n1192) );
  MUX2_X2 U1466 ( .A(n905), .B(n1101), .S(b[2]), .Z(n982) );
  NAND2_X2 U1467 ( .A1(b[1]), .A2(n982), .ZN(n932) );
  NAND2_X2 U1468 ( .A1(n689), .A2(a[25]), .ZN(n907) );
  NAND2_X2 U1469 ( .A1(n922), .A2(a[6]), .ZN(n906) );
  NAND3_X2 U1470 ( .A1(n907), .A2(n924), .A3(n906), .ZN(n1116) );
  NAND2_X2 U1471 ( .A1(n1116), .A2(b[4]), .ZN(n909) );
  NAND2_X2 U1472 ( .A1(n918), .A2(a[22]), .ZN(n908) );
  NAND3_X2 U1473 ( .A1(n582), .A2(n909), .A3(n908), .ZN(n979) );
  NAND2_X2 U1474 ( .A1(b[3]), .A2(n979), .ZN(n913) );
  NAND2_X2 U1475 ( .A1(n689), .A2(a[17]), .ZN(n911) );
  NAND2_X2 U1476 ( .A1(n922), .A2(a[14]), .ZN(n910) );
  NAND4_X2 U1477 ( .A1(n913), .A2(n924), .A3(n661), .A4(n912), .ZN(n914) );
  NAND2_X2 U1478 ( .A1(n1432), .A2(n914), .ZN(n931) );
  NAND2_X2 U1479 ( .A1(n915), .A2(a[5]), .ZN(n928) );
  NAND2_X2 U1480 ( .A1(n689), .A2(a[29]), .ZN(n917) );
  NAND2_X2 U1481 ( .A1(n922), .A2(a[2]), .ZN(n916) );
  NAND3_X2 U1482 ( .A1(n917), .A2(n631), .A3(n916), .ZN(n1010) );
  NAND2_X2 U1483 ( .A1(n1010), .A2(b[4]), .ZN(n920) );
  NAND2_X2 U1484 ( .A1(n918), .A2(a[18]), .ZN(n919) );
  NAND3_X2 U1485 ( .A1(n585), .A2(n920), .A3(n919), .ZN(n1103) );
  NAND2_X2 U1486 ( .A1(b[3]), .A2(n1103), .ZN(n927) );
  NAND2_X2 U1487 ( .A1(n689), .A2(a[21]), .ZN(n925) );
  NAND2_X2 U1488 ( .A1(n922), .A2(a[10]), .ZN(n923) );
  NAND3_X2 U1489 ( .A1(n925), .A2(n632), .A3(n923), .ZN(n1104) );
  NAND2_X2 U1490 ( .A1(n842), .A2(n1104), .ZN(n926) );
  NAND4_X2 U1491 ( .A1(n929), .A2(n928), .A3(n927), .A4(n926), .ZN(n1053) );
  NAND2_X2 U1492 ( .A1(n1430), .A2(n1053), .ZN(n930) );
  NAND3_X2 U1493 ( .A1(n932), .A2(n931), .A3(n930), .ZN(n1731) );
  MUX2_X2 U1494 ( .A(n933), .B(n1731), .S(b[0]), .Z(n934) );
  INV_X4 U1495 ( .A(n934), .ZN(n1848) );
  INV_X4 U1496 ( .A(alu_ctrl[2]), .ZN(n1817) );
  NAND2_X2 U1497 ( .A1(n640), .A2(alu_ctrl[1]), .ZN(n966) );
  INV_X4 U1498 ( .A(n1824), .ZN(n1827) );
  NAND2_X2 U1499 ( .A1(n1827), .A2(n1821), .ZN(n938) );
  INV_X4 U1500 ( .A(n938), .ZN(n943) );
  INV_X4 U1501 ( .A(n1821), .ZN(n935) );
  NAND3_X2 U1502 ( .A1(n1072), .A2(n1001), .A3(n1003), .ZN(n1028) );
  INV_X4 U1503 ( .A(n1028), .ZN(n939) );
  NAND2_X2 U1504 ( .A1(n657), .A2(n939), .ZN(n941) );
  NAND2_X2 U1505 ( .A1(n657), .A2(n1025), .ZN(n940) );
  OAI221_X2 U1506 ( .B1(n943), .B2(n942), .C1(n1027), .C2(n941), .A(n940), 
        .ZN(n944) );
  XNOR2_X2 U1507 ( .A(n944), .B(n1819), .ZN(n1794) );
  XNOR2_X2 U1508 ( .A(a[31]), .B(b[31]), .ZN(n1822) );
  NAND2_X2 U1509 ( .A1(n640), .A2(n949), .ZN(n1847) );
  INV_X4 U1510 ( .A(n1847), .ZN(n954) );
  INV_X4 U1511 ( .A(b[0]), .ZN(n967) );
  INV_X4 U1512 ( .A(n1840), .ZN(n995) );
  INV_X4 U1513 ( .A(n948), .ZN(n1211) );
  NAND2_X2 U1514 ( .A1(n995), .A2(n687), .ZN(n1140) );
  MUX2_X2 U1515 ( .A(n995), .B(n1117), .S(n1432), .Z(n1843) );
  NAND2_X2 U1516 ( .A1(n1732), .A2(alu_ctrl[0]), .ZN(n1711) );
  NAND2_X2 U1517 ( .A1(a[31]), .A2(b[31]), .ZN(n950) );
  NAND2_X2 U1518 ( .A1(n950), .A2(n1840), .ZN(n951) );
  NAND2_X2 U1519 ( .A1(n1732), .A2(n951), .ZN(n952) );
  AOI211_X2 U1520 ( .C1(n1722), .C2(n1843), .A(n955), .B(n665), .ZN(n956) );
  OAI211_X2 U1521 ( .C1(n1848), .C2(n966), .A(n957), .B(n956), .ZN(res[31]) );
  XNOR2_X2 U1522 ( .A(n958), .B(res[31]), .ZN(of) );
  NAND2_X2 U1523 ( .A1(b[30]), .A2(n959), .ZN(n978) );
  MUX2_X2 U1524 ( .A(n698), .B(n1732), .S(b[30]), .Z(n960) );
  INV_X4 U1525 ( .A(n649), .ZN(n965) );
  NAND2_X2 U1526 ( .A1(n961), .A2(n1698), .ZN(n962) );
  NAND2_X2 U1527 ( .A1(n1209), .A2(b[3]), .ZN(n1194) );
  NAND3_X2 U1528 ( .A1(n962), .A2(n670), .A3(n1194), .ZN(n1076) );
  AOI222_X4 U1529 ( .A1(n983), .A2(n1427), .B1(n1076), .B2(n690), .C1(n963), 
        .C2(n981), .ZN(n1727) );
  INV_X4 U1530 ( .A(n964), .ZN(n1222) );
  MUX2_X2 U1531 ( .A(n995), .B(n1141), .S(n1432), .Z(n1744) );
  AOI22_X2 U1532 ( .A1(n965), .A2(n1721), .B1(n1722), .B2(n1744), .ZN(n976) );
  INV_X4 U1533 ( .A(n1731), .ZN(n969) );
  INV_X4 U1534 ( .A(n966), .ZN(n968) );
  INV_X4 U1535 ( .A(n1843), .ZN(n1728) );
  INV_X4 U1536 ( .A(n970), .ZN(n971) );
  XNOR2_X2 U1537 ( .A(n971), .B(n1827), .ZN(n1803) );
  NAND4_X2 U1538 ( .A1(n978), .A2(n977), .A3(n976), .A4(n975), .ZN(res[30]) );
  NAND2_X2 U1539 ( .A1(n979), .A2(n1698), .ZN(n980) );
  NAND3_X2 U1540 ( .A1(n980), .A2(n1194), .A3(n667), .ZN(n1102) );
  NAND2_X2 U1541 ( .A1(n1432), .A2(n983), .ZN(n990) );
  NAND2_X2 U1542 ( .A1(n984), .A2(n1698), .ZN(n986) );
  INV_X4 U1543 ( .A(n985), .ZN(n1295) );
  INV_X4 U1544 ( .A(n1076), .ZN(n1157) );
  INV_X4 U1545 ( .A(n1680), .ZN(n1704) );
  INV_X4 U1546 ( .A(n994), .ZN(n1282) );
  NAND2_X2 U1547 ( .A1(n1432), .A2(n1223), .ZN(n997) );
  NAND2_X2 U1548 ( .A1(n1141), .A2(n1427), .ZN(n996) );
  NAND2_X2 U1549 ( .A1(n995), .A2(b[2]), .ZN(n1011) );
  NAND3_X2 U1550 ( .A1(n997), .A2(n996), .A3(n1011), .ZN(n1703) );
  NAND2_X2 U1551 ( .A1(n1722), .A2(n1703), .ZN(n1016) );
  INV_X4 U1552 ( .A(n998), .ZN(n1002) );
  OAI21_X4 U1553 ( .B1(n1002), .B2(n1050), .A(n1001), .ZN(n1004) );
  XNOR2_X2 U1554 ( .A(n1004), .B(n1003), .ZN(n1805) );
  MUX2_X2 U1555 ( .A(n698), .B(n1732), .S(b[28]), .Z(n1005) );
  NAND2_X2 U1556 ( .A1(n1117), .A2(n1427), .ZN(n1013) );
  INV_X4 U1557 ( .A(n1010), .ZN(n1270) );
  NAND2_X2 U1558 ( .A1(n1432), .A2(n1212), .ZN(n1012) );
  NAND3_X2 U1559 ( .A1(n1013), .A2(n1012), .A3(n1011), .ZN(n1715) );
  NAND3_X2 U1560 ( .A1(n1017), .A2(n1016), .A3(n1015), .ZN(res[28]) );
  MUX2_X2 U1561 ( .A(n696), .B(n1838), .S(b[29]), .Z(n1018) );
  NAND2_X2 U1562 ( .A1(n1018), .A2(n693), .ZN(n1024) );
  INV_X4 U1563 ( .A(n1715), .ZN(n1019) );
  INV_X4 U1564 ( .A(n1020), .ZN(n1021) );
  INV_X4 U1565 ( .A(n1025), .ZN(n1026) );
  OAI21_X4 U1566 ( .B1(n1028), .B2(n1027), .A(n1026), .ZN(n1030) );
  NAND2_X2 U1567 ( .A1(n1031), .A2(n1720), .ZN(n1036) );
  NAND2_X2 U1568 ( .A1(n1844), .A2(n1721), .ZN(n1035) );
  INV_X4 U1569 ( .A(n649), .ZN(n1033) );
  INV_X4 U1570 ( .A(n1714), .ZN(n1032) );
  AOI22_X2 U1571 ( .A1(n1033), .A2(n1032), .B1(n1659), .B2(n1744), .ZN(n1034)
         );
  NAND4_X2 U1572 ( .A1(n1037), .A2(n1036), .A3(n1035), .A4(n1034), .ZN(res[29]) );
  MUX2_X2 U1573 ( .A(n696), .B(n1838), .S(b[27]), .Z(n1038) );
  NAND2_X2 U1574 ( .A1(n1038), .A2(n693), .ZN(n1047) );
  NAND2_X2 U1575 ( .A1(n1212), .A2(n1427), .ZN(n1042) );
  INV_X4 U1576 ( .A(n1039), .ZN(n1310) );
  NAND2_X2 U1577 ( .A1(n1432), .A2(n1271), .ZN(n1041) );
  INV_X4 U1578 ( .A(n1660), .ZN(n1683) );
  INV_X4 U1579 ( .A(n1043), .ZN(n1044) );
  NAND2_X2 U1580 ( .A1(n1844), .A2(n1680), .ZN(n1064) );
  NAND2_X2 U1581 ( .A1(n1052), .A2(n1720), .ZN(n1063) );
  NAND2_X2 U1582 ( .A1(n1432), .A2(n1053), .ZN(n1061) );
  NAND2_X2 U1583 ( .A1(n1101), .A2(n1427), .ZN(n1060) );
  NAND2_X2 U1584 ( .A1(n1054), .A2(n1698), .ZN(n1056) );
  INV_X4 U1585 ( .A(n1055), .ZN(n1308) );
  INV_X4 U1586 ( .A(n1102), .ZN(n1198) );
  AOI22_X2 U1587 ( .A1(n1659), .A2(n1703), .B1(n1719), .B2(n1681), .ZN(n1062)
         );
  NAND4_X2 U1588 ( .A1(n1065), .A2(n1064), .A3(n1063), .A4(n1062), .ZN(res[27]) );
  NAND2_X2 U1589 ( .A1(n658), .A2(n1236), .ZN(n1123) );
  NAND2_X2 U1590 ( .A1(n1184), .A2(n1169), .ZN(n1124) );
  INV_X4 U1591 ( .A(n1068), .ZN(n1069) );
  OAI21_X4 U1592 ( .B1(n1167), .B2(n1070), .A(n1069), .ZN(n1131) );
  XNOR2_X2 U1593 ( .A(n1073), .B(n1072), .ZN(n1776) );
  AOI22_X2 U1594 ( .A1(n1720), .A2(n1074), .B1(n1844), .B2(n1681), .ZN(n1100)
         );
  NAND2_X2 U1595 ( .A1(n1659), .A2(n1660), .ZN(n1099) );
  NAND2_X2 U1596 ( .A1(n1076), .A2(n1427), .ZN(n1083) );
  INV_X4 U1597 ( .A(n1078), .ZN(n1281) );
  NOR2_X4 U1598 ( .A1(n646), .A2(n1079), .ZN(n1300) );
  MUX2_X2 U1599 ( .A(n698), .B(n1732), .S(b[26]), .Z(n1085) );
  NAND2_X2 U1600 ( .A1(n1430), .A2(n1141), .ZN(n1094) );
  INV_X4 U1601 ( .A(n1090), .ZN(n1296) );
  NAND2_X2 U1602 ( .A1(n1432), .A2(n1280), .ZN(n1093) );
  INV_X4 U1603 ( .A(n1657), .ZN(n1095) );
  NAND3_X2 U1604 ( .A1(n1100), .A2(n1099), .A3(n1098), .ZN(res[26]) );
  NAND2_X2 U1605 ( .A1(n1432), .A2(n1101), .ZN(n1110) );
  NAND2_X2 U1606 ( .A1(n1102), .A2(n1427), .ZN(n1109) );
  INV_X4 U1607 ( .A(n1104), .ZN(n1269) );
  NOR2_X4 U1608 ( .A1(n648), .A2(n1105), .ZN(n1314) );
  MUX2_X2 U1609 ( .A(n698), .B(n1732), .S(b[25]), .Z(n1111) );
  INV_X4 U1610 ( .A(n1116), .ZN(n1263) );
  AOI22_X2 U1611 ( .A1(n1432), .A2(n1342), .B1(n1271), .B2(n1427), .ZN(n1119)
         );
  AOI22_X2 U1612 ( .A1(n1430), .A2(n1212), .B1(n1117), .B2(n690), .ZN(n1118)
         );
  NAND2_X2 U1613 ( .A1(n1119), .A2(n1118), .ZN(n1640) );
  INV_X4 U1614 ( .A(n1640), .ZN(n1120) );
  NOR3_X4 U1615 ( .A1(n1181), .A2(n1124), .A3(n1123), .ZN(n1127) );
  INV_X4 U1616 ( .A(n1128), .ZN(n1130) );
  NAND2_X2 U1617 ( .A1(n1130), .A2(n1129), .ZN(n1132) );
  NAND2_X2 U1618 ( .A1(n1659), .A2(n1657), .ZN(n1134) );
  NAND2_X2 U1619 ( .A1(n1137), .A2(n1136), .ZN(res[25]) );
  MUX2_X2 U1620 ( .A(n696), .B(n1838), .S(b[24]), .Z(n1138) );
  NAND2_X2 U1621 ( .A1(n1138), .A2(n693), .ZN(n1151) );
  NAND2_X2 U1622 ( .A1(n1280), .A2(n1427), .ZN(n1145) );
  INV_X4 U1623 ( .A(n1139), .ZN(n1240) );
  NAND2_X2 U1624 ( .A1(n1432), .A2(n1353), .ZN(n1144) );
  NAND2_X2 U1625 ( .A1(n1430), .A2(n1223), .ZN(n1143) );
  NAND2_X2 U1626 ( .A1(n1141), .A2(n690), .ZN(n1142) );
  NAND4_X2 U1627 ( .A1(n1145), .A2(n1144), .A3(n1143), .A4(n1142), .ZN(n1607)
         );
  INV_X4 U1628 ( .A(n1607), .ZN(n1614) );
  INV_X4 U1629 ( .A(n1146), .ZN(n1148) );
  INV_X4 U1630 ( .A(b[24]), .ZN(n1147) );
  INV_X4 U1631 ( .A(n1153), .ZN(n1221) );
  NOR2_X4 U1632 ( .A1(n645), .A2(n1154), .ZN(n1370) );
  NAND2_X2 U1633 ( .A1(n1161), .A2(n1160), .ZN(n1627) );
  NAND2_X2 U1634 ( .A1(n1719), .A2(n1627), .ZN(n1175) );
  NAND2_X2 U1635 ( .A1(n1844), .A2(n1641), .ZN(n1174) );
  INV_X4 U1636 ( .A(n1162), .ZN(n1163) );
  NAND2_X2 U1637 ( .A1(n1232), .A2(n1236), .ZN(n1164) );
  NAND2_X2 U1638 ( .A1(n1164), .A2(n1237), .ZN(n1182) );
  INV_X4 U1639 ( .A(n1165), .ZN(n1185) );
  AOI21_X2 U1640 ( .B1(n1182), .B2(n1184), .A(n1185), .ZN(n1166) );
  OAI21_X4 U1641 ( .B1(n1168), .B2(n1167), .A(n1166), .ZN(n1189) );
  INV_X4 U1642 ( .A(n1170), .ZN(n1171) );
  XNOR2_X2 U1643 ( .A(n1172), .B(n1171), .ZN(n1778) );
  NAND4_X2 U1644 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), .ZN(res[24]) );
  NOR2_X4 U1645 ( .A1(n1179), .A2(n1254), .ZN(n1233) );
  NAND2_X2 U1646 ( .A1(n1259), .A2(n1236), .ZN(n1180) );
  NOR2_X4 U1647 ( .A1(n1181), .A2(n1180), .ZN(n1183) );
  NAND2_X2 U1648 ( .A1(n1185), .A2(n1184), .ZN(n1186) );
  NOR2_X4 U1649 ( .A1(n1187), .A2(n1186), .ZN(n1188) );
  INV_X4 U1650 ( .A(n1188), .ZN(n1190) );
  INV_X4 U1651 ( .A(n1191), .ZN(n1782) );
  INV_X4 U1652 ( .A(n1193), .ZN(n1210) );
  NOR2_X4 U1653 ( .A1(n647), .A2(n1195), .ZN(n1403) );
  NAND2_X2 U1654 ( .A1(n1202), .A2(n1201), .ZN(n1590) );
  MUX2_X2 U1655 ( .A(n698), .B(n1732), .S(b[23]), .Z(n1203) );
  INV_X4 U1656 ( .A(a[23]), .ZN(n1206) );
  AOI221_X2 U1657 ( .B1(n1782), .B2(n1720), .C1(n1719), .C2(n1590), .A(n1208), 
        .ZN(n1219) );
  INV_X4 U1658 ( .A(n1209), .ZN(n1307) );
  OAI221_X2 U1659 ( .B1(n1211), .B2(n1309), .C1(n1210), .C2(n687), .A(n1307), 
        .ZN(n1410) );
  INV_X4 U1660 ( .A(n1410), .ZN(n1215) );
  NAND2_X2 U1661 ( .A1(n1342), .A2(n1427), .ZN(n1214) );
  AOI22_X2 U1662 ( .A1(n1430), .A2(n1271), .B1(n1212), .B2(n690), .ZN(n1213)
         );
  OAI211_X2 U1663 ( .C1(n1215), .C2(n1406), .A(n1214), .B(n1213), .ZN(n1247)
         );
  INV_X4 U1664 ( .A(n1247), .ZN(n1609) );
  NAND2_X2 U1665 ( .A1(n1659), .A2(n1607), .ZN(n1216) );
  OAI21_X2 U1666 ( .B1(n1609), .B2(n636), .A(n1216), .ZN(n1217) );
  AOI21_X2 U1667 ( .B1(n1844), .B2(n1627), .A(n1217), .ZN(n1218) );
  NAND2_X2 U1668 ( .A1(n1219), .A2(n1218), .ZN(res[23]) );
  MUX2_X2 U1669 ( .A(n696), .B(n1838), .S(b[22]), .Z(n1220) );
  NAND2_X2 U1670 ( .A1(n1220), .A2(n693), .ZN(n1231) );
  OAI221_X2 U1671 ( .B1(n1222), .B2(n1309), .C1(n1221), .C2(n687), .A(n1307), 
        .ZN(n1433) );
  INV_X4 U1672 ( .A(n1433), .ZN(n1226) );
  NAND2_X2 U1673 ( .A1(n1353), .A2(n1427), .ZN(n1225) );
  AOI22_X2 U1674 ( .A1(n1430), .A2(n1280), .B1(n1223), .B2(n690), .ZN(n1224)
         );
  OAI211_X2 U1675 ( .C1(n1226), .C2(n1406), .A(n1225), .B(n1224), .ZN(n1558)
         );
  INV_X4 U1676 ( .A(n1558), .ZN(n1569) );
  INV_X4 U1677 ( .A(n1227), .ZN(n1228) );
  INV_X4 U1678 ( .A(n1232), .ZN(n1235) );
  NAND3_X4 U1679 ( .A1(n1256), .A2(n1259), .A3(n1233), .ZN(n1234) );
  XNOR2_X2 U1680 ( .A(n1238), .B(n1237), .ZN(n1775) );
  NAND2_X2 U1681 ( .A1(n1720), .A2(n1239), .ZN(n1250) );
  OAI221_X2 U1682 ( .B1(n1240), .B2(n1309), .C1(n641), .C2(n687), .A(n1307), 
        .ZN(n1431) );
  INV_X4 U1683 ( .A(n1431), .ZN(n1371) );
  NAND2_X2 U1684 ( .A1(n1246), .A2(n1245), .ZN(n1587) );
  NAND2_X2 U1685 ( .A1(n1719), .A2(n1587), .ZN(n1249) );
  AOI22_X2 U1686 ( .A1(n1716), .A2(n1247), .B1(n1844), .B2(n1590), .ZN(n1248)
         );
  NAND4_X2 U1687 ( .A1(n1251), .A2(n1250), .A3(n1249), .A4(n1248), .ZN(res[22]) );
  NAND2_X2 U1688 ( .A1(b[21]), .A2(n1252), .ZN(n1278) );
  MUX2_X2 U1689 ( .A(n698), .B(n1732), .S(b[21]), .Z(n1253) );
  OAI211_X2 U1690 ( .C1(n1260), .C2(n1293), .A(n1259), .B(n1258), .ZN(n1262)
         );
  OAI22_X2 U1691 ( .A1(n639), .A2(n1406), .B1(n246), .B2(n1314), .ZN(n1266) );
  OAI221_X2 U1692 ( .B1(n1263), .B2(n1309), .C1(n644), .C2(n687), .A(n1307), 
        .ZN(n1400) );
  INV_X4 U1693 ( .A(n1400), .ZN(n1407) );
  NAND2_X2 U1694 ( .A1(n1410), .A2(n1427), .ZN(n1274) );
  OAI221_X2 U1695 ( .B1(n1270), .B2(n1309), .C1(n1269), .C2(n687), .A(n1307), 
        .ZN(n1411) );
  NAND2_X2 U1696 ( .A1(n1432), .A2(n1411), .ZN(n1273) );
  AOI22_X2 U1697 ( .A1(n1430), .A2(n1342), .B1(n1271), .B2(n690), .ZN(n1272)
         );
  NAND4_X2 U1698 ( .A1(n1278), .A2(n1277), .A3(n1276), .A4(n1275), .ZN(res[21]) );
  MUX2_X2 U1699 ( .A(n696), .B(n1838), .S(b[20]), .Z(n1279) );
  NAND2_X2 U1700 ( .A1(n1279), .A2(n693), .ZN(n1292) );
  NAND2_X2 U1701 ( .A1(n1430), .A2(n1353), .ZN(n1286) );
  NAND2_X2 U1702 ( .A1(n1280), .A2(n690), .ZN(n1285) );
  OAI221_X2 U1703 ( .B1(n1282), .B2(n1309), .C1(n1281), .C2(n687), .A(n1307), 
        .ZN(n1429) );
  NAND2_X2 U1704 ( .A1(n1432), .A2(n1429), .ZN(n1284) );
  NAND2_X2 U1705 ( .A1(n1433), .A2(n1427), .ZN(n1283) );
  NAND4_X2 U1706 ( .A1(n1286), .A2(n1285), .A3(n1284), .A4(n1283), .ZN(n1536)
         );
  INV_X4 U1707 ( .A(n1536), .ZN(n1315) );
  INV_X4 U1708 ( .A(n1287), .ZN(n1289) );
  INV_X4 U1709 ( .A(b[20]), .ZN(n1288) );
  XNOR2_X2 U1710 ( .A(n1294), .B(n1293), .ZN(n1781) );
  NAND2_X2 U1711 ( .A1(n1720), .A2(n1781), .ZN(n1305) );
  OAI221_X2 U1712 ( .B1(n1296), .B2(n1309), .C1(n1295), .C2(n687), .A(n1307), 
        .ZN(n1428) );
  INV_X4 U1713 ( .A(n1428), .ZN(n1366) );
  OAI221_X2 U1714 ( .B1(n246), .B2(n1370), .C1(n1300), .C2(n1406), .A(n1299), 
        .ZN(n1544) );
  INV_X4 U1715 ( .A(n1559), .ZN(n1545) );
  NAND4_X2 U1716 ( .A1(n1306), .A2(n1305), .A3(n1304), .A4(n1303), .ZN(res[20]) );
  OAI221_X2 U1717 ( .B1(n1310), .B2(n1309), .C1(n1308), .C2(n687), .A(n1307), 
        .ZN(n1401) );
  INV_X4 U1718 ( .A(n1401), .ZN(n1405) );
  OAI221_X2 U1719 ( .B1(n246), .B2(n1403), .C1(n1314), .C2(n1406), .A(n1313), 
        .ZN(n1521) );
  AOI21_X2 U1720 ( .B1(n1719), .B2(n1521), .A(n1316), .ZN(n1351) );
  INV_X4 U1721 ( .A(n1459), .ZN(n1390) );
  INV_X4 U1722 ( .A(n1318), .ZN(n1321) );
  INV_X4 U1723 ( .A(n1333), .ZN(n1324) );
  NAND2_X2 U1724 ( .A1(n652), .A2(n1376), .ZN(n1332) );
  INV_X4 U1725 ( .A(n1332), .ZN(n1323) );
  NAND3_X2 U1726 ( .A1(n1324), .A2(n1335), .A3(n1323), .ZN(n1325) );
  NAND2_X2 U1727 ( .A1(n1326), .A2(n1325), .ZN(n1784) );
  INV_X4 U1728 ( .A(n1784), .ZN(n1327) );
  INV_X4 U1729 ( .A(n1380), .ZN(n1330) );
  OAI211_X2 U1730 ( .C1(n1333), .C2(n1332), .A(n1378), .B(n1331), .ZN(n1336)
         );
  NAND3_X2 U1731 ( .A1(n1336), .A2(n1335), .A3(n1334), .ZN(n1347) );
  MUX2_X2 U1732 ( .A(n698), .B(n1732), .S(b[19]), .Z(n1337) );
  AOI22_X2 U1733 ( .A1(n1432), .A2(n1401), .B1(n1411), .B2(n1427), .ZN(n1344)
         );
  AOI22_X2 U1734 ( .A1(n1430), .A2(n1410), .B1(n1342), .B2(n690), .ZN(n1343)
         );
  NAND2_X2 U1735 ( .A1(n1344), .A2(n1343), .ZN(n1500) );
  INV_X4 U1736 ( .A(n1500), .ZN(n1514) );
  NAND3_X2 U1737 ( .A1(n1351), .A2(n1350), .A3(n1349), .ZN(res[19]) );
  MUX2_X2 U1738 ( .A(n697), .B(n1838), .S(b[18]), .Z(n1352) );
  NAND2_X2 U1739 ( .A1(n1352), .A2(n693), .ZN(n1363) );
  NAND2_X2 U1740 ( .A1(n1430), .A2(n1433), .ZN(n1355) );
  NAND2_X2 U1741 ( .A1(n1353), .A2(n690), .ZN(n1354) );
  NAND2_X2 U1742 ( .A1(n1355), .A2(n1354), .ZN(n1357) );
  INV_X4 U1743 ( .A(n1429), .ZN(n1364) );
  OAI22_X2 U1744 ( .A1(n1366), .A2(n1406), .B1(n246), .B2(n1364), .ZN(n1356)
         );
  INV_X4 U1745 ( .A(n1358), .ZN(n1360) );
  INV_X4 U1746 ( .A(b[18]), .ZN(n1359) );
  OAI221_X2 U1747 ( .B1(n246), .B2(n1371), .C1(n1370), .C2(n1406), .A(n1369), 
        .ZN(n1509) );
  NAND2_X2 U1748 ( .A1(n1719), .A2(n1509), .ZN(n1383) );
  NAND2_X2 U1749 ( .A1(n1844), .A2(n1521), .ZN(n1382) );
  NAND2_X2 U1750 ( .A1(n1373), .A2(n1372), .ZN(n1374) );
  INV_X4 U1751 ( .A(n1374), .ZN(n1396) );
  INV_X4 U1752 ( .A(n1426), .ZN(n1377) );
  NAND4_X2 U1753 ( .A1(n1384), .A2(n1383), .A3(n1382), .A4(n1381), .ZN(res[18]) );
  INV_X4 U1754 ( .A(n1385), .ZN(n1578) );
  NAND2_X2 U1755 ( .A1(n679), .A2(n1448), .ZN(n1495) );
  INV_X4 U1756 ( .A(n1495), .ZN(n1393) );
  NAND3_X2 U1757 ( .A1(n1499), .A2(n1389), .A3(n1454), .ZN(n1391) );
  NAND3_X2 U1758 ( .A1(n1393), .A2(n655), .A3(n1392), .ZN(n1394) );
  INV_X4 U1759 ( .A(n1397), .ZN(n1399) );
  OAI22_X2 U1760 ( .A1(n736), .A2(n1399), .B1(n1398), .B2(n1397), .ZN(n1787)
         );
  INV_X4 U1761 ( .A(n1411), .ZN(n1404) );
  AOI22_X2 U1762 ( .A1(n1430), .A2(n1401), .B1(n1400), .B2(n1427), .ZN(n1402)
         );
  AOI22_X2 U1763 ( .A1(n1430), .A2(n1411), .B1(n1410), .B2(n690), .ZN(n1412)
         );
  NAND2_X2 U1764 ( .A1(n1413), .A2(n1412), .ZN(n1489) );
  INV_X4 U1765 ( .A(n1489), .ZN(n1424) );
  MUX2_X2 U1766 ( .A(n698), .B(n1732), .S(b[17]), .Z(n1415) );
  INV_X4 U1767 ( .A(a[17]), .ZN(n1418) );
  AOI211_X2 U1768 ( .C1(n1844), .C2(n1509), .A(n1421), .B(n1420), .ZN(n1422)
         );
  OAI211_X2 U1769 ( .C1(n633), .C2(n1787), .A(n1423), .B(n1422), .ZN(res[17])
         );
  NAND2_X2 U1770 ( .A1(n1720), .A2(n1750), .ZN(n1446) );
  NAND2_X2 U1771 ( .A1(n636), .A2(n649), .ZN(n1444) );
  NAND2_X2 U1772 ( .A1(n1428), .A2(n1427), .ZN(n1437) );
  NAND2_X2 U1773 ( .A1(n1430), .A2(n1429), .ZN(n1436) );
  NAND2_X2 U1774 ( .A1(n1432), .A2(n1431), .ZN(n1435) );
  NAND2_X2 U1775 ( .A1(n1433), .A2(n690), .ZN(n1434) );
  NAND4_X2 U1776 ( .A1(n1437), .A2(n1436), .A3(n1435), .A4(n1434), .ZN(n1467)
         );
  MUX2_X2 U1777 ( .A(n697), .B(n1838), .S(b[16]), .Z(n1438) );
  AOI21_X2 U1778 ( .B1(n1438), .B2(n693), .A(n1439), .ZN(n1443) );
  NAND2_X2 U1779 ( .A1(n698), .A2(n1439), .ZN(n1441) );
  AOI21_X2 U1780 ( .B1(n1441), .B2(n693), .A(n1440), .ZN(n1442) );
  NAND3_X2 U1781 ( .A1(n1447), .A2(n1446), .A3(n1445), .ZN(res[16]) );
  NAND2_X2 U1782 ( .A1(n1722), .A2(n1488), .ZN(n1472) );
  NAND2_X2 U1783 ( .A1(n1719), .A2(n1489), .ZN(n1471) );
  INV_X4 U1784 ( .A(n1449), .ZN(n1451) );
  NAND2_X2 U1785 ( .A1(n1451), .A2(n1450), .ZN(n1456) );
  NAND2_X2 U1786 ( .A1(n1458), .A2(n1459), .ZN(n1457) );
  INV_X4 U1787 ( .A(n1752), .ZN(n1460) );
  NAND2_X2 U1788 ( .A1(n1460), .A2(n1720), .ZN(n1470) );
  NAND2_X2 U1789 ( .A1(n637), .A2(n634), .ZN(n1468) );
  MUX2_X2 U1790 ( .A(n697), .B(n1838), .S(b[15]), .Z(n1461) );
  INV_X4 U1791 ( .A(a[15]), .ZN(n1462) );
  AOI21_X2 U1792 ( .B1(n1461), .B2(n693), .A(n1462), .ZN(n1466) );
  NAND2_X2 U1793 ( .A1(n698), .A2(n1462), .ZN(n1464) );
  AOI21_X2 U1794 ( .B1(n1464), .B2(n693), .A(n1463), .ZN(n1465) );
  NAND4_X2 U1795 ( .A1(n1472), .A2(n1471), .A3(n1470), .A4(n1469), .ZN(res[15]) );
  MUX2_X2 U1796 ( .A(n697), .B(n1838), .S(b[14]), .Z(n1473) );
  NAND2_X2 U1797 ( .A1(n1473), .A2(n693), .ZN(n1479) );
  INV_X4 U1798 ( .A(n1474), .ZN(n1476) );
  INV_X4 U1799 ( .A(b[14]), .ZN(n1475) );
  NAND2_X2 U1800 ( .A1(n1722), .A2(n1509), .ZN(n1492) );
  XNOR2_X2 U1801 ( .A(n1486), .B(n1485), .ZN(n1768) );
  NAND2_X2 U1802 ( .A1(n1720), .A2(n1487), .ZN(n1491) );
  AOI22_X2 U1803 ( .A1(n1844), .A2(n1489), .B1(n1659), .B2(n1488), .ZN(n1490)
         );
  NAND4_X2 U1804 ( .A1(n1493), .A2(n1492), .A3(n1491), .A4(n1490), .ZN(res[14]) );
  INV_X4 U1805 ( .A(n1498), .ZN(n1497) );
  AOI22_X2 U1806 ( .A1(n672), .A2(n1720), .B1(n1719), .B2(n1500), .ZN(n1512)
         );
  NAND2_X2 U1807 ( .A1(n1722), .A2(n1521), .ZN(n1511) );
  MUX2_X2 U1808 ( .A(n698), .B(n1732), .S(b[13]), .Z(n1501) );
  AOI211_X2 U1809 ( .C1(n1659), .C2(n1509), .A(n1508), .B(n1507), .ZN(n1510)
         );
  NAND3_X2 U1810 ( .A1(n1512), .A2(n1511), .A3(n1510), .ZN(res[13]) );
  MUX2_X2 U1811 ( .A(n697), .B(n1838), .S(b[12]), .Z(n1513) );
  NAND2_X2 U1812 ( .A1(n1513), .A2(n693), .ZN(n1520) );
  INV_X4 U1813 ( .A(n1515), .ZN(n1517) );
  INV_X4 U1814 ( .A(b[12]), .ZN(n1516) );
  NAND2_X2 U1815 ( .A1(n1659), .A2(n1521), .ZN(n1532) );
  INV_X4 U1816 ( .A(n1525), .ZN(n1538) );
  NAND2_X2 U1817 ( .A1(n1583), .A2(n1523), .ZN(n1557) );
  NAND2_X2 U1818 ( .A1(n1525), .A2(n1556), .ZN(n1526) );
  OAI211_X2 U1819 ( .C1(n1538), .C2(n1557), .A(n1539), .B(n1526), .ZN(n1542)
         );
  NAND2_X2 U1820 ( .A1(n1542), .A2(n1527), .ZN(n1529) );
  XNOR2_X2 U1821 ( .A(n1529), .B(n1528), .ZN(n1774) );
  AOI22_X2 U1822 ( .A1(n965), .A2(n1536), .B1(n1720), .B2(n1774), .ZN(n1530)
         );
  NAND4_X2 U1823 ( .A1(n1533), .A2(n1532), .A3(n1531), .A4(n1530), .ZN(res[12]) );
  NAND2_X2 U1824 ( .A1(b[11]), .A2(n1534), .ZN(n1552) );
  MUX2_X2 U1825 ( .A(n698), .B(n1732), .S(b[11]), .Z(n1535) );
  INV_X4 U1826 ( .A(n1555), .ZN(n1537) );
  AOI22_X2 U1827 ( .A1(n1722), .A2(n1537), .B1(n1844), .B2(n1536), .ZN(n1550)
         );
  INV_X4 U1828 ( .A(n1557), .ZN(n1541) );
  NAND2_X2 U1829 ( .A1(n1543), .A2(n1542), .ZN(n1783) );
  INV_X4 U1830 ( .A(n1544), .ZN(n1546) );
  OAI22_X2 U1831 ( .A1(n1546), .A2(n637), .B1(n1545), .B2(n649), .ZN(n1547) );
  NAND4_X2 U1832 ( .A1(n1552), .A2(n1551), .A3(n1550), .A4(n1549), .ZN(res[11]) );
  NAND2_X2 U1833 ( .A1(b[10]), .A2(n1553), .ZN(n1563) );
  MUX2_X2 U1834 ( .A(n698), .B(n1732), .S(b[10]), .Z(n1554) );
  XNOR2_X2 U1835 ( .A(n1557), .B(n1556), .ZN(n1766) );
  AOI22_X2 U1836 ( .A1(n1716), .A2(n1537), .B1(n1720), .B2(n1766), .ZN(n1561)
         );
  NAND4_X2 U1837 ( .A1(n1563), .A2(n1562), .A3(n1561), .A4(n1560), .ZN(res[10]) );
  MUX2_X2 U1838 ( .A(n698), .B(n1732), .S(b[9]), .Z(n1564) );
  AOI211_X2 U1839 ( .C1(n1722), .C2(n1590), .A(n1571), .B(n1570), .ZN(n1589)
         );
  INV_X4 U1840 ( .A(n1572), .ZN(n1576) );
  NAND3_X2 U1841 ( .A1(n1582), .A2(n1581), .A3(n1580), .ZN(n1584) );
  NAND2_X2 U1842 ( .A1(n1584), .A2(n1583), .ZN(n1754) );
  AOI211_X2 U1843 ( .C1(n1659), .C2(n1587), .A(n1586), .B(n1585), .ZN(n1588)
         );
  NAND2_X2 U1844 ( .A1(n1589), .A2(n1588), .ZN(res[9]) );
  INV_X4 U1845 ( .A(n1590), .ZN(n1599) );
  INV_X4 U1846 ( .A(n1639), .ZN(n1594) );
  NAND2_X2 U1847 ( .A1(n1595), .A2(n1621), .ZN(n1624) );
  NAND2_X2 U1848 ( .A1(n1624), .A2(n1596), .ZN(n1598) );
  OAI22_X2 U1849 ( .A1(n1599), .A2(n637), .B1(n1749), .B2(n633), .ZN(n1606) );
  MUX2_X2 U1850 ( .A(n1732), .B(n698), .S(n109), .Z(n1600) );
  NOR2_X2 U1851 ( .A1(n1606), .A2(n1605), .ZN(n1612) );
  NAND2_X2 U1852 ( .A1(n1719), .A2(n1607), .ZN(n1608) );
  OAI21_X2 U1853 ( .B1(n1609), .B2(n634), .A(n1608), .ZN(n1610) );
  AOI21_X2 U1854 ( .B1(n1722), .B2(n1627), .A(n1610), .ZN(n1611) );
  NAND2_X2 U1855 ( .A1(n1612), .A2(n1611), .ZN(res[8]) );
  MUX2_X2 U1856 ( .A(n696), .B(n1838), .S(b[7]), .Z(n1613) );
  NAND2_X2 U1857 ( .A1(n1613), .A2(n693), .ZN(n1620) );
  INV_X4 U1858 ( .A(n1615), .ZN(n1617) );
  INV_X4 U1859 ( .A(b[7]), .ZN(n1616) );
  INV_X4 U1860 ( .A(n1621), .ZN(n1623) );
  NAND2_X2 U1861 ( .A1(n1623), .A2(n1622), .ZN(n1625) );
  NAND2_X2 U1862 ( .A1(n1625), .A2(n1624), .ZN(n1769) );
  INV_X4 U1863 ( .A(n1769), .ZN(n1626) );
  NAND2_X2 U1864 ( .A1(n1626), .A2(n1720), .ZN(n1630) );
  NAND2_X2 U1865 ( .A1(n1722), .A2(n1641), .ZN(n1629) );
  AOI22_X2 U1866 ( .A1(n965), .A2(n1640), .B1(n1659), .B2(n1627), .ZN(n1628)
         );
  NAND4_X2 U1867 ( .A1(n1631), .A2(n1630), .A3(n1629), .A4(n1628), .ZN(res[7])
         );
  MUX2_X2 U1868 ( .A(n1838), .B(n697), .S(n111), .Z(n1633) );
  INV_X4 U1869 ( .A(a[6]), .ZN(n1632) );
  INV_X4 U1870 ( .A(n1634), .ZN(n1635) );
  AOI22_X2 U1871 ( .A1(n1765), .A2(n1720), .B1(n1844), .B2(n1640), .ZN(n1644)
         );
  NAND2_X2 U1872 ( .A1(n1722), .A2(n1658), .ZN(n1643) );
  AOI22_X2 U1873 ( .A1(n1033), .A2(n1657), .B1(n1659), .B2(n1641), .ZN(n1642)
         );
  NAND4_X2 U1874 ( .A1(n1645), .A2(n1644), .A3(n1643), .A4(n1642), .ZN(res[6])
         );
  NAND2_X2 U1875 ( .A1(n1648), .A2(n1647), .ZN(n1650) );
  NAND2_X2 U1876 ( .A1(n1650), .A2(n1649), .ZN(n1762) );
  NAND2_X2 U1877 ( .A1(n1732), .A2(a[5]), .ZN(n1651) );
  NAND2_X2 U1878 ( .A1(n1844), .A2(n1657), .ZN(n1663) );
  NAND2_X2 U1879 ( .A1(n1722), .A2(n1681), .ZN(n1662) );
  AOI22_X2 U1880 ( .A1(n1033), .A2(n1660), .B1(n1659), .B2(n1658), .ZN(n1661)
         );
  NAND4_X2 U1881 ( .A1(n1664), .A2(n1663), .A3(n1662), .A4(n1661), .ZN(res[5])
         );
  MUX2_X2 U1882 ( .A(n1838), .B(n697), .S(n115), .Z(n1665) );
  NAND2_X2 U1883 ( .A1(n1665), .A2(n693), .ZN(n1679) );
  INV_X4 U1884 ( .A(n1666), .ZN(n1667) );
  INV_X4 U1885 ( .A(n1672), .ZN(n1673) );
  XNOR2_X2 U1886 ( .A(n1674), .B(n1673), .ZN(n1755) );
  INV_X4 U1887 ( .A(n1675), .ZN(n1676) );
  NAND2_X2 U1888 ( .A1(n1722), .A2(n1680), .ZN(n1688) );
  INV_X4 U1889 ( .A(n1681), .ZN(n1682) );
  INV_X4 U1890 ( .A(n1703), .ZN(n1684) );
  OAI22_X2 U1891 ( .A1(n1684), .A2(n649), .B1(n1683), .B2(n634), .ZN(n1685) );
  MUX2_X2 U1892 ( .A(n696), .B(n1838), .S(b[3]), .Z(n1690) );
  NAND2_X2 U1893 ( .A1(n1690), .A2(n693), .ZN(n1702) );
  INV_X4 U1894 ( .A(n1718), .ZN(n1694) );
  INV_X4 U1895 ( .A(n1697), .ZN(n1699) );
  INV_X4 U1896 ( .A(b[3]), .ZN(n1698) );
  NAND2_X2 U1897 ( .A1(n1719), .A2(n1715), .ZN(n1709) );
  NAND2_X2 U1898 ( .A1(n1844), .A2(n1703), .ZN(n1708) );
  NAND4_X2 U1899 ( .A1(n1710), .A2(n1709), .A3(n1708), .A4(n1707), .ZN(res[3])
         );
  NAND2_X2 U1900 ( .A1(b[2]), .A2(n1712), .ZN(n1726) );
  MUX2_X2 U1901 ( .A(n698), .B(n1732), .S(b[2]), .Z(n1713) );
  INV_X4 U1902 ( .A(n637), .ZN(n1716) );
  AOI22_X2 U1903 ( .A1(n1716), .A2(n1032), .B1(n1844), .B2(n1715), .ZN(n1724)
         );
  INV_X4 U1904 ( .A(n636), .ZN(n1722) );
  XNOR2_X2 U1905 ( .A(n1718), .B(n1717), .ZN(n1759) );
  AOI222_X4 U1906 ( .A1(n1722), .A2(n1721), .B1(n1720), .B2(n1759), .C1(n1719), 
        .C2(n1744), .ZN(n1723) );
  NAND4_X2 U1907 ( .A1(n1726), .A2(n1725), .A3(n1724), .A4(n1723), .ZN(res[2])
         );
  NAND2_X2 U1908 ( .A1(n1722), .A2(n1731), .ZN(n1746) );
  MUX2_X2 U1909 ( .A(n698), .B(n1732), .S(b[1]), .Z(n1733) );
  INV_X4 U1910 ( .A(a[1]), .ZN(n1737) );
  AOI211_X2 U1911 ( .C1(n1844), .C2(n1744), .A(n1743), .B(n1742), .ZN(n1745)
         );
  NAND3_X2 U1912 ( .A1(n1747), .A2(n1746), .A3(n1745), .ZN(res[1]) );
  NAND2_X2 U1913 ( .A1(n1749), .A2(n1748), .ZN(n1773) );
  INV_X4 U1914 ( .A(n1750), .ZN(n1751) );
  INV_X4 U1915 ( .A(n1754), .ZN(n1764) );
  INV_X4 U1916 ( .A(n1755), .ZN(n1760) );
  NAND2_X2 U1917 ( .A1(n642), .A2(n656), .ZN(n1758) );
  NAND3_X2 U1918 ( .A1(n654), .A2(n1762), .A3(n1761), .ZN(n1763) );
  INV_X4 U1919 ( .A(n1766), .ZN(n1767) );
  NAND4_X2 U1920 ( .A1(n1770), .A2(n1769), .A3(n1768), .A4(n1767), .ZN(n1771)
         );
  NAND2_X2 U1921 ( .A1(n1776), .A2(n1775), .ZN(n1780) );
  INV_X4 U1922 ( .A(n1777), .ZN(n1779) );
  NOR3_X4 U1923 ( .A1(n1780), .A2(n1779), .A3(n1778), .ZN(n1792) );
  NOR2_X4 U1924 ( .A1(n1782), .A2(n1781), .ZN(n1788) );
  INV_X4 U1925 ( .A(n1783), .ZN(n1785) );
  NOR2_X4 U1926 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  NAND3_X2 U1927 ( .A1(n1788), .A2(n1787), .A3(n1786), .ZN(n1789) );
  NAND3_X4 U1928 ( .A1(n1793), .A2(n1792), .A3(n1791), .ZN(n1807) );
  INV_X4 U1929 ( .A(n1822), .ZN(n1798) );
  NAND2_X2 U1930 ( .A1(b[31]), .A2(n1798), .ZN(n1812) );
  INV_X4 U1931 ( .A(n1812), .ZN(n1820) );
  AOI21_X4 U1932 ( .B1(n1802), .B2(n1801), .A(n1800), .ZN(n1816) );
  INV_X4 U1933 ( .A(n1803), .ZN(n1804) );
  NOR3_X4 U1934 ( .A1(n1804), .A2(n1806), .A3(n1805), .ZN(n1810) );
  NAND3_X4 U1935 ( .A1(n1810), .A2(n1809), .A3(n1808), .ZN(n1814) );
  MUX2_X2 U1936 ( .A(n1816), .B(n1815), .S(inverse_set), .Z(n1818) );
  INV_X4 U1937 ( .A(inverse_set), .ZN(n1829) );
  NAND2_X2 U1938 ( .A1(n1822), .A2(n1821), .ZN(n1823) );
  OAI21_X4 U1939 ( .B1(n1827), .B2(n1826), .A(n1825), .ZN(n1828) );
  FA_X1 U1940 ( .A(n1830), .B(n1829), .CI(n1828), .S(n1831) );
  MUX2_X2 U1941 ( .A(n1832), .B(n1831), .S(alu_ctrl[2]), .Z(n1833) );
  MUX2_X2 U1942 ( .A(n1835), .B(n1834), .S(alu_ctrl[1]), .Z(n1836) );
  NAND2_X2 U1943 ( .A1(alu_ctrl[3]), .A2(n1836), .ZN(n1880) );
  INV_X4 U1944 ( .A(n1880), .ZN(n1877) );
  NAND2_X2 U1945 ( .A1(a[0]), .A2(b[0]), .ZN(n1837) );
  AOI211_X2 U1946 ( .C1(n1844), .C2(n1843), .A(n1842), .B(n1841), .ZN(n1845)
         );
  OAI211_X2 U1947 ( .C1(n1848), .C2(n1847), .A(n1846), .B(n1845), .ZN(n1878)
         );
  INV_X4 U1948 ( .A(res[28]), .ZN(n1874) );
  NOR2_X4 U1949 ( .A1(res[2]), .A2(res[3]), .ZN(n1860) );
  INV_X4 U1950 ( .A(res[1]), .ZN(n1859) );
  NOR4_X2 U1951 ( .A1(res[4]), .A2(res[5]), .A3(res[6]), .A4(res[7]), .ZN(
        n1858) );
  INV_X4 U1952 ( .A(res[10]), .ZN(n1851) );
  INV_X4 U1953 ( .A(res[9]), .ZN(n1850) );
  INV_X4 U1954 ( .A(res[8]), .ZN(n1849) );
  INV_X4 U1955 ( .A(res[12]), .ZN(n1854) );
  INV_X4 U1956 ( .A(res[11]), .ZN(n1853) );
  NOR2_X4 U1957 ( .A1(res[13]), .A2(res[14]), .ZN(n1852) );
  NAND3_X2 U1958 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1855) );
  NOR2_X2 U1959 ( .A1(n1856), .A2(n1855), .ZN(n1857) );
  NAND4_X2 U1960 ( .A1(n1860), .A2(n1859), .A3(n1858), .A4(n1857), .ZN(n1871)
         );
  INV_X4 U1961 ( .A(res[19]), .ZN(n1864) );
  INV_X4 U1962 ( .A(res[18]), .ZN(n1863) );
  NAND4_X2 U1963 ( .A1(n1864), .A2(n1863), .A3(n1862), .A4(n1861), .ZN(n1870)
         );
  INV_X4 U1964 ( .A(res[29]), .ZN(n1868) );
  INV_X4 U1965 ( .A(res[27]), .ZN(n1867) );
  NAND4_X2 U1966 ( .A1(n1868), .A2(n1867), .A3(n1866), .A4(n1865), .ZN(n1869)
         );
  INV_X4 U1967 ( .A(res[31]), .ZN(n1872) );
  NAND4_X2 U1968 ( .A1(n1875), .A2(n1874), .A3(n1873), .A4(n1872), .ZN(n1876)
         );
  INV_X4 U1969 ( .A(n1878), .ZN(n1879) );
endmodule

