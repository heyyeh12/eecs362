`ifndef _alu_const_vh_
`define _alu_const_vh_

`define alu_sll 4'b0010
`define alu_srl 4'b0000
`define alu_sra 4'b0001
`define alu_add 4'b0100
`define alu_sub 4`b0101
`define alu_and 4'b1000
`define alu_or  4'b1001
`define alu_xor 4'b1010
`define alu_seq 4'b1100
`define alu_sgt 4'b1101
`define alu_sge 4'b1110

`endif // _alu_const_vh_