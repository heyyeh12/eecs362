
module multiplier ( a, b, control, product_in, product_out );
  input [31:0] a;
  input [31:0] b;
  input [1:0] control;
  input [31:0] product_in;
  output [31:0] product_out;
  wire   net86661, net293924, net293927, net293929, net293931, net293933,
         net293935, net293986, net293988, net293989, net293991, net293992,
         net294000, net294004, net294006, net294010, net294012, net294016,
         net294039, net294040, net294043, net294044, net294045, net294048,
         net294051, net294052, net294053, net294054, net294068, net294080,
         net294081, net294082, net294087, net294088, net294092, net294093,
         net294100, net294101, net294102, net294117, net294126, net294137,
         net294153, net294154, net294155, net294156, net294171, net294175,
         net294188, net294194, net294196, net294217, net294220, net294234,
         net294241, net294250, net294251, net294252, net294253, net294285,
         net294298, net294299, net294301, net294303, net294305, net294307,
         net294308, net294309, net294310, net294314, net294320, net294321,
         net294322, net294326, net294329, net294330, net294331, net294332,
         net294333, net294346, net294349, net294353, net294354, net294356,
         net294358, net294359, net294360, net294362, net294364, net294366,
         net294367, net294379, net294388, net294393, net294394, net294425,
         net294426, net294439, net294446, net294448, net294450, net294479,
         net294484, net294485, net294506, net294507, net294510, net294515,
         net294519, net294525, net294526, net294543, net294544, net294573,
         net294574, net294575, net294576, net294577, net294578, net294580,
         net294611, net294628, net294636, net294640, net294642, net294643,
         net294645, net294646, net294649, net294650, net294651, net294652,
         net294656, net294694, net294696, net294698, net294701, net294770,
         net294772, net294779, net294784, net294786, net294787, net294788,
         net294790, net294791, net294792, net294795, net294800, net294801,
         net294808, net294809, net294810, net294815, net294816, net294840,
         net294842, net294843, net294844, net294879, net294881, net294882,
         net294883, net294888, net294889, net294901, net294905, net294907,
         net294908, net294909, net294910, net294911, net294913, net294918,
         net294940, net294980, net294981, net294993, net294994, net294995,
         net295008, net295010, net295012, net295013, net295017, net295020,
         net295156, net295158, net295167, net295168, net295175, net295176,
         net295271, net295273, net295274, net295277, net295278, net295291,
         net295372, net295380, net295387, net295393, net295494, net295495,
         net295496, net295506, net295585, net295587, net295618, net295621,
         net295624, net295626, net295732, net295733, net295734, net295736,
         net295737, net295738, net295748, net295749, net295750, net295754,
         net295755, net295756, net295757, net295759, net295864, net295866,
         net295934, net295978, net295982, net295983, net295989, net295990,
         net295991, net295995, net295996, net296097, net296098, net296099,
         net296104, net296105, net296106, net296216, net296221, net296222,
         net296230, net296324, net296325, net296326, net296333, net296334,
         net296337, net296416, net296417, net296418, net296419, net296424,
         net296430, net296472, net296524, net296529, net296530, net296535,
         net296536, net296544, net296547, net296554, net296672, net296771,
         net296781, net296788, net296808, net296842, net296909, net296910,
         net296911, net296932, net297002, net297009, net297022, net297061,
         net297086, net297128, net297172, net297170, net297168, net297166,
         net297184, net297182, net297180, net297196, net297190, net297188,
         net297210, net297204, net297202, net297222, net297218, net297216,
         net297234, net297230, net297228, net297226, net297250, net297246,
         net297244, net297254, net297268, net297262, net297260, net297276,
         net297274, net297272, net297279, net297278, net297281, net297481,
         net297485, net297515, net297526, net297616, net297615, net297774,
         net297862, net298051, net298149, net298226, net298225, net298392,
         net298389, net298388, net298483, net298482, net298605, net298655,
         net298716, net298730, net298731, net298829, net298857, net298860,
         net298880, net298907, net298909, net298912, net298937, net298969,
         net299021, net299020, net299044, net299047, net299046, net299066,
         net299073, net299089, net299137, net299191, net299241, net299240,
         net299300, net299323, net299325, net299331, net299334, net295379,
         net295377, net295275, net295032, net295031, net295030, net294655,
         net295019, net294334, net294438, net294406, net294653, net295745,
         net295743, net294372, net294371, net294370, net294369, net294042,
         net294657, net298916, net297071, net294219, net294200, net298959,
         net297640, net297100, net294930, net295385, net295288, net294804,
         net294803, net296540, net294931, net294841, net294818, net294817,
         net294532, net294530, net294529, net294405, net297593, net294802,
         net294793, net294680, net294541, net294540, net294539, net294538,
         net294537, net294536, net294535, net294437, net295622, net295509,
         net295508, net295504, net294228, net294218, net294083, net298632,
         net297270, net295165, net295163, net295018, net298968, net295507,
         net295503, net295502, net295500, net295499, net295498, net296539,
         net294407, net294402, net294400, net294249, net299052, net294399,
         net294317, net294313, net294300, net299321, net296553, net296537,
         net296432, net296427, net296426, net296329, net295501, net295382,
         net295289, net296425, net296328, net295752, net295742, net295162,
         net295161, net295160, net295159, net295029, net295028, net294932,
         net294820, net294819, net295287, net295286, net295283, net295282,
         net295281, net295279, net297068, net295280, net295172, net295170,
         net297200, net297198, net294839, net294837, net294806, net294658,
         net293950, net299335, net294205, net297484, net295870, net295869,
         net295868, net295867, net295741, net295739, net295628, net295516,
         net295515, net295514, net295513, net295510, net294447, net294442,
         net294441, net294401, net294248, net294247, net294520, net294509,
         net294396, net294365, net294639, net294531, net294528, net294527,
         net294444, net294440, net297153, net297152, net297070, net294187,
         net297154, net294355, net294347, net294327, net294325, net294324,
         net294199, net294198, net294086, net294085, net294084, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1984, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3270, n3271, n3272, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304;
  wire   [31:0] \set_product_in_sig/z1 ;
  assign \set_product_in_sig/z1  [31] = product_in[31];
  assign \set_product_in_sig/z1  [30] = product_in[30];
  assign \set_product_in_sig/z1  [29] = product_in[29];
  assign \set_product_in_sig/z1  [28] = product_in[28];
  assign \set_product_in_sig/z1  [27] = product_in[27];
  assign \set_product_in_sig/z1  [26] = product_in[26];
  assign \set_product_in_sig/z1  [25] = product_in[25];
  assign \set_product_in_sig/z1  [24] = product_in[24];
  assign \set_product_in_sig/z1  [23] = product_in[23];
  assign \set_product_in_sig/z1  [22] = product_in[22];
  assign \set_product_in_sig/z1  [21] = product_in[21];
  assign \set_product_in_sig/z1  [20] = product_in[20];
  assign \set_product_in_sig/z1  [19] = product_in[19];
  assign \set_product_in_sig/z1  [18] = product_in[18];
  assign \set_product_in_sig/z1  [17] = product_in[17];
  assign \set_product_in_sig/z1  [16] = product_in[16];
  assign \set_product_in_sig/z1  [15] = product_in[15];
  assign \set_product_in_sig/z1  [14] = product_in[14];
  assign \set_product_in_sig/z1  [13] = product_in[13];
  assign \set_product_in_sig/z1  [12] = product_in[12];
  assign \set_product_in_sig/z1  [11] = product_in[11];
  assign \set_product_in_sig/z1  [10] = product_in[10];
  assign \set_product_in_sig/z1  [9] = product_in[9];
  assign \set_product_in_sig/z1  [8] = product_in[8];
  assign \set_product_in_sig/z1  [7] = product_in[7];
  assign \set_product_in_sig/z1  [6] = product_in[6];
  assign \set_product_in_sig/z1  [5] = product_in[5];
  assign \set_product_in_sig/z1  [4] = product_in[4];
  assign \set_product_in_sig/z1  [3] = product_in[3];
  assign \set_product_in_sig/z1  [2] = product_in[2];
  assign \set_product_in_sig/z1  [1] = product_in[1];
  assign \set_product_in_sig/z1  [0] = product_in[0];
  assign product_out[29] = net86661;

  INV_X4 U1134 ( .A(net295271), .ZN(net295273) );
  OAI21_X4 U1135 ( .B1(net295502), .B2(net295503), .A(net295504), .ZN(n1104)
         );
  OAI21_X2 U1136 ( .B1(net295502), .B2(net295503), .A(net295504), .ZN(
        net295500) );
  CLKBUF_X3 U1137 ( .A(n2863), .Z(n1105) );
  INV_X4 U1138 ( .A(n2109), .ZN(n2204) );
  NAND2_X2 U1139 ( .A1(n1977), .A2(n4203), .ZN(n1145) );
  INV_X4 U1141 ( .A(n1876), .ZN(n1219) );
  XOR2_X2 U1144 ( .A(n2311), .B(n2080), .Z(n1106) );
  NAND2_X4 U1145 ( .A1(n2079), .A2(n1109), .ZN(n2080) );
  INV_X1 U1146 ( .A(n1855), .ZN(n1107) );
  INV_X4 U1147 ( .A(n1371), .ZN(n1855) );
  NAND2_X2 U1148 ( .A1(net294396), .A2(n1388), .ZN(n1392) );
  NAND2_X4 U1149 ( .A1(n3168), .A2(n3169), .ZN(n1108) );
  NAND2_X2 U1150 ( .A1(n1496), .A2(n2020), .ZN(n1109) );
  NAND2_X4 U1151 ( .A1(a[3]), .A2(net297230), .ZN(n2020) );
  BUF_X8 U1152 ( .A(net295030), .Z(n1110) );
  OAI21_X4 U1153 ( .B1(net294694), .B2(n3733), .A(net294696), .ZN(n3735) );
  NAND2_X2 U1157 ( .A1(n2881), .A2(n2884), .ZN(n2743) );
  NAND2_X4 U1158 ( .A1(n2915), .A2(n2916), .ZN(n2884) );
  XNOR2_X1 U1160 ( .A(net294841), .B(net294840), .ZN(net294839) );
  INV_X8 U1161 ( .A(n2579), .ZN(n2580) );
  NAND2_X2 U1163 ( .A1(a[13]), .A2(net297485), .ZN(n2588) );
  NAND2_X1 U1164 ( .A1(a[0]), .A2(net297485), .ZN(n3618) );
  INV_X1 U1165 ( .A(net295281), .ZN(net295283) );
  INV_X2 U1167 ( .A(n1630), .ZN(n1372) );
  XNOR2_X1 U1168 ( .A(n2254), .B(n2288), .ZN(n1309) );
  NAND3_X1 U1169 ( .A1(n1514), .A2(n3577), .A3(n1530), .ZN(n1112) );
  INV_X2 U1171 ( .A(n1205), .ZN(n1113) );
  INV_X2 U1172 ( .A(n3403), .ZN(n1205) );
  NAND2_X4 U1173 ( .A1(n3104), .A2(n3105), .ZN(n1120) );
  INV_X4 U1174 ( .A(n3311), .ZN(n1543) );
  XNOR2_X2 U1177 ( .A(n3972), .B(n3971), .ZN(n1114) );
  NAND2_X4 U1178 ( .A1(n4027), .A2(n4026), .ZN(n3971) );
  INV_X8 U1179 ( .A(n4078), .ZN(n4088) );
  NOR2_X2 U1180 ( .A1(n1116), .A2(n3167), .ZN(n1115) );
  INV_X32 U1181 ( .A(n3169), .ZN(n1116) );
  NAND4_X2 U1182 ( .A1(n2767), .A2(n2766), .A3(n2868), .A4(n1312), .ZN(n2768)
         );
  NAND2_X4 U1184 ( .A1(n3083), .A2(n1280), .ZN(n1118) );
  INV_X2 U1185 ( .A(n3396), .ZN(n1119) );
  OAI21_X4 U1186 ( .B1(n2931), .B2(n1347), .A(n3116), .ZN(n3105) );
  INV_X4 U1187 ( .A(net294509), .ZN(net294365) );
  NAND2_X4 U1188 ( .A1(n1494), .A2(n2604), .ZN(n2750) );
  NAND2_X2 U1189 ( .A1(n2604), .A2(n1494), .ZN(n1573) );
  AOI221_X4 U1191 ( .B1(net294051), .B2(n3295), .C1(n1122), .C2(n1129), .A(
        n1123), .ZN(n1121) );
  INV_X4 U1192 ( .A(n1121), .ZN(net294220) );
  XOR2_X2 U1193 ( .A(n3349), .B(n3348), .Z(n1122) );
  AND2_X2 U1194 ( .A1(net294053), .A2(n1618), .ZN(n1123) );
  NAND2_X1 U1195 ( .A1(net297172), .A2(net298226), .ZN(net294126) );
  INV_X8 U1196 ( .A(net294126), .ZN(net294051) );
  NAND2_X1 U1197 ( .A1(n1974), .A2(n2043), .ZN(n3994) );
  INV_X4 U1198 ( .A(net297278), .ZN(n1129) );
  OAI21_X4 U1199 ( .B1(n4032), .B2(n4034), .A(n4031), .ZN(n4075) );
  INV_X2 U1200 ( .A(n3479), .ZN(n1124) );
  INV_X2 U1201 ( .A(n3482), .ZN(n3479) );
  BUF_X4 U1202 ( .A(n4289), .Z(n1683) );
  NAND2_X4 U1203 ( .A1(n3538), .A2(n3536), .ZN(n3607) );
  NOR2_X2 U1204 ( .A1(n1126), .A2(net298731), .ZN(n3674) );
  NAND2_X2 U1205 ( .A1(n1268), .A2(n2066), .ZN(n1168) );
  INV_X1 U1206 ( .A(net294779), .ZN(net294889) );
  OAI21_X1 U1207 ( .B1(n3993), .B2(net297188), .A(n3351), .ZN(n1125) );
  NAND3_X2 U1208 ( .A1(b[24]), .A2(net298226), .A3(n1999), .ZN(n2001) );
  NAND2_X4 U1209 ( .A1(n2482), .A2(n2481), .ZN(n2484) );
  INV_X4 U1210 ( .A(n2199), .ZN(n1561) );
  NOR2_X2 U1211 ( .A1(n3532), .A2(n3604), .ZN(n1126) );
  INV_X2 U1212 ( .A(n3604), .ZN(n3531) );
  NAND2_X4 U1213 ( .A1(a[18]), .A2(net297216), .ZN(n3604) );
  NAND2_X4 U1214 ( .A1(n3229), .A2(n3228), .ZN(n1127) );
  CLKBUF_X2 U1215 ( .A(n1629), .Z(n1160) );
  AOI211_X4 U1216 ( .C1(net295585), .C2(n1129), .A(n1130), .B(n1131), .ZN(
        n1128) );
  AND2_X2 U1217 ( .A1(net294053), .A2(n1421), .ZN(n1130) );
  AND2_X2 U1218 ( .A1(n1420), .A2(net294051), .ZN(n1131) );
  NAND2_X4 U1221 ( .A1(net294448), .A2(n3801), .ZN(n3679) );
  INV_X1 U1222 ( .A(n2282), .ZN(n2189) );
  BUF_X8 U1223 ( .A(n2956), .Z(n1132) );
  NOR2_X2 U1224 ( .A1(net298880), .A2(net294485), .ZN(n3847) );
  NOR3_X2 U1225 ( .A1(n3045), .A2(n2937), .A3(n2936), .ZN(n1133) );
  INV_X8 U1227 ( .A(n1946), .ZN(n1936) );
  INV_X4 U1229 ( .A(n2046), .ZN(n2051) );
  NAND3_X2 U1230 ( .A1(n2079), .A2(n1109), .A3(n2093), .ZN(n2075) );
  INV_X2 U1231 ( .A(net294045), .ZN(net294043) );
  NAND2_X2 U1233 ( .A1(n2475), .A2(n2474), .ZN(n1134) );
  OAI21_X2 U1234 ( .B1(n2283), .B2(n2149), .A(n2282), .ZN(n2147) );
  OAI21_X1 U1236 ( .B1(n3810), .B2(n1173), .A(n3811), .ZN(n3813) );
  NAND2_X2 U1237 ( .A1(n3812), .A2(n3885), .ZN(n3947) );
  NAND2_X1 U1238 ( .A1(n3263), .A2(n3264), .ZN(n1137) );
  INV_X1 U1242 ( .A(n3264), .ZN(n1136) );
  NAND2_X1 U1243 ( .A1(n3770), .A2(n3769), .ZN(n1141) );
  NAND2_X2 U1244 ( .A1(n1139), .A2(n1140), .ZN(n1142) );
  NAND2_X2 U1245 ( .A1(n1141), .A2(n1142), .ZN(n3833) );
  INV_X4 U1246 ( .A(n3770), .ZN(n1139) );
  INV_X2 U1247 ( .A(n3769), .ZN(n1140) );
  INV_X8 U1249 ( .A(n2516), .ZN(n2518) );
  NAND2_X4 U1250 ( .A1(n3970), .A2(n3969), .ZN(n4026) );
  NAND2_X2 U1251 ( .A1(n3670), .A2(n3669), .ZN(n1701) );
  INV_X8 U1252 ( .A(n3048), .ZN(n2947) );
  NAND4_X4 U1253 ( .A1(n3227), .A2(n3374), .A3(n3226), .A4(n1521), .ZN(n3459)
         );
  NAND2_X4 U1254 ( .A1(net294085), .A2(net294086), .ZN(net294081) );
  INV_X4 U1257 ( .A(n1115), .ZN(n1595) );
  INV_X2 U1260 ( .A(n3488), .ZN(n3373) );
  OAI211_X4 U1261 ( .C1(n3130), .C2(n3129), .A(n3128), .B(n3127), .ZN(n3228)
         );
  INV_X8 U1262 ( .A(n1508), .ZN(n3808) );
  NAND3_X2 U1263 ( .A1(n2555), .A2(n2516), .A3(n2515), .ZN(n2399) );
  NAND2_X4 U1264 ( .A1(n1143), .A2(n1144), .ZN(n1146) );
  NAND2_X4 U1265 ( .A1(n1145), .A2(n1146), .ZN(n1978) );
  INV_X4 U1266 ( .A(n1977), .ZN(n1143) );
  NAND2_X4 U1268 ( .A1(n1978), .A2(n1979), .ZN(n2099) );
  INV_X8 U1269 ( .A(n2958), .ZN(n2961) );
  INV_X4 U1271 ( .A(net294085), .ZN(net294198) );
  NAND2_X4 U1273 ( .A1(n3183), .A2(n3185), .ZN(n3003) );
  NOR2_X2 U1274 ( .A1(n3195), .A2(n3194), .ZN(n3196) );
  CLKBUF_X2 U1275 ( .A(n3194), .Z(n1572) );
  INV_X8 U1276 ( .A(n2818), .ZN(n2819) );
  NAND2_X4 U1277 ( .A1(net295934), .A2(n2815), .ZN(n2823) );
  NAND2_X4 U1279 ( .A1(n1304), .A2(n1572), .ZN(n2822) );
  CLKBUF_X3 U1280 ( .A(n2993), .Z(n1148) );
  NAND2_X4 U1281 ( .A1(n2823), .A2(n3191), .ZN(n2824) );
  OAI21_X2 U1282 ( .B1(n2820), .B2(n2821), .A(n2819), .ZN(n1304) );
  NOR2_X4 U1283 ( .A1(n3202), .A2(n3201), .ZN(n3209) );
  XNOR2_X1 U1284 ( .A(n3356), .B(n3447), .ZN(product_out[20]) );
  INV_X2 U1285 ( .A(n3473), .ZN(n1149) );
  XNOR2_X1 U1286 ( .A(n4286), .B(n3624), .ZN(product_out[24]) );
  INV_X8 U1289 ( .A(n3441), .ZN(n1226) );
  INV_X4 U1291 ( .A(n1422), .ZN(n1152) );
  INV_X4 U1293 ( .A(n3334), .ZN(n1153) );
  INV_X4 U1294 ( .A(n1153), .ZN(n1154) );
  INV_X4 U1296 ( .A(n1691), .ZN(n1155) );
  AOI21_X2 U1298 ( .B1(n1175), .B2(n2797), .A(n2846), .ZN(n2804) );
  NAND2_X4 U1299 ( .A1(n3541), .A2(n3574), .ZN(n1161) );
  INV_X8 U1300 ( .A(n2688), .ZN(n2414) );
  OAI21_X4 U1301 ( .B1(n3180), .B2(net297188), .A(n3179), .ZN(n3451) );
  XNOR2_X2 U1302 ( .A(n2812), .B(n2831), .ZN(n1156) );
  INV_X4 U1303 ( .A(n1156), .ZN(n1366) );
  INV_X4 U1304 ( .A(n2812), .ZN(n2832) );
  XNOR2_X2 U1305 ( .A(n2966), .B(n3138), .ZN(n1157) );
  INV_X4 U1306 ( .A(n1199), .ZN(n1158) );
  INV_X8 U1307 ( .A(n1158), .ZN(n1159) );
  NAND2_X4 U1308 ( .A1(net294770), .A2(n3800), .ZN(n3744) );
  NAND4_X2 U1309 ( .A1(n2126), .A2(n1370), .A3(n2229), .A4(n2220), .ZN(n2128)
         );
  NAND2_X2 U1311 ( .A1(n3365), .A2(n3570), .ZN(n3366) );
  NAND2_X4 U1312 ( .A1(n3541), .A2(n3574), .ZN(n1162) );
  NAND2_X4 U1313 ( .A1(n1252), .A2(n1253), .ZN(n3541) );
  INV_X2 U1314 ( .A(n2185), .ZN(n1634) );
  NAND2_X2 U1315 ( .A1(n3476), .A2(n4293), .ZN(n3544) );
  INV_X4 U1316 ( .A(n3777), .ZN(n1197) );
  INV_X4 U1317 ( .A(n3768), .ZN(n3769) );
  NAND2_X4 U1318 ( .A1(n1344), .A2(n1517), .ZN(n3768) );
  NAND2_X4 U1319 ( .A1(n2296), .A2(n2140), .ZN(n1163) );
  NAND2_X2 U1320 ( .A1(n2296), .A2(n2140), .ZN(n2481) );
  INV_X8 U1321 ( .A(n2139), .ZN(n2140) );
  INV_X2 U1322 ( .A(n3336), .ZN(n1164) );
  INV_X2 U1323 ( .A(n1164), .ZN(n1165) );
  INV_X2 U1327 ( .A(net294698), .ZN(net294694) );
  OAI21_X4 U1328 ( .B1(n1638), .B2(n3699), .A(n3698), .ZN(n3705) );
  AOI22_X4 U1329 ( .A1(n3719), .A2(n3718), .B1(n3717), .B2(n3718), .ZN(n3784)
         );
  INV_X2 U1330 ( .A(n1607), .ZN(n1190) );
  NAND2_X4 U1331 ( .A1(n2360), .A2(n2361), .ZN(n2625) );
  XNOR2_X2 U1332 ( .A(n3421), .B(n3420), .ZN(n1169) );
  AOI21_X2 U1334 ( .B1(n2355), .B2(n2515), .A(n2354), .ZN(n2356) );
  NAND2_X2 U1335 ( .A1(n2515), .A2(n2353), .ZN(n2257) );
  XNOR2_X2 U1336 ( .A(n2612), .B(n1194), .ZN(n1555) );
  AND2_X2 U1337 ( .A1(a[23]), .A2(net297485), .ZN(n1170) );
  AND2_X2 U1338 ( .A1(a[27]), .A2(net297485), .ZN(n1171) );
  AND2_X2 U1339 ( .A1(a[29]), .A2(net297485), .ZN(n1172) );
  NOR2_X4 U1340 ( .A1(net296328), .A2(net296329), .ZN(net296430) );
  NOR2_X4 U1341 ( .A1(n2231), .A2(n2230), .ZN(n2072) );
  AND2_X2 U1342 ( .A1(n1508), .A2(n3809), .ZN(n1173) );
  INV_X4 U1343 ( .A(n2956), .ZN(n2757) );
  INV_X2 U1344 ( .A(n1238), .ZN(n1585) );
  INV_X8 U1345 ( .A(n2959), .ZN(n1238) );
  INV_X8 U1346 ( .A(n2490), .ZN(n2338) );
  INV_X8 U1347 ( .A(n1879), .ZN(n1713) );
  INV_X8 U1348 ( .A(n1949), .ZN(n2098) );
  INV_X4 U1349 ( .A(n1775), .ZN(n1194) );
  OAI22_X2 U1350 ( .A1(n2697), .A2(n2757), .B1(n2757), .B2(n2766), .ZN(n1524)
         );
  NAND2_X4 U1351 ( .A1(n3133), .A2(n3132), .ZN(n3065) );
  NAND2_X4 U1352 ( .A1(n2967), .A2(n2968), .ZN(n1199) );
  NAND2_X4 U1353 ( .A1(n2528), .A2(n2527), .ZN(n2626) );
  NOR3_X4 U1354 ( .A1(n3045), .A2(n2937), .A3(n2936), .ZN(n1582) );
  NAND2_X2 U1355 ( .A1(n3324), .A2(n3323), .ZN(n3514) );
  NAND2_X4 U1356 ( .A1(net294843), .A2(net294795), .ZN(net294792) );
  NAND2_X4 U1357 ( .A1(net294317), .A2(n1448), .ZN(net294040) );
  NAND2_X4 U1358 ( .A1(net294300), .A2(net294313), .ZN(net294329) );
  INV_X8 U1359 ( .A(n3877), .ZN(n1334) );
  NOR2_X4 U1360 ( .A1(net294365), .A2(net294308), .ZN(n1400) );
  NAND2_X4 U1361 ( .A1(n3280), .A2(n3283), .ZN(n3014) );
  AND2_X2 U1362 ( .A1(net294068), .A2(net294137), .ZN(n1174) );
  AOI22_X4 U1365 ( .A1(n3624), .A2(n3791), .B1(n3717), .B2(n3791), .ZN(n3714)
         );
  INV_X4 U1366 ( .A(net294042), .ZN(n1233) );
  NAND2_X2 U1367 ( .A1(n1960), .A2(n1959), .ZN(n1965) );
  NAND2_X4 U1369 ( .A1(net294540), .A2(net294541), .ZN(net294801) );
  NAND2_X1 U1370 ( .A1(a[22]), .A2(net297254), .ZN(n1176) );
  NAND2_X4 U1371 ( .A1(n1177), .A2(n3991), .ZN(net294068) );
  INV_X4 U1372 ( .A(n1176), .ZN(n1177) );
  NAND2_X1 U1373 ( .A1(n2708), .A2(n2709), .ZN(n1180) );
  NAND2_X2 U1374 ( .A1(n4236), .A2(n1179), .ZN(n1181) );
  NAND2_X2 U1375 ( .A1(n1180), .A2(n1181), .ZN(n1375) );
  INV_X2 U1377 ( .A(n2709), .ZN(n1179) );
  OAI21_X4 U1379 ( .B1(n2838), .B2(n2839), .A(n1375), .ZN(n2840) );
  AND2_X4 U1380 ( .A1(n2526), .A2(n2654), .ZN(n1690) );
  NOR2_X2 U1381 ( .A1(n2615), .A2(n2563), .ZN(n2513) );
  NAND2_X4 U1384 ( .A1(n3249), .A2(n3065), .ZN(n3137) );
  OAI21_X4 U1385 ( .B1(n2801), .B2(n1231), .A(n2845), .ZN(n2802) );
  NAND2_X2 U1386 ( .A1(net294334), .A2(net294329), .ZN(n1185) );
  NAND2_X4 U1387 ( .A1(n1183), .A2(n1184), .ZN(n1186) );
  NAND2_X4 U1388 ( .A1(n1185), .A2(n1186), .ZN(net294369) );
  INV_X8 U1389 ( .A(net294334), .ZN(n1183) );
  INV_X4 U1390 ( .A(net294329), .ZN(n1184) );
  NAND2_X1 U1391 ( .A1(a[21]), .A2(net297254), .ZN(net294334) );
  INV_X4 U1392 ( .A(n1324), .ZN(n1187) );
  NAND2_X1 U1394 ( .A1(net299066), .A2(net294101), .ZN(n1417) );
  INV_X1 U1398 ( .A(n1677), .ZN(n1188) );
  INV_X4 U1399 ( .A(n1677), .ZN(n1678) );
  AOI21_X2 U1400 ( .B1(n3141), .B2(n3140), .A(n3238), .ZN(n3146) );
  INV_X4 U1401 ( .A(n2971), .ZN(n1239) );
  INV_X4 U1402 ( .A(n3312), .ZN(n1192) );
  CLKBUF_X3 U1403 ( .A(n3786), .Z(n1189) );
  XNOR2_X2 U1404 ( .A(n2241), .B(n2408), .ZN(n1607) );
  NAND2_X4 U1405 ( .A1(n2399), .A2(n1298), .ZN(n2446) );
  INV_X4 U1406 ( .A(n2568), .ZN(n1191) );
  INV_X4 U1407 ( .A(n2568), .ZN(n2469) );
  INV_X1 U1408 ( .A(n1387), .ZN(net298880) );
  NAND2_X2 U1409 ( .A1(n4045), .A2(n3471), .ZN(n3434) );
  NAND2_X2 U1410 ( .A1(n3514), .A2(n3510), .ZN(n3399) );
  NAND2_X4 U1411 ( .A1(n3517), .A2(n3400), .ZN(n3250) );
  NAND2_X2 U1412 ( .A1(n2612), .A2(n1775), .ZN(n1195) );
  NAND2_X4 U1413 ( .A1(n1193), .A2(n1194), .ZN(n1196) );
  NAND2_X4 U1414 ( .A1(n1195), .A2(n1196), .ZN(n1544) );
  INV_X4 U1415 ( .A(n2612), .ZN(n1193) );
  INV_X4 U1416 ( .A(n2196), .ZN(n1526) );
  XNOR2_X2 U1417 ( .A(net294200), .B(n1341), .ZN(net86661) );
  INV_X8 U1419 ( .A(n2749), .ZN(n1339) );
  AOI21_X1 U1421 ( .B1(net294657), .B2(net294656), .A(net294652), .ZN(
        net294649) );
  OAI21_X2 U1422 ( .B1(n2480), .B2(n1626), .A(n1602), .ZN(n2485) );
  CLKBUF_X3 U1423 ( .A(n3163), .Z(n1198) );
  NAND2_X2 U1424 ( .A1(n3672), .A2(net294779), .ZN(net294786) );
  NAND2_X4 U1425 ( .A1(n2334), .A2(n1505), .ZN(n2073) );
  INV_X4 U1427 ( .A(n3173), .ZN(n3223) );
  NAND2_X2 U1428 ( .A1(net295501), .A2(n1104), .ZN(net295382) );
  NAND3_X2 U1429 ( .A1(n1593), .A2(n3569), .A3(n3497), .ZN(n3498) );
  INV_X8 U1430 ( .A(net296337), .ZN(net296416) );
  NAND2_X4 U1431 ( .A1(n2247), .A2(n2248), .ZN(n2249) );
  INV_X4 U1432 ( .A(n2364), .ZN(n2365) );
  XNOR2_X2 U1433 ( .A(n3783), .B(n3782), .ZN(n1623) );
  NAND2_X2 U1434 ( .A1(n2691), .A2(n2690), .ZN(n2761) );
  NAND2_X4 U1435 ( .A1(n2992), .A2(n1148), .ZN(n2826) );
  NAND2_X4 U1436 ( .A1(n2145), .A2(n2146), .ZN(n1493) );
  INV_X8 U1437 ( .A(n1620), .ZN(n1621) );
  NAND2_X4 U1438 ( .A1(n1350), .A2(n4174), .ZN(n4178) );
  AOI21_X4 U1439 ( .B1(net294539), .B2(net294540), .A(net294536), .ZN(n1459)
         );
  INV_X4 U1440 ( .A(net294541), .ZN(net294536) );
  INV_X4 U1441 ( .A(net295029), .ZN(net295028) );
  NAND2_X4 U1442 ( .A1(n1707), .A2(n1708), .ZN(n1710) );
  INV_X8 U1443 ( .A(n1601), .ZN(n1602) );
  NAND2_X1 U1444 ( .A1(net295621), .A2(net295503), .ZN(n1202) );
  NAND2_X2 U1445 ( .A1(n1200), .A2(n1201), .ZN(n1203) );
  NAND2_X2 U1446 ( .A1(n1202), .A2(n1203), .ZN(net295618) );
  INV_X2 U1447 ( .A(net295621), .ZN(n1200) );
  INV_X1 U1448 ( .A(net295503), .ZN(n1201) );
  NAND2_X2 U1449 ( .A1(n3322), .A2(n1113), .ZN(n1206) );
  NAND2_X4 U1450 ( .A1(n1204), .A2(n1205), .ZN(n1207) );
  NAND2_X4 U1451 ( .A1(n1206), .A2(n1207), .ZN(n3324) );
  INV_X4 U1452 ( .A(n3322), .ZN(n1204) );
  NAND2_X2 U1453 ( .A1(n3149), .A2(n3237), .ZN(n1210) );
  NAND2_X4 U1454 ( .A1(n1208), .A2(n1209), .ZN(n1211) );
  NAND2_X4 U1455 ( .A1(n1210), .A2(n1211), .ZN(n3152) );
  INV_X4 U1456 ( .A(n3149), .ZN(n1208) );
  INV_X2 U1457 ( .A(n3237), .ZN(n1209) );
  INV_X2 U1458 ( .A(n3152), .ZN(n3150) );
  INV_X8 U1459 ( .A(n2463), .ZN(n3824) );
  XNOR2_X2 U1460 ( .A(n1297), .B(n2543), .ZN(n2463) );
  OAI21_X4 U1461 ( .B1(n2462), .B2(n2461), .A(n2460), .ZN(n1297) );
  NAND2_X4 U1462 ( .A1(n1701), .A2(n1702), .ZN(n3736) );
  NAND2_X4 U1463 ( .A1(net294784), .A2(n3668), .ZN(n3669) );
  NOR2_X2 U1464 ( .A1(n1934), .A2(n1942), .ZN(n1212) );
  NAND2_X2 U1465 ( .A1(n3392), .A2(n3331), .ZN(n3332) );
  INV_X8 U1466 ( .A(n2009), .ZN(n1951) );
  AOI21_X4 U1467 ( .B1(n2253), .B2(n2252), .A(n2401), .ZN(n2403) );
  NAND2_X4 U1468 ( .A1(n3428), .A2(n3427), .ZN(n3438) );
  INV_X2 U1469 ( .A(n3920), .ZN(n3292) );
  NOR2_X2 U1470 ( .A1(n2530), .A2(n2659), .ZN(n2664) );
  NAND2_X1 U1471 ( .A1(n2565), .A2(n2564), .ZN(n2566) );
  NAND2_X4 U1472 ( .A1(n2793), .A2(n2792), .ZN(n2794) );
  NAND2_X2 U1473 ( .A1(n3579), .A2(n4284), .ZN(n3387) );
  NAND2_X2 U1474 ( .A1(n3335), .A2(n1154), .ZN(n3255) );
  NAND2_X4 U1475 ( .A1(n1216), .A2(n2104), .ZN(n1213) );
  INV_X2 U1476 ( .A(n2777), .ZN(n2776) );
  NAND2_X4 U1477 ( .A1(n2013), .A2(n1627), .ZN(n2058) );
  INV_X8 U1478 ( .A(n1936), .ZN(n1214) );
  INV_X8 U1479 ( .A(n2301), .ZN(n2303) );
  NAND2_X2 U1480 ( .A1(n2670), .A2(n2669), .ZN(n1215) );
  NAND2_X4 U1481 ( .A1(n2018), .A2(n2019), .ZN(n1216) );
  NAND2_X1 U1482 ( .A1(n2018), .A2(n2019), .ZN(n1217) );
  INV_X8 U1483 ( .A(n2021), .ZN(n2018) );
  NAND2_X2 U1484 ( .A1(n1877), .A2(n1876), .ZN(n1220) );
  NAND2_X4 U1485 ( .A1(n1218), .A2(n1219), .ZN(n1221) );
  NAND2_X4 U1486 ( .A1(n1220), .A2(n1221), .ZN(n1642) );
  INV_X4 U1487 ( .A(n1877), .ZN(n1218) );
  INV_X8 U1488 ( .A(n3702), .ZN(n3708) );
  INV_X32 U1489 ( .A(control[1]), .ZN(net297172) );
  NAND2_X2 U1490 ( .A1(n2115), .A2(n2114), .ZN(n1227) );
  NAND2_X4 U1492 ( .A1(n1672), .A2(n1673), .ZN(n1675) );
  INV_X4 U1493 ( .A(n3038), .ZN(n3041) );
  AND3_X4 U1495 ( .A1(n1629), .A2(n2407), .A3(n2432), .ZN(n2340) );
  INV_X4 U1496 ( .A(n3474), .ZN(n1222) );
  NOR2_X4 U1497 ( .A1(n1413), .A2(net293929), .ZN(n1223) );
  NOR2_X4 U1498 ( .A1(net293931), .A2(n1224), .ZN(net293927) );
  INV_X4 U1499 ( .A(n1223), .ZN(n1224) );
  INV_X4 U1500 ( .A(net294100), .ZN(net293929) );
  NAND2_X4 U1502 ( .A1(n1882), .A2(n1940), .ZN(n1225) );
  NAND2_X2 U1503 ( .A1(n1669), .A2(n2234), .ZN(n2017) );
  NAND3_X1 U1505 ( .A1(n3720), .A2(n3785), .A3(n3692), .ZN(n3693) );
  NAND2_X2 U1506 ( .A1(net294701), .A2(n3911), .ZN(n3689) );
  NAND2_X1 U1507 ( .A1(n1387), .A2(net294349), .ZN(net294353) );
  NAND2_X2 U1508 ( .A1(net294349), .A2(n3916), .ZN(net294356) );
  OAI21_X4 U1509 ( .B1(n2462), .B2(n2461), .A(n2460), .ZN(n2541) );
  INV_X8 U1510 ( .A(n2458), .ZN(n2462) );
  NAND2_X4 U1511 ( .A1(n2041), .A2(n2040), .ZN(n2161) );
  INV_X8 U1512 ( .A(n2667), .ZN(n2881) );
  NAND3_X4 U1513 ( .A1(n1569), .A2(n1930), .A3(n1228), .ZN(n1946) );
  INV_X4 U1514 ( .A(n1227), .ZN(n1228) );
  NAND2_X4 U1515 ( .A1(n1946), .A2(n1947), .ZN(n1567) );
  INV_X4 U1516 ( .A(n2692), .ZN(n2584) );
  OAI21_X1 U1517 ( .B1(n1962), .B2(n1961), .A(n1963), .ZN(n1574) );
  INV_X4 U1518 ( .A(n3259), .ZN(n3067) );
  NAND2_X4 U1519 ( .A1(n2760), .A2(n2412), .ZN(n2408) );
  NAND3_X2 U1520 ( .A1(n2758), .A2(n2493), .A3(n1625), .ZN(n1229) );
  NAND3_X2 U1521 ( .A1(n2758), .A2(n2493), .A3(n1625), .ZN(n2692) );
  NAND2_X2 U1522 ( .A1(n2320), .A2(net296672), .ZN(n2205) );
  NAND2_X4 U1523 ( .A1(n3318), .A2(n1645), .ZN(n3322) );
  INV_X8 U1524 ( .A(n1858), .ZN(n1846) );
  INV_X4 U1525 ( .A(n2858), .ZN(n1230) );
  OAI21_X4 U1526 ( .B1(n2704), .B2(n1339), .A(n2788), .ZN(n2858) );
  BUF_X4 U1528 ( .A(n2800), .Z(n1231) );
  NOR2_X4 U1529 ( .A1(n3771), .A2(net297188), .ZN(n3781) );
  NAND2_X4 U1530 ( .A1(n3595), .A2(n3596), .ZN(n3597) );
  NAND2_X4 U1531 ( .A1(n3528), .A2(n3527), .ZN(net294795) );
  INV_X2 U1532 ( .A(n3132), .ZN(n3063) );
  INV_X8 U1533 ( .A(n2789), .ZN(n2753) );
  OAI21_X4 U1536 ( .B1(n2584), .B2(n2497), .A(n2579), .ZN(n2503) );
  NOR2_X2 U1537 ( .A1(n2833), .A2(n2707), .ZN(n1311) );
  NAND2_X4 U1538 ( .A1(n3478), .A2(n1240), .ZN(n3342) );
  INV_X1 U1539 ( .A(n1108), .ZN(n1255) );
  INV_X1 U1540 ( .A(net297862), .ZN(n1232) );
  INV_X2 U1541 ( .A(net293933), .ZN(net297862) );
  INV_X2 U1542 ( .A(n2083), .ZN(n2185) );
  INV_X2 U1543 ( .A(net294770), .ZN(n1408) );
  NAND2_X4 U1544 ( .A1(n1652), .A2(n1653), .ZN(n1655) );
  NAND2_X4 U1545 ( .A1(n2048), .A2(n2047), .ZN(n2029) );
  AND2_X4 U1546 ( .A1(net294313), .A2(n1233), .ZN(net294301) );
  NAND2_X4 U1547 ( .A1(net294217), .A2(n1343), .ZN(n1342) );
  NOR2_X4 U1549 ( .A1(n1868), .A2(n1869), .ZN(n1841) );
  NAND2_X2 U1550 ( .A1(n1919), .A2(n1918), .ZN(n1868) );
  NAND4_X4 U1552 ( .A1(b[25]), .A2(net297172), .A3(a[2]), .A4(net298226), .ZN(
        n1920) );
  OAI21_X2 U1553 ( .B1(net294042), .B2(net294043), .A(net294044), .ZN(
        net294039) );
  OAI21_X4 U1554 ( .B1(net294155), .B2(net294154), .A(net294298), .ZN(n3972)
         );
  AOI21_X4 U1555 ( .B1(n1104), .B2(net295501), .A(n1384), .ZN(net295286) );
  NAND2_X1 U1556 ( .A1(n2347), .A2(n2348), .ZN(n1236) );
  NAND2_X2 U1557 ( .A1(n1234), .A2(n1235), .ZN(n1237) );
  NAND2_X2 U1558 ( .A1(n1237), .A2(n1236), .ZN(n1619) );
  INV_X8 U1559 ( .A(n2347), .ZN(n1234) );
  INV_X4 U1560 ( .A(n2348), .ZN(n1235) );
  INV_X8 U1562 ( .A(n2978), .ZN(n2971) );
  INV_X2 U1563 ( .A(n1161), .ZN(n3738) );
  NAND2_X2 U1564 ( .A1(n1856), .A2(n1855), .ZN(n1849) );
  NAND3_X2 U1565 ( .A1(n2689), .A2(n2687), .A3(n2688), .ZN(n2690) );
  INV_X2 U1566 ( .A(n2952), .ZN(n1542) );
  OAI221_X2 U1567 ( .B1(n3029), .B2(n2669), .C1(n3026), .C2(n2615), .A(n2670), 
        .ZN(n2616) );
  INV_X8 U1568 ( .A(n2287), .ZN(n2401) );
  BUF_X4 U1569 ( .A(n1578), .Z(n1759) );
  NOR2_X2 U1570 ( .A1(n1498), .A2(n3117), .ZN(n3119) );
  NAND2_X4 U1571 ( .A1(n2858), .A2(n2857), .ZN(n2705) );
  NAND2_X4 U1572 ( .A1(n3103), .A2(n1111), .ZN(n2987) );
  NAND2_X4 U1574 ( .A1(n3469), .A2(n3470), .ZN(n1512) );
  NAND2_X2 U1575 ( .A1(n2607), .A2(n2703), .ZN(n2506) );
  NAND2_X4 U1576 ( .A1(n2984), .A2(n2983), .ZN(n3073) );
  NAND2_X4 U1577 ( .A1(n1342), .A2(n1415), .ZN(n1341) );
  INV_X4 U1578 ( .A(n3136), .ZN(n1241) );
  NAND3_X2 U1579 ( .A1(n2949), .A2(n2789), .A3(n2788), .ZN(n2793) );
  INV_X2 U1580 ( .A(n2224), .ZN(n1735) );
  AOI21_X4 U1582 ( .B1(net294326), .B2(net294325), .A(net294198), .ZN(n1385)
         );
  INV_X4 U1583 ( .A(net295032), .ZN(n1435) );
  INV_X8 U1584 ( .A(n3378), .ZN(n3492) );
  INV_X2 U1585 ( .A(n1365), .ZN(n1638) );
  NAND2_X4 U1586 ( .A1(n2930), .A2(n2929), .ZN(n3104) );
  NAND2_X4 U1587 ( .A1(a[2]), .A2(net299325), .ZN(n1834) );
  INV_X4 U1588 ( .A(n2745), .ZN(n1328) );
  INV_X8 U1589 ( .A(n3215), .ZN(n3217) );
  INV_X2 U1590 ( .A(n1887), .ZN(n1888) );
  NAND3_X2 U1591 ( .A1(n2941), .A2(n2940), .A3(n3043), .ZN(n1243) );
  INV_X32 U1592 ( .A(control[0]), .ZN(net297184) );
  INV_X4 U1593 ( .A(n1900), .ZN(n1558) );
  NAND3_X4 U1594 ( .A1(n3281), .A2(n1615), .A3(n1245), .ZN(n3285) );
  INV_X8 U1595 ( .A(n3014), .ZN(n1245) );
  NAND2_X4 U1596 ( .A1(n1485), .A2(net294544), .ZN(net294438) );
  NAND2_X4 U1597 ( .A1(net297002), .A2(n1923), .ZN(n1871) );
  NAND4_X4 U1598 ( .A1(b[24]), .A2(net297640), .A3(a[3]), .A4(net297180), .ZN(
        net297002) );
  INV_X8 U1599 ( .A(net296333), .ZN(n1441) );
  INV_X8 U1600 ( .A(net294841), .ZN(net294930) );
  CLKBUF_X3 U1601 ( .A(n2765), .Z(n1312) );
  NAND2_X2 U1602 ( .A1(n2698), .A2(n1155), .ZN(n1248) );
  NAND2_X4 U1603 ( .A1(n1246), .A2(n1247), .ZN(n1249) );
  NAND2_X4 U1604 ( .A1(n1248), .A2(n1249), .ZN(n1800) );
  INV_X4 U1605 ( .A(n2698), .ZN(n1246) );
  INV_X1 U1606 ( .A(n2755), .ZN(n1247) );
  NOR2_X2 U1607 ( .A1(n1800), .A2(n2850), .ZN(n2853) );
  INV_X2 U1608 ( .A(net296104), .ZN(net296216) );
  OAI21_X4 U1609 ( .B1(n3584), .B2(n3583), .A(n1604), .ZN(n3600) );
  INV_X2 U1611 ( .A(n1599), .ZN(n1895) );
  NAND2_X4 U1612 ( .A1(n3316), .A2(n3315), .ZN(n3478) );
  NAND2_X4 U1613 ( .A1(net296334), .A2(net296333), .ZN(net295990) );
  NAND2_X4 U1614 ( .A1(a[12]), .A2(net297485), .ZN(net296333) );
  INV_X4 U1616 ( .A(n2725), .ZN(n2723) );
  INV_X2 U1617 ( .A(n4251), .ZN(n1477) );
  NAND2_X2 U1618 ( .A1(n3535), .A2(n3534), .ZN(n1252) );
  NAND2_X2 U1619 ( .A1(n1250), .A2(n1251), .ZN(n1253) );
  INV_X4 U1620 ( .A(n3535), .ZN(n1250) );
  INV_X4 U1621 ( .A(n3534), .ZN(n1251) );
  NAND3_X1 U1622 ( .A1(net294137), .A2(net294068), .A3(n4090), .ZN(n4042) );
  NAND2_X4 U1623 ( .A1(n3498), .A2(n3499), .ZN(n3542) );
  NAND2_X4 U1624 ( .A1(net294437), .A2(net294438), .ZN(net294405) );
  AOI21_X2 U1625 ( .B1(net294153), .B2(net294154), .A(net294155), .ZN(n4028)
         );
  NAND2_X4 U1627 ( .A1(n3735), .A2(n3734), .ZN(n3776) );
  NOR2_X2 U1628 ( .A1(n4239), .A2(net299021), .ZN(net294346) );
  INV_X8 U1629 ( .A(n2328), .ZN(n1795) );
  NAND2_X1 U1630 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  NAND2_X4 U1632 ( .A1(n3140), .A2(n3141), .ZN(n2966) );
  OAI22_X4 U1633 ( .A1(b[1]), .A2(net298225), .B1(b[9]), .B2(control[0]), .ZN(
        n1835) );
  OAI21_X4 U1634 ( .B1(n1313), .B2(net297188), .A(n2999), .ZN(n3215) );
  AOI21_X4 U1635 ( .B1(n1953), .B2(n1954), .A(n1952), .ZN(n1955) );
  INV_X4 U1636 ( .A(n3836), .ZN(n3771) );
  NOR2_X4 U1637 ( .A1(n3913), .A2(n3912), .ZN(n3741) );
  NAND2_X2 U1638 ( .A1(net294527), .A2(net294440), .ZN(n1257) );
  INV_X2 U1639 ( .A(net294444), .ZN(n1258) );
  NAND2_X4 U1640 ( .A1(net294531), .A2(net294530), .ZN(net294527) );
  NAND2_X2 U1641 ( .A1(net294527), .A2(net294440), .ZN(net294439) );
  INV_X8 U1642 ( .A(net294440), .ZN(net294444) );
  INV_X8 U1643 ( .A(n2283), .ZN(n1721) );
  NAND2_X2 U1644 ( .A1(n3681), .A2(n3565), .ZN(n3420) );
  NAND2_X4 U1645 ( .A1(n1674), .A2(n1675), .ZN(n2618) );
  NAND2_X2 U1646 ( .A1(n2617), .A2(n2616), .ZN(n1674) );
  NAND2_X2 U1647 ( .A1(n3081), .A2(n1187), .ZN(n1325) );
  NAND3_X2 U1648 ( .A1(n2309), .A2(n1377), .A3(n2310), .ZN(n1609) );
  NAND3_X4 U1649 ( .A1(n1858), .A2(n1859), .A3(n1857), .ZN(n2009) );
  INV_X4 U1650 ( .A(n3826), .ZN(n3180) );
  INV_X4 U1652 ( .A(n2026), .ZN(n2028) );
  AND2_X2 U1653 ( .A1(n3121), .A2(n3231), .ZN(n1500) );
  NAND2_X2 U1654 ( .A1(n4044), .A2(n3560), .ZN(n3348) );
  INV_X8 U1655 ( .A(n3560), .ZN(n3474) );
  INV_X4 U1656 ( .A(net299335), .ZN(net294519) );
  NAND2_X2 U1657 ( .A1(a[10]), .A2(net294188), .ZN(net296539) );
  INV_X4 U1658 ( .A(n2788), .ZN(n1712) );
  INV_X1 U1659 ( .A(n3805), .ZN(n1509) );
  INV_X4 U1662 ( .A(n1404), .ZN(n1403) );
  INV_X4 U1663 ( .A(n1403), .ZN(n1409) );
  OAI21_X2 U1664 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4018) );
  INV_X4 U1665 ( .A(n1853), .ZN(n1554) );
  NOR2_X2 U1666 ( .A1(net294194), .A2(n4034), .ZN(n3983) );
  NAND2_X1 U1668 ( .A1(control[1]), .A2(net297184), .ZN(net297278) );
  NAND2_X1 U1669 ( .A1(control[1]), .A2(net297180), .ZN(net297279) );
  AOI21_X2 U1670 ( .B1(net294515), .B2(n3615), .A(n2896), .ZN(n2897) );
  NOR2_X1 U1671 ( .A1(net294519), .A2(n3618), .ZN(n2896) );
  NOR2_X2 U1672 ( .A1(n1279), .A2(n1413), .ZN(n1418) );
  NAND3_X2 U1673 ( .A1(a[6]), .A2(control[0]), .A3(n1995), .ZN(n2003) );
  INV_X4 U1674 ( .A(n2194), .ZN(n2197) );
  INV_X16 U1675 ( .A(a[8]), .ZN(net298483) );
  INV_X4 U1676 ( .A(net296432), .ZN(net296553) );
  INV_X4 U1677 ( .A(net296221), .ZN(net295991) );
  INV_X4 U1678 ( .A(n2588), .ZN(n2677) );
  NAND2_X2 U1679 ( .A1(n2224), .A2(n1561), .ZN(n1736) );
  NAND2_X1 U1681 ( .A1(net298632), .A2(net295163), .ZN(net295160) );
  INV_X2 U1682 ( .A(n3647), .ZN(n1538) );
  INV_X4 U1683 ( .A(n1793), .ZN(n1794) );
  INV_X4 U1684 ( .A(n2707), .ZN(n2839) );
  OAI21_X2 U1685 ( .B1(n2281), .B2(n2280), .A(n2282), .ZN(n2286) );
  NAND2_X2 U1686 ( .A1(n3317), .A2(n3401), .ZN(n1645) );
  INV_X4 U1687 ( .A(n3159), .ZN(n3162) );
  NAND2_X2 U1688 ( .A1(a[12]), .A2(net297216), .ZN(n3117) );
  NAND2_X2 U1689 ( .A1(a[13]), .A2(net297216), .ZN(n3070) );
  NOR2_X1 U1690 ( .A1(n2922), .A2(n2921), .ZN(n2927) );
  INV_X4 U1691 ( .A(n3230), .ZN(n3384) );
  INV_X4 U1692 ( .A(n3382), .ZN(n3383) );
  INV_X4 U1694 ( .A(n3952), .ZN(n1587) );
  NAND2_X2 U1695 ( .A1(a[17]), .A2(net297216), .ZN(n3415) );
  INV_X8 U1696 ( .A(net297234), .ZN(net297228) );
  INV_X2 U1697 ( .A(n3536), .ZN(n1774) );
  INV_X4 U1698 ( .A(n4011), .ZN(n4141) );
  NAND2_X2 U1699 ( .A1(n1820), .A2(n1819), .ZN(n1825) );
  NOR2_X2 U1700 ( .A1(n4141), .A2(n4140), .ZN(n4142) );
  INV_X4 U1701 ( .A(net297250), .ZN(net297246) );
  INV_X4 U1702 ( .A(net293992), .ZN(net297222) );
  INV_X4 U1703 ( .A(net297222), .ZN(net297218) );
  NAND2_X2 U1704 ( .A1(n2664), .A2(n2663), .ZN(n2666) );
  INV_X4 U1705 ( .A(net294307), .ZN(net294379) );
  OAI21_X2 U1706 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4107) );
  INV_X16 U1708 ( .A(net297250), .ZN(net297244) );
  INV_X16 U1709 ( .A(net297222), .ZN(net297216) );
  INV_X4 U1710 ( .A(net297210), .ZN(net297202) );
  NOR2_X2 U1712 ( .A1(n3462), .A2(n3461), .ZN(n3466) );
  NOR2_X1 U1713 ( .A1(net294126), .A2(n4049), .ZN(n4050) );
  NAND3_X2 U1714 ( .A1(net296808), .A2(n1454), .A3(n1455), .ZN(n1452) );
  NOR2_X2 U1715 ( .A1(n1334), .A2(n1335), .ZN(n1336) );
  INV_X4 U1716 ( .A(net297279), .ZN(net299241) );
  NOR2_X1 U1717 ( .A1(net294126), .A2(n3922), .ZN(n3923) );
  AOI21_X2 U1718 ( .B1(net294039), .B2(net294040), .A(n4098), .ZN(n4099) );
  NOR2_X2 U1719 ( .A1(n3921), .A2(n3290), .ZN(n3291) );
  NOR2_X2 U1720 ( .A1(n1334), .A2(net297188), .ZN(n3619) );
  INV_X4 U1721 ( .A(net294092), .ZN(n1358) );
  NOR2_X2 U1722 ( .A1(n4056), .A2(n4055), .ZN(n4066) );
  NOR2_X2 U1723 ( .A1(n1287), .A2(n3178), .ZN(n3179) );
  INV_X4 U1724 ( .A(net293950), .ZN(net297200) );
  AND2_X4 U1725 ( .A1(a[8]), .A2(net297202), .ZN(n1259) );
  AND2_X2 U1726 ( .A1(a[16]), .A2(net297216), .ZN(n1260) );
  INV_X8 U1727 ( .A(net297200), .ZN(net297198) );
  AND2_X2 U1728 ( .A1(a[24]), .A2(net297204), .ZN(n1261) );
  AND2_X4 U1729 ( .A1(a[6]), .A2(net297254), .ZN(n1262) );
  AND2_X4 U1730 ( .A1(\set_product_in_sig/z1 [25]), .A2(net297190), .ZN(n1263)
         );
  AND2_X2 U1731 ( .A1(a[10]), .A2(net297216), .ZN(n1264) );
  NAND3_X2 U1732 ( .A1(n1893), .A2(n1892), .A3(n1891), .ZN(net294000) );
  INV_X8 U1733 ( .A(net294000), .ZN(net297250) );
  NAND3_X2 U1734 ( .A1(n1969), .A2(n1968), .A3(n1967), .ZN(net293992) );
  AND2_X2 U1735 ( .A1(a[20]), .A2(net297244), .ZN(n1265) );
  NAND3_X2 U1736 ( .A1(n2037), .A2(n2036), .A3(n2035), .ZN(net293989) );
  INV_X4 U1737 ( .A(net293989), .ZN(net297210) );
  NAND2_X1 U1738 ( .A1(a[23]), .A2(net297204), .ZN(net294250) );
  INV_X2 U1739 ( .A(net299020), .ZN(net299021) );
  XOR2_X2 U1740 ( .A(n2873), .B(n1585), .Z(n1266) );
  INV_X4 U1741 ( .A(n2651), .ZN(n2530) );
  AND2_X2 U1742 ( .A1(net295030), .A2(net295377), .ZN(n1267) );
  AND2_X2 U1743 ( .A1(n2324), .A2(n2118), .ZN(n1268) );
  AND2_X4 U1744 ( .A1(a[14]), .A2(net297272), .ZN(n1269) );
  AND2_X2 U1745 ( .A1(net296221), .A2(net297526), .ZN(n1270) );
  XOR2_X2 U1746 ( .A(n3069), .B(n3335), .Z(n1271) );
  AND2_X2 U1747 ( .A1(n2551), .A2(n2638), .ZN(n1272) );
  AND2_X2 U1748 ( .A1(n3511), .A2(n3512), .ZN(n1273) );
  INV_X4 U1749 ( .A(net293924), .ZN(net294093) );
  AND2_X2 U1750 ( .A1(n2064), .A2(n1168), .ZN(n1274) );
  AND2_X2 U1751 ( .A1(n3910), .A2(n4215), .ZN(n1275) );
  AND3_X4 U1753 ( .A1(n2323), .A2(n1556), .A3(n2212), .ZN(n1277) );
  INV_X4 U1755 ( .A(n2099), .ZN(n1770) );
  AND2_X2 U1756 ( .A1(net295742), .A2(n1438), .ZN(n1278) );
  INV_X2 U1757 ( .A(n2367), .ZN(n2370) );
  INV_X8 U1758 ( .A(n1423), .ZN(n1426) );
  INV_X8 U1759 ( .A(net297230), .ZN(net297234) );
  AND2_X4 U1760 ( .A1(\set_product_in_sig/z1 [26]), .A2(net297190), .ZN(n1279)
         );
  AND2_X4 U1761 ( .A1(a[11]), .A2(net297254), .ZN(n1280) );
  AND2_X4 U1762 ( .A1(n3754), .A2(n3805), .ZN(n1281) );
  INV_X4 U1763 ( .A(net297196), .ZN(net297188) );
  AND2_X2 U1764 ( .A1(a[21]), .A2(net297226), .ZN(n1282) );
  AND2_X2 U1765 ( .A1(a[8]), .A2(net297216), .ZN(n1283) );
  AND2_X2 U1766 ( .A1(a[3]), .A2(a[4]), .ZN(n1284) );
  AND2_X4 U1767 ( .A1(\set_product_in_sig/z1 [28]), .A2(net297190), .ZN(n1285)
         );
  AND2_X4 U1768 ( .A1(\set_product_in_sig/z1 [8]), .A2(net297190), .ZN(n1286)
         );
  AND2_X4 U1769 ( .A1(\set_product_in_sig/z1 [19]), .A2(net297188), .ZN(n1287)
         );
  AND2_X4 U1770 ( .A1(\set_product_in_sig/z1 [30]), .A2(net297190), .ZN(n1288)
         );
  AND2_X4 U1771 ( .A1(a[0]), .A2(net297254), .ZN(n1289) );
  XOR2_X2 U1772 ( .A(n1516), .B(n2647), .Z(n1290) );
  AND2_X2 U1773 ( .A1(a[16]), .A2(net297272), .ZN(n1291) );
  AND2_X4 U1774 ( .A1(a[20]), .A2(net297272), .ZN(n1292) );
  AND2_X2 U1775 ( .A1(n3451), .A2(n3439), .ZN(n1293) );
  INV_X2 U1776 ( .A(n2052), .ZN(n2151) );
  AND2_X2 U1777 ( .A1(net295748), .A2(net297526), .ZN(n1294) );
  INV_X4 U1778 ( .A(n1364), .ZN(net297526) );
  INV_X1 U1779 ( .A(net293989), .ZN(n1451) );
  INV_X4 U1780 ( .A(net297210), .ZN(net297204) );
  INV_X8 U1781 ( .A(n1452), .ZN(n1456) );
  INV_X16 U1782 ( .A(n1456), .ZN(net297254) );
  XNOR2_X1 U1783 ( .A(n2898), .B(n3002), .ZN(product_out[16]) );
  XNOR2_X1 U1784 ( .A(n3004), .B(n3006), .ZN(product_out[17]) );
  INV_X4 U1785 ( .A(n2822), .ZN(n2825) );
  NOR2_X4 U1786 ( .A1(n2572), .A2(n2571), .ZN(n2576) );
  NAND2_X2 U1787 ( .A1(n2987), .A2(n2986), .ZN(n1660) );
  INV_X4 U1788 ( .A(n2986), .ZN(n1659) );
  AND2_X2 U1789 ( .A1(n2620), .A2(n2621), .ZN(n1295) );
  NAND2_X4 U1790 ( .A1(a[7]), .A2(net297202), .ZN(n2621) );
  NAND2_X2 U1791 ( .A1(n1303), .A2(n2716), .ZN(n2717) );
  INV_X4 U1792 ( .A(n2729), .ZN(n2737) );
  INV_X8 U1793 ( .A(n2622), .ZN(n2620) );
  NAND2_X4 U1794 ( .A1(n2798), .A2(n1231), .ZN(n2676) );
  NAND2_X4 U1795 ( .A1(n1658), .A2(n1659), .ZN(n1661) );
  INV_X4 U1796 ( .A(n2987), .ZN(n1658) );
  AOI21_X2 U1797 ( .B1(n3182), .B2(n3184), .A(n3181), .ZN(n3189) );
  NAND2_X4 U1798 ( .A1(n2618), .A2(n1283), .ZN(n2667) );
  NAND2_X4 U1799 ( .A1(n3001), .A2(n3002), .ZN(n3183) );
  INV_X2 U1800 ( .A(n3001), .ZN(n2898) );
  OAI21_X4 U1801 ( .B1(n2825), .B2(n2824), .A(n2823), .ZN(n3001) );
  NAND2_X4 U1802 ( .A1(n2811), .A2(n2913), .ZN(n2831) );
  NOR2_X2 U1803 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  CLKBUF_X3 U1805 ( .A(n2276), .Z(n1296) );
  NAND2_X4 U1806 ( .A1(n2366), .A2(n2365), .ZN(n2460) );
  CLKBUF_X2 U1807 ( .A(n2517), .Z(n1298) );
  XNOR2_X2 U1808 ( .A(n2523), .B(n2524), .ZN(n1305) );
  NAND2_X2 U1809 ( .A1(n2476), .A2(n1577), .ZN(n2487) );
  NAND2_X4 U1810 ( .A1(n2181), .A2(n2180), .ZN(n2182) );
  NAND2_X2 U1811 ( .A1(n2152), .A2(n2185), .ZN(n2089) );
  NAND3_X1 U1812 ( .A1(n2477), .A2(n2479), .A3(n2093), .ZN(n2074) );
  XNOR2_X1 U1813 ( .A(n2822), .B(n2824), .ZN(product_out[15]) );
  NAND3_X2 U1814 ( .A1(n3183), .A2(n3184), .A3(n3185), .ZN(n3188) );
  NAND2_X4 U1815 ( .A1(n1798), .A2(n3279), .ZN(n3176) );
  XNOR2_X2 U1817 ( .A(n2808), .B(n2807), .ZN(n1299) );
  CLKBUF_X3 U1818 ( .A(n3181), .Z(n1300) );
  INV_X1 U1820 ( .A(n3045), .ZN(n1301) );
  NAND2_X4 U1821 ( .A1(n3126), .A2(n3125), .ZN(n3071) );
  INV_X2 U1822 ( .A(n1732), .ZN(n1302) );
  INV_X2 U1823 ( .A(n2496), .ZN(n1732) );
  NAND2_X2 U1824 ( .A1(n1550), .A2(n3460), .ZN(n3461) );
  NAND2_X2 U1825 ( .A1(n3222), .A2(n3374), .ZN(n3460) );
  INV_X4 U1826 ( .A(n3494), .ZN(n1549) );
  XOR2_X2 U1827 ( .A(n2713), .B(n2714), .Z(n1303) );
  NAND2_X4 U1828 ( .A1(n2279), .A2(n2278), .ZN(n2149) );
  INV_X4 U1829 ( .A(n1688), .ZN(n2733) );
  INV_X2 U1830 ( .A(n3434), .ZN(n3427) );
  XNOR2_X1 U1831 ( .A(n3443), .B(n3555), .ZN(product_out[22]) );
  NAND2_X4 U1832 ( .A1(n3555), .A2(n4059), .ZN(n3862) );
  INV_X1 U1833 ( .A(net298860), .ZN(n1421) );
  INV_X1 U1834 ( .A(n2636), .ZN(n1618) );
  NAND2_X4 U1835 ( .A1(n2258), .A2(n2259), .ZN(n2527) );
  NAND2_X2 U1837 ( .A1(n1354), .A2(n1760), .ZN(n1762) );
  NOR2_X2 U1838 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
  INV_X8 U1839 ( .A(n2817), .ZN(n2820) );
  NAND3_X4 U1841 ( .A1(n3160), .A2(n3162), .A3(n4269), .ZN(n1540) );
  INV_X2 U1842 ( .A(n3246), .ZN(n3155) );
  NAND3_X2 U1843 ( .A1(n2662), .A2(n2660), .A3(n2661), .ZN(n2663) );
  NAND3_X2 U1844 ( .A1(n2661), .A2(n2528), .A3(n2527), .ZN(n2451) );
  NOR2_X1 U1845 ( .A1(n1387), .A2(net294485), .ZN(net294484) );
  INV_X4 U1846 ( .A(n2251), .ZN(n2252) );
  INV_X4 U1847 ( .A(n3257), .ZN(n1307) );
  INV_X4 U1848 ( .A(n2495), .ZN(n2421) );
  INV_X2 U1849 ( .A(n1362), .ZN(n3238) );
  XNOR2_X2 U1851 ( .A(n2311), .B(n2080), .ZN(n1308) );
  NAND2_X4 U1852 ( .A1(n2287), .A2(n2285), .ZN(n2178) );
  NAND2_X4 U1853 ( .A1(n3236), .A2(n3237), .ZN(n3241) );
  INV_X4 U1854 ( .A(n2525), .ZN(n2526) );
  XNOR2_X2 U1855 ( .A(n2347), .B(n2348), .ZN(n1310) );
  NAND2_X4 U1856 ( .A1(n2678), .A2(n2677), .ZN(net295749) );
  NAND2_X4 U1857 ( .A1(n1269), .A2(n1468), .ZN(net295750) );
  CLKBUF_X3 U1858 ( .A(n2841), .Z(n1776) );
  INV_X2 U1859 ( .A(n2556), .ZN(n2444) );
  INV_X8 U1860 ( .A(n3123), .ZN(n3229) );
  NAND2_X4 U1861 ( .A1(n2289), .A2(n2290), .ZN(n2348) );
  OAI21_X2 U1862 ( .B1(n1270), .B2(n2593), .A(net295754), .ZN(n2591) );
  OAI211_X2 U1863 ( .C1(n1270), .C2(n2593), .A(n2771), .B(net295754), .ZN(
        n2594) );
  XNOR2_X2 U1864 ( .A(n2997), .B(n2998), .ZN(n1313) );
  NAND2_X4 U1865 ( .A1(n3113), .A2(n3114), .ZN(n3121) );
  OAI211_X4 U1866 ( .C1(n3442), .C2(n3449), .A(n3441), .B(n3858), .ZN(n1353)
         );
  NAND2_X2 U1867 ( .A1(n2235), .A2(n2234), .ZN(n2236) );
  NAND2_X1 U1868 ( .A1(n2131), .A2(n2234), .ZN(n2132) );
  AOI21_X2 U1869 ( .B1(n3636), .B2(n3635), .A(n3634), .ZN(n3696) );
  NAND2_X2 U1870 ( .A1(n3876), .A2(n1336), .ZN(n1337) );
  INV_X8 U1871 ( .A(n2755), .ZN(n1691) );
  INV_X4 U1872 ( .A(net294324), .ZN(net294199) );
  NAND2_X4 U1873 ( .A1(n1704), .A2(n1314), .ZN(n2342) );
  CLKBUF_X3 U1874 ( .A(net294309), .Z(net298857) );
  NAND2_X2 U1875 ( .A1(net294388), .A2(n3767), .ZN(n1344) );
  INV_X2 U1876 ( .A(n2693), .ZN(n1801) );
  NAND3_X2 U1877 ( .A1(n3987), .A2(net299137), .A3(n3988), .ZN(n3986) );
  NOR2_X1 U1878 ( .A1(net296419), .A2(net296418), .ZN(n2420) );
  NAND2_X2 U1880 ( .A1(n2183), .A2(n2182), .ZN(n1317) );
  NAND2_X4 U1881 ( .A1(n1315), .A2(n1316), .ZN(n1318) );
  NAND2_X2 U1882 ( .A1(n1317), .A2(n1318), .ZN(n2187) );
  INV_X4 U1883 ( .A(n2183), .ZN(n1315) );
  INV_X4 U1884 ( .A(n2182), .ZN(n1316) );
  NAND2_X2 U1885 ( .A1(n1671), .A2(n2138), .ZN(n1321) );
  NAND2_X4 U1886 ( .A1(n1319), .A2(n1320), .ZN(n1322) );
  NAND2_X4 U1887 ( .A1(n1321), .A2(n1322), .ZN(n2139) );
  INV_X4 U1888 ( .A(n2138), .ZN(n1319) );
  INV_X4 U1889 ( .A(n1671), .ZN(n1320) );
  INV_X2 U1890 ( .A(n1670), .ZN(n1671) );
  NAND2_X2 U1891 ( .A1(n2298), .A2(n2139), .ZN(n2248) );
  INV_X2 U1892 ( .A(n3137), .ZN(n1653) );
  NAND2_X2 U1893 ( .A1(n1323), .A2(n1324), .ZN(n1326) );
  NAND2_X4 U1894 ( .A1(n1325), .A2(n1326), .ZN(n3082) );
  INV_X4 U1895 ( .A(n3081), .ZN(n1323) );
  NAND2_X4 U1896 ( .A1(n1327), .A2(n1328), .ZN(n1330) );
  NAND2_X4 U1897 ( .A1(n1330), .A2(n1329), .ZN(n2622) );
  INV_X4 U1898 ( .A(n2619), .ZN(n1327) );
  INV_X2 U1899 ( .A(n1760), .ZN(n1331) );
  NAND2_X4 U1901 ( .A1(n3056), .A2(n3141), .ZN(n3236) );
  NAND2_X4 U1902 ( .A1(n4098), .A2(n4085), .ZN(n4086) );
  NAND2_X2 U1903 ( .A1(net294326), .A2(net294325), .ZN(net294324) );
  INV_X1 U1904 ( .A(net295737), .ZN(net295736) );
  INV_X8 U1905 ( .A(n3873), .ZN(n3876) );
  NAND2_X4 U1906 ( .A1(n3079), .A2(n3078), .ZN(n1332) );
  NAND2_X2 U1908 ( .A1(n3791), .A2(n4061), .ZN(n3716) );
  NAND2_X2 U1909 ( .A1(n3623), .A2(n1611), .ZN(n3791) );
  NOR2_X4 U1910 ( .A1(n3786), .A2(n1333), .ZN(n3795) );
  NAND2_X1 U1911 ( .A1(n1335), .A2(n1263), .ZN(n1333) );
  NOR2_X4 U1912 ( .A1(n3795), .A2(n3794), .ZN(n3796) );
  INV_X4 U1915 ( .A(n3785), .ZN(n1335) );
  NAND2_X2 U1916 ( .A1(n2655), .A2(n2656), .ZN(n2657) );
  OAI22_X4 U1917 ( .A1(b[1]), .A2(net297182), .B1(b[9]), .B2(control[0]), .ZN(
        n1815) );
  OAI21_X2 U1918 ( .B1(n2097), .B2(n2098), .A(n2096), .ZN(n2101) );
  OAI211_X2 U1919 ( .C1(n4063), .C2(n4062), .A(n4060), .B(n4061), .ZN(n4064)
         );
  OAI21_X4 U1920 ( .B1(n2704), .B2(n1339), .A(n2788), .ZN(n1338) );
  INV_X8 U1921 ( .A(n2747), .ZN(n2749) );
  INV_X2 U1922 ( .A(n2111), .ZN(n1564) );
  NAND2_X4 U1923 ( .A1(a[10]), .A2(net297244), .ZN(n2707) );
  NAND2_X4 U1925 ( .A1(n2032), .A2(n2031), .ZN(n2044) );
  INV_X2 U1926 ( .A(net294308), .ZN(net294320) );
  NAND2_X2 U1927 ( .A1(n2883), .A2(n2917), .ZN(n2919) );
  OAI21_X4 U1928 ( .B1(n1536), .B2(n3379), .A(n3377), .ZN(n3380) );
  INV_X2 U1929 ( .A(n3514), .ZN(n3583) );
  INV_X8 U1930 ( .A(n1798), .ZN(n3468) );
  AOI21_X2 U1931 ( .B1(n1262), .B2(n2732), .A(n2731), .ZN(n2735) );
  NAND2_X4 U1932 ( .A1(n2732), .A2(n1262), .ZN(n2718) );
  INV_X4 U1933 ( .A(net295503), .ZN(net298907) );
  NAND3_X2 U1934 ( .A1(n3630), .A2(n3629), .A3(n3475), .ZN(n3476) );
  NAND2_X4 U1935 ( .A1(n1279), .A2(n1422), .ZN(net294100) );
  NAND2_X2 U1936 ( .A1(n2671), .A2(n3027), .ZN(n2617) );
  INV_X8 U1937 ( .A(n3281), .ZN(n3096) );
  INV_X4 U1938 ( .A(n3235), .ZN(n3243) );
  XNOR2_X2 U1939 ( .A(n2710), .B(n2801), .ZN(n1340) );
  NAND2_X4 U1940 ( .A1(net297774), .A2(n1405), .ZN(net294882) );
  NAND2_X4 U1941 ( .A1(n3533), .A2(net297774), .ZN(n3606) );
  NAND2_X2 U1942 ( .A1(n2849), .A2(n2938), .ZN(n2924) );
  INV_X4 U1943 ( .A(n1414), .ZN(n1343) );
  OAI21_X2 U1944 ( .B1(n1418), .B2(n1419), .A(net299066), .ZN(n1414) );
  NAND2_X2 U1945 ( .A1(n1729), .A2(n1730), .ZN(n2880) );
  INV_X4 U1946 ( .A(n1768), .ZN(n3907) );
  XNOR2_X2 U1947 ( .A(net296530), .B(net296425), .ZN(n1345) );
  NAND2_X4 U1950 ( .A1(n2482), .A2(n2481), .ZN(n1793) );
  OAI21_X2 U1951 ( .B1(n2556), .B2(n2557), .A(n2555), .ZN(n2559) );
  INV_X4 U1952 ( .A(n1635), .ZN(n3613) );
  NOR2_X4 U1953 ( .A1(n1402), .A2(net294450), .ZN(net294441) );
  NOR2_X4 U1954 ( .A1(n1348), .A2(n1264), .ZN(n1347) );
  INV_X8 U1955 ( .A(n1347), .ZN(n3128) );
  XNOR2_X2 U1956 ( .A(n2805), .B(n1776), .ZN(n1348) );
  NAND3_X2 U1957 ( .A1(n4078), .A2(net294040), .A3(n4077), .ZN(n4081) );
  XNOR2_X2 U1958 ( .A(n4152), .B(n1261), .ZN(n1349) );
  XNOR2_X2 U1959 ( .A(n4173), .B(n1288), .ZN(n1350) );
  NAND2_X2 U1960 ( .A1(net294346), .A2(net299047), .ZN(n3927) );
  INV_X4 U1961 ( .A(n2616), .ZN(n1673) );
  XNOR2_X2 U1962 ( .A(n2190), .B(n2052), .ZN(n2082) );
  INV_X4 U1963 ( .A(n2190), .ZN(n2283) );
  NAND2_X2 U1964 ( .A1(n3128), .A2(n3124), .ZN(n2807) );
  NAND2_X2 U1965 ( .A1(n1449), .A2(net294249), .ZN(net294402) );
  XNOR2_X2 U1966 ( .A(n2142), .B(n2141), .ZN(n1351) );
  XNOR2_X2 U1967 ( .A(n3417), .B(net299334), .ZN(n1352) );
  NAND2_X4 U1968 ( .A1(n2478), .A2(n2477), .ZN(n2311) );
  NAND2_X2 U1969 ( .A1(n3017), .A2(n3099), .ZN(n3019) );
  INV_X2 U1970 ( .A(n2881), .ZN(n1720) );
  INV_X4 U1971 ( .A(n3855), .ZN(n3442) );
  NOR2_X2 U1972 ( .A1(n4072), .A2(n4071), .ZN(n1355) );
  NAND2_X4 U1973 ( .A1(n4070), .A2(n1357), .ZN(n1356) );
  NAND2_X2 U1974 ( .A1(n1358), .A2(net293924), .ZN(n1357) );
  XNOR2_X2 U1975 ( .A(n2714), .B(n2713), .ZN(n1359) );
  NAND2_X4 U1976 ( .A1(n1628), .A2(n3271), .ZN(n1360) );
  OAI22_X4 U1978 ( .A1(n2268), .A2(net297278), .B1(n3637), .B2(net297190), 
        .ZN(n2270) );
  NAND2_X4 U1979 ( .A1(n3700), .A2(n3699), .ZN(n3625) );
  OAI21_X2 U1980 ( .B1(n3700), .B2(n3699), .A(n3697), .ZN(n3704) );
  OAI21_X4 U1982 ( .B1(n1763), .B2(n3877), .A(net297196), .ZN(n3724) );
  NAND2_X4 U1984 ( .A1(n2622), .A2(n2623), .ZN(n2908) );
  NAND2_X2 U1985 ( .A1(n2700), .A2(n1134), .ZN(n2488) );
  NAND2_X2 U1986 ( .A1(n1622), .A2(n2903), .ZN(n2739) );
  OAI21_X4 U1987 ( .B1(n2903), .B2(n1690), .A(n1622), .ZN(n2714) );
  NOR2_X4 U1989 ( .A1(n3138), .A2(n3139), .ZN(n1362) );
  NAND2_X4 U1992 ( .A1(n3294), .A2(n3293), .ZN(n3447) );
  NAND2_X4 U1993 ( .A1(n4059), .A2(n3552), .ZN(n3863) );
  NAND2_X4 U1994 ( .A1(\set_product_in_sig/z1 [21]), .A2(n3350), .ZN(n3552) );
  NAND2_X4 U1995 ( .A1(n2668), .A2(n1720), .ZN(n2712) );
  NAND2_X4 U1996 ( .A1(n4161), .A2(n4160), .ZN(n4169) );
  NAND2_X4 U1997 ( .A1(a[3]), .A2(net297218), .ZN(n2180) );
  INV_X4 U1998 ( .A(n3167), .ZN(n3168) );
  NOR2_X4 U1999 ( .A1(n1230), .A2(n2834), .ZN(n2836) );
  INV_X2 U2000 ( .A(n1714), .ZN(n1715) );
  NOR2_X4 U2001 ( .A1(net296424), .A2(n1483), .ZN(n1364) );
  NAND2_X4 U2002 ( .A1(n2996), .A2(n1502), .ZN(n2997) );
  INV_X4 U2003 ( .A(n3103), .ZN(n3020) );
  AOI21_X2 U2004 ( .B1(n3847), .B2(n3848), .A(n4069), .ZN(n3851) );
  NOR2_X4 U2005 ( .A1(n1938), .A2(n1941), .ZN(n1939) );
  NAND2_X2 U2006 ( .A1(n3509), .A2(n1165), .ZN(n3337) );
  XNOR2_X2 U2007 ( .A(n4034), .B(n4037), .ZN(n3997) );
  NAND2_X4 U2008 ( .A1(n3549), .A2(n3789), .ZN(n4055) );
  NAND2_X4 U2009 ( .A1(n3548), .A2(n3547), .ZN(n3789) );
  NOR2_X2 U2010 ( .A1(n3089), .A2(n3011), .ZN(n2998) );
  NAND2_X4 U2011 ( .A1(n3018), .A2(n3017), .ZN(n2986) );
  NAND2_X4 U2012 ( .A1(n3107), .A2(n2985), .ZN(n3017) );
  XNOR2_X2 U2013 ( .A(n3542), .B(n3738), .ZN(n1365) );
  NAND2_X4 U2014 ( .A1(n3298), .A2(n3425), .ZN(n3299) );
  INV_X4 U2015 ( .A(n3528), .ZN(n3529) );
  INV_X8 U2016 ( .A(n3227), .ZN(n3308) );
  INV_X2 U2017 ( .A(net294332), .ZN(n1478) );
  AOI21_X4 U2018 ( .B1(n3928), .B2(n3927), .A(n3996), .ZN(n3929) );
  INV_X1 U2019 ( .A(n1501), .ZN(n3996) );
  OAI22_X4 U2021 ( .A1(n3096), .A2(n3014), .B1(n3015), .B2(n3016), .ZN(n3085)
         );
  NAND2_X4 U2022 ( .A1(n1635), .A2(n3697), .ZN(n3877) );
  NAND3_X2 U2023 ( .A1(n1217), .A2(n2053), .A3(n1771), .ZN(n2079) );
  NAND2_X4 U2024 ( .A1(n3390), .A2(n3389), .ZN(n3417) );
  NOR2_X4 U2025 ( .A1(n3376), .A2(n3375), .ZN(n3377) );
  NAND4_X2 U2026 ( .A1(n2585), .A2(net297526), .A3(net295748), .A4(n2499), 
        .ZN(n2500) );
  XNOR2_X2 U2027 ( .A(n4290), .B(n3910), .ZN(n1635) );
  NAND2_X4 U2028 ( .A1(net294080), .A2(net294082), .ZN(n1367) );
  NAND2_X4 U2029 ( .A1(net294081), .A2(net294083), .ZN(n1368) );
  NOR2_X4 U2030 ( .A1(n1367), .A2(n1368), .ZN(n1369) );
  CLKBUF_X3 U2031 ( .A(n3280), .Z(n1502) );
  NAND2_X1 U2032 ( .A1(n1470), .A2(net293935), .ZN(net294219) );
  OAI21_X4 U2033 ( .B1(n3259), .B2(n1307), .A(n3258), .ZN(n3328) );
  AOI21_X4 U2034 ( .B1(n3071), .B2(n3128), .A(n3072), .ZN(n2886) );
  NOR2_X2 U2035 ( .A1(n3072), .A2(n2928), .ZN(n2929) );
  NAND2_X2 U2037 ( .A1(n2700), .A2(n2701), .ZN(n2486) );
  NAND2_X4 U2038 ( .A1(n1735), .A2(n2199), .ZN(n1737) );
  INV_X1 U2039 ( .A(n2937), .ZN(n1714) );
  OAI211_X4 U2040 ( .C1(n1801), .C2(n2954), .A(n1132), .B(n2957), .ZN(n2869)
         );
  NAND3_X2 U2041 ( .A1(n2119), .A2(n2117), .A3(n1643), .ZN(n1370) );
  NAND2_X4 U2042 ( .A1(a[2]), .A2(net297230), .ZN(n1975) );
  NAND2_X4 U2043 ( .A1(n1920), .A2(n1928), .ZN(n1869) );
  XNOR2_X1 U2044 ( .A(n1818), .B(n1372), .ZN(n1371) );
  INV_X8 U2045 ( .A(n1817), .ZN(n1630) );
  OAI21_X2 U2046 ( .B1(n2098), .B2(n2097), .A(n2096), .ZN(n1711) );
  NAND2_X4 U2047 ( .A1(n1555), .A2(n2613), .ZN(n3027) );
  NAND2_X4 U2048 ( .A1(n2440), .A2(n2439), .ZN(n1373) );
  NAND2_X4 U2049 ( .A1(n2248), .A2(n1163), .ZN(n2141) );
  NOR2_X4 U2050 ( .A1(n1632), .A2(n2303), .ZN(n2307) );
  NAND2_X2 U2051 ( .A1(n3520), .A2(n3596), .ZN(n3407) );
  INV_X4 U2052 ( .A(n2917), .ZN(n1518) );
  NAND2_X2 U2053 ( .A1(n2009), .A2(n1642), .ZN(n2011) );
  XNOR2_X1 U2054 ( .A(n2612), .B(n1775), .ZN(n1374) );
  INV_X2 U2056 ( .A(n4061), .ZN(n3866) );
  NAND2_X1 U2057 ( .A1(net295756), .A2(net295750), .ZN(net295513) );
  NAND2_X2 U2058 ( .A1(n2067), .A2(n1556), .ZN(n2068) );
  INV_X4 U2059 ( .A(n2533), .ZN(n2536) );
  INV_X2 U2060 ( .A(n3374), .ZN(n3375) );
  INV_X1 U2061 ( .A(net294054), .ZN(net294981) );
  XNOR2_X2 U2062 ( .A(n3799), .B(n3831), .ZN(n3691) );
  NAND2_X1 U2063 ( .A1(a[18]), .A2(net297254), .ZN(n3830) );
  XNOR2_X2 U2065 ( .A(n3171), .B(n3170), .ZN(n1376) );
  OAI22_X4 U2066 ( .A1(n2308), .A2(n2307), .B1(n2306), .B2(n1213), .ZN(n1377)
         );
  OAI22_X4 U2067 ( .A1(b[0]), .A2(net297184), .B1(b[8]), .B2(control[0]), .ZN(
        n1831) );
  INV_X4 U2068 ( .A(n2491), .ZN(n2336) );
  NAND2_X2 U2069 ( .A1(n3144), .A2(n3059), .ZN(n3062) );
  NAND2_X4 U2070 ( .A1(n2225), .A2(net296324), .ZN(n2320) );
  NAND2_X4 U2071 ( .A1(n1604), .A2(n3513), .ZN(n3413) );
  XNOR2_X2 U2073 ( .A(n2333), .B(n2493), .ZN(n1378) );
  NAND2_X4 U2074 ( .A1(n3987), .A2(n3988), .ZN(n3989) );
  NAND2_X4 U2076 ( .A1(n1360), .A2(n1361), .ZN(n3463) );
  NAND2_X4 U2077 ( .A1(n4208), .A2(n1602), .ZN(n2142) );
  OAI22_X2 U2079 ( .A1(net294980), .A2(net294519), .B1(net294981), .B2(
        net297278), .ZN(n3547) );
  XNOR2_X2 U2080 ( .A(n2168), .B(n1289), .ZN(net294980) );
  NAND2_X4 U2081 ( .A1(n2870), .A2(n2869), .ZN(n2873) );
  NAND2_X4 U2082 ( .A1(n1529), .A2(n1527), .ZN(n1942) );
  INV_X2 U2083 ( .A(n2053), .ZN(n1962) );
  OAI21_X2 U2084 ( .B1(n2206), .B2(n1796), .A(n2212), .ZN(n2207) );
  NAND2_X4 U2085 ( .A1(n1169), .A2(n3422), .ZN(n3630) );
  INV_X4 U2086 ( .A(net295759), .ZN(net295864) );
  NAND2_X4 U2087 ( .A1(n4289), .A2(n3536), .ZN(net299334) );
  NAND3_X2 U2088 ( .A1(n4262), .A2(n2287), .A3(n2400), .ZN(n2290) );
  NAND2_X4 U2090 ( .A1(n2404), .A2(n2400), .ZN(n2288) );
  INV_X8 U2091 ( .A(n2112), .ZN(n2126) );
  NOR2_X4 U2092 ( .A1(n2835), .A2(n2707), .ZN(n2709) );
  NOR2_X2 U2093 ( .A1(net295514), .A2(net295515), .ZN(n1412) );
  OAI22_X4 U2096 ( .A1(b[17]), .A2(net297182), .B1(b[25]), .B2(control[0]), 
        .ZN(n1813) );
  NAND2_X2 U2097 ( .A1(n2191), .A2(n1721), .ZN(n2181) );
  OAI21_X4 U2098 ( .B1(n1875), .B2(n1874), .A(net297009), .ZN(n2195) );
  INV_X2 U2099 ( .A(n1650), .ZN(n1874) );
  OAI221_X4 U2101 ( .B1(n3243), .B2(n3242), .C1(n3241), .C2(n3240), .A(
        net295393), .ZN(net295291) );
  OAI221_X4 U2102 ( .B1(n1490), .B2(net295275), .C1(n1435), .C2(n1436), .A(
        net295028), .ZN(net294820) );
  NAND3_X2 U2103 ( .A1(n1127), .A2(n3314), .A3(n3382), .ZN(n3315) );
  NAND2_X4 U2104 ( .A1(n3409), .A2(n3410), .ZN(n3513) );
  XNOR2_X2 U2105 ( .A(n2362), .B(n2626), .ZN(n2364) );
  AOI21_X4 U2106 ( .B1(n2327), .B2(n2198), .A(net296427), .ZN(n2332) );
  NAND3_X4 U2107 ( .A1(n1379), .A2(n1380), .A3(b[25]), .ZN(net297154) );
  INV_X8 U2108 ( .A(control[0]), .ZN(n1379) );
  INV_X32 U2109 ( .A(control[1]), .ZN(n1380) );
  INV_X2 U2110 ( .A(n2250), .ZN(n2253) );
  NAND2_X2 U2111 ( .A1(n3157), .A2(n1592), .ZN(n3336) );
  OAI211_X4 U2112 ( .C1(n1381), .C2(n3599), .A(n3598), .B(net294913), .ZN(
        net294908) );
  INV_X1 U2113 ( .A(n3526), .ZN(n1381) );
  NAND3_X4 U2114 ( .A1(n1729), .A2(n1730), .A3(n2923), .ZN(n3116) );
  INV_X2 U2115 ( .A(n2922), .ZN(n2923) );
  NAND3_X2 U2116 ( .A1(net294088), .A2(net294085), .A3(net294087), .ZN(
        net294080) );
  NAND2_X4 U2117 ( .A1(n1661), .A2(n1660), .ZN(n2989) );
  XNOR2_X2 U2118 ( .A(n2065), .B(net296842), .ZN(n2328) );
  NAND2_X4 U2119 ( .A1(n2512), .A2(n2563), .ZN(n2560) );
  NAND2_X4 U2120 ( .A1(n4202), .A2(n2684), .ZN(n2765) );
  NAND2_X4 U2121 ( .A1(n3160), .A2(n3047), .ZN(n3331) );
  OAI211_X2 U2122 ( .C1(net294652), .C2(net294653), .A(net294651), .B(n1488), 
        .ZN(net294650) );
  XNOR2_X2 U2124 ( .A(n2441), .B(n2442), .ZN(n2556) );
  NOR2_X4 U2125 ( .A1(n1934), .A2(n1942), .ZN(n1935) );
  INV_X4 U2126 ( .A(n1933), .ZN(n1934) );
  NOR2_X4 U2127 ( .A1(n4205), .A2(n1260), .ZN(n1382) );
  INV_X8 U2128 ( .A(n1382), .ZN(net294779) );
  AOI22_X2 U2129 ( .A1(n3682), .A2(n3683), .B1(n3418), .B2(n3419), .ZN(n3729)
         );
  INV_X4 U2130 ( .A(n3540), .ZN(n3683) );
  NAND2_X2 U2131 ( .A1(n1764), .A2(n2004), .ZN(n1783) );
  NOR2_X2 U2132 ( .A1(n3708), .A2(n3707), .ZN(n1383) );
  INV_X2 U2133 ( .A(n1383), .ZN(n3568) );
  INV_X1 U2134 ( .A(n1442), .ZN(n1384) );
  OAI22_X4 U2135 ( .A1(n4048), .A2(net293950), .B1(n4049), .B2(net297279), 
        .ZN(n2725) );
  OAI21_X4 U2136 ( .B1(n3506), .B2(n3505), .A(n3683), .ZN(n3535) );
  XNOR2_X2 U2137 ( .A(n2997), .B(n2998), .ZN(n3642) );
  INV_X1 U2138 ( .A(net295277), .ZN(n1490) );
  INV_X4 U2139 ( .A(net295278), .ZN(net295275) );
  OAI21_X2 U2141 ( .B1(net294199), .B2(n4238), .A(net294083), .ZN(net294137)
         );
  NAND2_X4 U2142 ( .A1(n1386), .A2(net294327), .ZN(net294085) );
  NAND2_X2 U2143 ( .A1(net298730), .A2(net294085), .ZN(net294082) );
  XNOR2_X2 U2144 ( .A(net294196), .B(n4285), .ZN(n1386) );
  INV_X4 U2145 ( .A(net294334), .ZN(net294327) );
  NOR2_X4 U2146 ( .A1(net294086), .A2(net294084), .ZN(net294325) );
  XNOR2_X2 U2147 ( .A(net294369), .B(net294355), .ZN(net294084) );
  NAND3_X2 U2148 ( .A1(net294372), .A2(net294371), .A3(net294370), .ZN(
        net294355) );
  INV_X8 U2149 ( .A(net294347), .ZN(net294086) );
  NAND2_X4 U2150 ( .A1(n1387), .A2(net294349), .ZN(net294347) );
  NAND2_X4 U2154 ( .A1(n1388), .A2(net294396), .ZN(net294314) );
  XNOR2_X2 U2155 ( .A(net294526), .B(n1257), .ZN(n1393) );
  NAND2_X4 U2156 ( .A1(net297153), .A2(net297154), .ZN(net297152) );
  NAND2_X2 U2157 ( .A1(a[9]), .A2(net297272), .ZN(n1394) );
  NAND2_X2 U2158 ( .A1(n1394), .A2(net296539), .ZN(net296537) );
  INV_X32 U2159 ( .A(net297276), .ZN(net297272) );
  INV_X16 U2160 ( .A(net294187), .ZN(net297276) );
  NAND2_X4 U2161 ( .A1(net297070), .A2(net297071), .ZN(net294187) );
  NAND2_X4 U2162 ( .A1(net294187), .A2(a[6]), .ZN(net296842) );
  INV_X8 U2163 ( .A(net297152), .ZN(net297070) );
  NAND2_X4 U2164 ( .A1(net297070), .A2(net297071), .ZN(net296932) );
  NAND2_X4 U2165 ( .A1(net297070), .A2(net298916), .ZN(net297515) );
  NAND3_X2 U2166 ( .A1(control[0]), .A2(net299325), .A3(b[17]), .ZN(net297153)
         );
  INV_X32 U2167 ( .A(control[1]), .ZN(net299325) );
  NOR2_X4 U2168 ( .A1(net294444), .A2(n1396), .ZN(n1395) );
  OAI21_X4 U2169 ( .B1(net294441), .B2(net294442), .A(n1395), .ZN(net294247)
         );
  NAND2_X4 U2171 ( .A1(net298716), .A2(n1397), .ZN(net294639) );
  NAND2_X4 U2172 ( .A1(net294577), .A2(net294639), .ZN(net294636) );
  INV_X4 U2173 ( .A(net294640), .ZN(n1397) );
  NAND2_X2 U2174 ( .A1(n1397), .A2(net298716), .ZN(net294446) );
  NAND2_X4 U2175 ( .A1(net294529), .A2(net294528), .ZN(net294440) );
  NAND2_X4 U2176 ( .A1(net294439), .A2(n1258), .ZN(net294248) );
  INV_X4 U2177 ( .A(net294530), .ZN(net294528) );
  INV_X2 U2179 ( .A(net294529), .ZN(net294531) );
  INV_X4 U2180 ( .A(net294525), .ZN(net294396) );
  OAI21_X2 U2181 ( .B1(n1400), .B2(n1401), .A(net294322), .ZN(net294520) );
  NAND2_X1 U2182 ( .A1(n1399), .A2(net294310), .ZN(n1401) );
  INV_X8 U2183 ( .A(n1398), .ZN(n1399) );
  AOI21_X4 U2184 ( .B1(n1399), .B2(net294310), .A(net294364), .ZN(net294362)
         );
  NAND2_X4 U2185 ( .A1(net294393), .A2(net294307), .ZN(n1398) );
  NOR2_X4 U2186 ( .A1(net294365), .A2(net294507), .ZN(net294506) );
  NAND2_X4 U2187 ( .A1(net294510), .A2(net298857), .ZN(net294509) );
  NAND2_X4 U2188 ( .A1(net294247), .A2(net294248), .ZN(net294401) );
  XNOR2_X2 U2189 ( .A(net294401), .B(net294402), .ZN(net294399) );
  NAND3_X2 U2190 ( .A1(net294247), .A2(net294248), .A3(net294249), .ZN(
        net294241) );
  INV_X8 U2192 ( .A(net294636), .ZN(net294447) );
  INV_X8 U2194 ( .A(n1406), .ZN(n1402) );
  OAI21_X4 U2195 ( .B1(n1402), .B2(net294573), .A(net294574), .ZN(net294526)
         );
  OAI21_X4 U2196 ( .B1(n1402), .B2(net294883), .A(net294881), .ZN(net294701)
         );
  OAI211_X4 U2197 ( .C1(n1407), .C2(net294882), .A(n1409), .B(n1408), .ZN(
        n1406) );
  OAI21_X2 U2198 ( .B1(n1403), .B2(net294770), .A(net294787), .ZN(net294784)
         );
  OAI21_X2 U2199 ( .B1(n1403), .B2(net294770), .A(net294879), .ZN(net294698)
         );
  NAND3_X2 U2200 ( .A1(n1405), .A2(net297774), .A3(net299334), .ZN(n1404) );
  INV_X8 U2201 ( .A(net298731), .ZN(n1405) );
  OAI21_X2 U2202 ( .B1(net294889), .B2(net299334), .A(n1405), .ZN(net294888)
         );
  NAND3_X4 U2203 ( .A1(net294994), .A2(n1405), .A3(net294940), .ZN(net294993)
         );
  INV_X4 U2204 ( .A(net294786), .ZN(n1407) );
  NOR2_X4 U2205 ( .A1(net295510), .A2(n1411), .ZN(n1410) );
  AOI21_X4 U2206 ( .B1(n1410), .B2(net298968), .A(net295507), .ZN(net295502)
         );
  NAND2_X2 U2207 ( .A1(n1412), .A2(net295513), .ZN(n1411) );
  INV_X4 U2208 ( .A(net295516), .ZN(net295510) );
  NAND3_X2 U2209 ( .A1(net295506), .A2(net295516), .A3(net295513), .ZN(
        net295741) );
  XNOR2_X2 U2210 ( .A(n1291), .B(net295628), .ZN(net295514) );
  NAND2_X2 U2211 ( .A1(net295736), .A2(net295514), .ZN(net295732) );
  INV_X4 U2212 ( .A(net295514), .ZN(net295738) );
  INV_X4 U2213 ( .A(net295739), .ZN(net295628) );
  NAND2_X2 U2214 ( .A1(n1291), .A2(net295628), .ZN(net295509) );
  NAND2_X2 U2215 ( .A1(a[17]), .A2(net297485), .ZN(net295739) );
  INV_X16 U2216 ( .A(net297484), .ZN(net297485) );
  INV_X4 U2217 ( .A(net297068), .ZN(net297484) );
  OAI21_X4 U2218 ( .B1(net295867), .B2(net295868), .A(net295508), .ZN(
        net295515) );
  XNOR2_X2 U2219 ( .A(net295866), .B(net295515), .ZN(net299089) );
  OAI21_X4 U2220 ( .B1(net295741), .B2(net295515), .A(net295508), .ZN(
        net295737) );
  XNOR2_X2 U2221 ( .A(net295866), .B(net295515), .ZN(net295759) );
  NOR2_X1 U2222 ( .A1(net297276), .A2(net295869), .ZN(net295868) );
  INV_X4 U2223 ( .A(a[15]), .ZN(net295869) );
  INV_X4 U2224 ( .A(net295870), .ZN(net295867) );
  NAND3_X4 U2225 ( .A1(a[15]), .A2(net295867), .A3(net297272), .ZN(net295508)
         );
  NAND2_X1 U2226 ( .A1(a[16]), .A2(net297485), .ZN(net295870) );
  NAND3_X2 U2227 ( .A1(net295745), .A2(net295743), .A3(n1278), .ZN(net295516)
         );
  OAI21_X4 U2228 ( .B1(net294205), .B2(net293933), .A(n1416), .ZN(n1415) );
  NAND2_X1 U2229 ( .A1(n1417), .A2(net294117), .ZN(n1416) );
  INV_X2 U2230 ( .A(net294117), .ZN(net294205) );
  NOR2_X1 U2231 ( .A1(n1413), .A2(n1422), .ZN(n1419) );
  XNOR2_X1 U2232 ( .A(n1152), .B(n1279), .ZN(net299044) );
  XNOR2_X2 U2233 ( .A(n1128), .B(n1279), .ZN(net294102) );
  INV_X4 U2234 ( .A(net296472), .ZN(n1420) );
  MUX2_X2 U2235 ( .A(\set_product_in_sig/z1 [2]), .B(n1420), .S(net297196), 
        .Z(product_out[2]) );
  NAND2_X2 U2236 ( .A1(n1420), .A2(net294053), .ZN(net295587) );
  INV_X8 U2237 ( .A(net294519), .ZN(net294053) );
  NOR2_X4 U2238 ( .A1(net297184), .A2(control[1]), .ZN(net299335) );
  INV_X4 U2239 ( .A(net294101), .ZN(n1413) );
  XNOR2_X2 U2241 ( .A(net294806), .B(net294655), .ZN(net294803) );
  NAND3_X2 U2242 ( .A1(net294653), .A2(net294656), .A3(net294657), .ZN(
        net294837) );
  NAND3_X2 U2243 ( .A1(n4283), .A2(net294837), .A3(n1265), .ZN(net294842) );
  INV_X2 U2244 ( .A(net294837), .ZN(net294909) );
  NAND2_X2 U2245 ( .A1(net294839), .A2(n1282), .ZN(net294658) );
  XNOR2_X2 U2246 ( .A(n1282), .B(net294930), .ZN(net298959) );
  XNOR2_X2 U2247 ( .A(n1282), .B(net294930), .ZN(net294918) );
  INV_X32 U2248 ( .A(n1425), .ZN(net297226) );
  INV_X16 U2249 ( .A(net297230), .ZN(n1425) );
  NAND2_X4 U2250 ( .A1(net297100), .A2(n1424), .ZN(n1423) );
  AOI22_X2 U2251 ( .A1(b[3]), .A2(net297196), .B1(b[11]), .B2(net294515), .ZN(
        n1424) );
  INV_X16 U2252 ( .A(net294048), .ZN(net294515) );
  INV_X32 U2253 ( .A(net297198), .ZN(net297196) );
  NAND2_X2 U2254 ( .A1(control[0]), .A2(net297166), .ZN(net293950) );
  INV_X16 U2255 ( .A(net297640), .ZN(net297166) );
  INV_X32 U2256 ( .A(control[1]), .ZN(net297640) );
  NAND2_X2 U2257 ( .A1(a[3]), .A2(net297640), .ZN(net297086) );
  NAND2_X4 U2258 ( .A1(n1427), .A2(net295172), .ZN(net295170) );
  XNOR2_X2 U2259 ( .A(net295170), .B(net295165), .ZN(net298632) );
  INV_X4 U2260 ( .A(net295170), .ZN(net295018) );
  NAND2_X2 U2261 ( .A1(n1292), .A2(n1428), .ZN(n1427) );
  INV_X4 U2262 ( .A(n1429), .ZN(n1428) );
  XNOR2_X2 U2263 ( .A(n1292), .B(n1428), .ZN(net295282) );
  NAND2_X2 U2264 ( .A1(a[21]), .A2(net297485), .ZN(n1429) );
  NAND2_X4 U2265 ( .A1(net295280), .A2(net295281), .ZN(net295172) );
  NAND2_X2 U2266 ( .A1(net295279), .A2(net295172), .ZN(net295278) );
  INV_X4 U2267 ( .A(net295282), .ZN(net295280) );
  NAND2_X4 U2268 ( .A1(net297061), .A2(n1430), .ZN(net297068) );
  NAND2_X2 U2269 ( .A1(a[9]), .A2(net297068), .ZN(net296432) );
  NAND3_X2 U2270 ( .A1(net297068), .A2(net297515), .A3(n1284), .ZN(net297009)
         );
  INV_X8 U2271 ( .A(n1431), .ZN(n1430) );
  NAND2_X4 U2272 ( .A1(n1430), .A2(net297061), .ZN(net297481) );
  NAND2_X4 U2273 ( .A1(n1430), .A2(net297061), .ZN(net294188) );
  NAND2_X4 U2274 ( .A1(n1430), .A2(net297061), .ZN(net297281) );
  NAND2_X4 U2275 ( .A1(n1432), .A2(n1433), .ZN(n1431) );
  NAND2_X4 U2276 ( .A1(n1434), .A2(b[24]), .ZN(n1433) );
  NOR2_X4 U2277 ( .A1(control[0]), .A2(control[1]), .ZN(n1434) );
  NAND3_X2 U2278 ( .A1(control[0]), .A2(net299325), .A3(b[16]), .ZN(n1432) );
  OAI21_X4 U2279 ( .B1(net295286), .B2(net295287), .A(net295288), .ZN(
        net295281) );
  NAND2_X2 U2280 ( .A1(net295283), .A2(net295282), .ZN(net295279) );
  XNOR2_X2 U2281 ( .A(net295287), .B(net295289), .ZN(net295380) );
  NAND2_X2 U2282 ( .A1(net295385), .A2(net295288), .ZN(net295287) );
  NAND2_X4 U2283 ( .A1(net294820), .A2(net294819), .ZN(net294932) );
  INV_X4 U2284 ( .A(net294932), .ZN(net294931) );
  XNOR2_X2 U2285 ( .A(net294932), .B(net294817), .ZN(net295008) );
  NAND3_X2 U2286 ( .A1(net294820), .A2(net294819), .A3(net294818), .ZN(
        net294815) );
  NAND2_X1 U2287 ( .A1(net295030), .A2(net295031), .ZN(n1436) );
  NAND2_X4 U2288 ( .A1(net295161), .A2(net295162), .ZN(net294819) );
  NAND2_X4 U2289 ( .A1(net295160), .A2(net294819), .ZN(net295029) );
  INV_X4 U2290 ( .A(net298632), .ZN(net295162) );
  INV_X4 U2291 ( .A(net295163), .ZN(net295161) );
  XNOR2_X2 U2292 ( .A(net295159), .B(net295029), .ZN(net295156) );
  NAND2_X4 U2293 ( .A1(net295032), .A2(n1110), .ZN(net295176) );
  OAI21_X4 U2294 ( .B1(net295175), .B2(n1437), .A(net295031), .ZN(net295159)
         );
  NAND2_X4 U2295 ( .A1(net295274), .A2(net295031), .ZN(n1437) );
  XNOR2_X2 U2296 ( .A(net295176), .B(n1437), .ZN(net295271) );
  NOR2_X2 U2297 ( .A1(net295752), .A2(n1439), .ZN(net295742) );
  INV_X4 U2298 ( .A(net295754), .ZN(n1439) );
  INV_X4 U2299 ( .A(net295755), .ZN(net295752) );
  NAND3_X4 U2300 ( .A1(n1346), .A2(net296426), .A3(net296427), .ZN(n1438) );
  NAND2_X4 U2301 ( .A1(net296222), .A2(n1438), .ZN(net296106) );
  NAND2_X4 U2302 ( .A1(n1438), .A2(net295748), .ZN(net295995) );
  NAND3_X4 U2304 ( .A1(n1441), .A2(a[11]), .A3(net297274), .ZN(net295754) );
  INV_X8 U2305 ( .A(net297276), .ZN(net297274) );
  NAND3_X4 U2306 ( .A1(n1440), .A2(a[13]), .A3(net297274), .ZN(net295755) );
  INV_X4 U2307 ( .A(net296099), .ZN(n1440) );
  INV_X4 U2308 ( .A(net296426), .ZN(net296328) );
  INV_X8 U2309 ( .A(net296427), .ZN(net296544) );
  NOR2_X1 U2310 ( .A1(net296529), .A2(n4282), .ZN(net296536) );
  NAND2_X2 U2311 ( .A1(net296098), .A2(net296099), .ZN(net296097) );
  NAND2_X4 U2312 ( .A1(n1442), .A2(net295382), .ZN(net295289) );
  NAND2_X2 U2313 ( .A1(n1443), .A2(n1444), .ZN(n1442) );
  INV_X4 U2314 ( .A(n1445), .ZN(n1444) );
  XNOR2_X2 U2315 ( .A(n1443), .B(n1444), .ZN(net295499) );
  NAND2_X2 U2316 ( .A1(a[19]), .A2(net297485), .ZN(n1445) );
  INV_X4 U2317 ( .A(n1446), .ZN(n1443) );
  NAND2_X2 U2318 ( .A1(a[18]), .A2(net297274), .ZN(n1446) );
  NAND4_X2 U2319 ( .A1(a[17]), .A2(net295382), .A3(net295494), .A4(net297260), 
        .ZN(net295393) );
  INV_X1 U2320 ( .A(net295382), .ZN(net295495) );
  INV_X4 U2321 ( .A(net295499), .ZN(net295501) );
  NAND2_X4 U2322 ( .A1(net299321), .A2(n1447), .ZN(net296426) );
  NAND2_X2 U2323 ( .A1(a[8]), .A2(net297274), .ZN(n1447) );
  INV_X1 U2324 ( .A(net296553), .ZN(net299321) );
  XNOR2_X2 U2325 ( .A(net298482), .B(net296553), .ZN(net299323) );
  NAND2_X4 U2326 ( .A1(net298482), .A2(net296553), .ZN(net296325) );
  XNOR2_X2 U2327 ( .A(net298482), .B(net296553), .ZN(net296554) );
  NAND3_X4 U2328 ( .A1(net296326), .A2(net296325), .A3(net296324), .ZN(
        net296427) );
  NAND2_X4 U2329 ( .A1(net295748), .A2(net296537), .ZN(net296329) );
  NAND2_X2 U2330 ( .A1(net294400), .A2(net299052), .ZN(net294300) );
  NAND2_X4 U2331 ( .A1(net294317), .A2(n1448), .ZN(net294313) );
  INV_X4 U2332 ( .A(net294399), .ZN(net294317) );
  INV_X4 U2333 ( .A(net294400), .ZN(n1448) );
  XNOR2_X2 U2334 ( .A(net294407), .B(n1450), .ZN(n1449) );
  NOR2_X2 U2335 ( .A1(net294253), .A2(net294156), .ZN(n1450) );
  AOI21_X2 U2336 ( .B1(net294405), .B2(net294406), .A(net294253), .ZN(
        net294407) );
  NAND2_X2 U2337 ( .A1(a[22]), .A2(net297204), .ZN(net294400) );
  NOR2_X4 U2338 ( .A1(n1451), .A2(net293988), .ZN(net293986) );
  INV_X4 U2339 ( .A(net294253), .ZN(net294251) );
  NAND2_X4 U2340 ( .A1(net299073), .A2(net294253), .ZN(net294249) );
  NAND2_X2 U2341 ( .A1(net294156), .A2(net294299), .ZN(net294298) );
  INV_X4 U2342 ( .A(net294156), .ZN(net294153) );
  NAND2_X4 U2343 ( .A1(net294405), .A2(net294406), .ZN(net294154) );
  INV_X4 U2345 ( .A(net296539), .ZN(net296540) );
  INV_X1 U2346 ( .A(net295500), .ZN(net295498) );
  NAND2_X2 U2347 ( .A1(net295508), .A2(net295509), .ZN(net295507) );
  NAND3_X2 U2348 ( .A1(net295750), .A2(net295755), .A3(net295757), .ZN(
        net298968) );
  NAND2_X2 U2349 ( .A1(net295498), .A2(net295499), .ZN(net295494) );
  NAND2_X4 U2350 ( .A1(net295622), .A2(net295504), .ZN(net295503) );
  INV_X4 U2351 ( .A(net295019), .ZN(net295165) );
  NAND2_X2 U2352 ( .A1(a[20]), .A2(net297260), .ZN(net295163) );
  INV_X16 U2353 ( .A(net297270), .ZN(net297260) );
  INV_X4 U2354 ( .A(net294175), .ZN(net297270) );
  NOR2_X4 U2355 ( .A1(net297270), .A2(net294006), .ZN(net294004) );
  INV_X8 U2356 ( .A(net297128), .ZN(net294175) );
  OAI21_X4 U2357 ( .B1(net295018), .B2(net295019), .A(net295020), .ZN(
        net295017) );
  OAI21_X4 U2358 ( .B1(net297128), .B2(net293991), .A(net294425), .ZN(
        net294171) );
  NAND2_X4 U2360 ( .A1(net294234), .A2(n1453), .ZN(net294083) );
  NAND2_X2 U2361 ( .A1(a[22]), .A2(net297254), .ZN(n1453) );
  NOR2_X4 U2362 ( .A1(n1456), .A2(net294012), .ZN(net294010) );
  AOI22_X2 U2363 ( .A1(b[31]), .A2(net294051), .B1(b[23]), .B2(net294053), 
        .ZN(n1455) );
  NAND2_X2 U2364 ( .A1(b[7]), .A2(net297196), .ZN(n1454) );
  NAND2_X2 U2365 ( .A1(n1458), .A2(net295624), .ZN(net295622) );
  NAND2_X2 U2366 ( .A1(a[17]), .A2(net297272), .ZN(n1458) );
  NAND3_X2 U2367 ( .A1(n1457), .A2(a[17]), .A3(net297274), .ZN(net295504) );
  INV_X4 U2368 ( .A(net295624), .ZN(n1457) );
  NAND2_X4 U2369 ( .A1(net295626), .A2(net295509), .ZN(net295621) );
  OAI21_X4 U2370 ( .B1(n1459), .B2(n1460), .A(n4279), .ZN(net294437) );
  XNOR2_X2 U2371 ( .A(net294532), .B(net294437), .ZN(net294529) );
  OAI21_X4 U2372 ( .B1(net294536), .B2(net294537), .A(net294538), .ZN(n1460)
         );
  NAND2_X2 U2373 ( .A1(net294645), .A2(n1461), .ZN(net294535) );
  NAND2_X4 U2374 ( .A1(net294538), .A2(net294535), .ZN(net294643) );
  INV_X4 U2375 ( .A(net294646), .ZN(n1461) );
  NAND2_X4 U2376 ( .A1(net294793), .A2(net297593), .ZN(net294537) );
  NAND3_X2 U2377 ( .A1(net294539), .A2(net294540), .A3(net294537), .ZN(
        net294680) );
  NAND2_X4 U2378 ( .A1(net294539), .A2(net294537), .ZN(net294800) );
  NAND3_X4 U2380 ( .A1(net294843), .A2(net297593), .A3(net294795), .ZN(
        net294539) );
  NAND2_X4 U2381 ( .A1(n1462), .A2(net294646), .ZN(net294538) );
  NAND2_X4 U2383 ( .A1(net294803), .A2(net294802), .ZN(net294541) );
  NAND2_X4 U2384 ( .A1(net294680), .A2(net294541), .ZN(net294642) );
  INV_X4 U2385 ( .A(net294804), .ZN(net294802) );
  NAND2_X4 U2386 ( .A1(n4206), .A2(net294804), .ZN(net294540) );
  XNOR2_X2 U2389 ( .A(net294793), .B(net294772), .ZN(net294905) );
  OAI21_X4 U2390 ( .B1(n1265), .B2(net294907), .A(net294842), .ZN(net294793)
         );
  NAND2_X4 U2391 ( .A1(net294795), .A2(net294844), .ZN(net294901) );
  NAND2_X2 U2392 ( .A1(a[22]), .A2(net297216), .ZN(net294530) );
  OAI21_X4 U2393 ( .B1(net294931), .B2(net294817), .A(net294818), .ZN(
        net294841) );
  NAND2_X4 U2394 ( .A1(net294818), .A2(n1463), .ZN(net294817) );
  NAND2_X2 U2395 ( .A1(net294817), .A2(net294818), .ZN(net294816) );
  NAND2_X2 U2396 ( .A1(net295012), .A2(net295013), .ZN(n1463) );
  NAND2_X4 U2397 ( .A1(n1464), .A2(n1465), .ZN(net294818) );
  INV_X4 U2398 ( .A(net295012), .ZN(n1465) );
  INV_X4 U2399 ( .A(net295013), .ZN(n1464) );
  NAND3_X4 U2400 ( .A1(net296540), .A2(a[9]), .A3(net297272), .ZN(net295748)
         );
  NAND2_X2 U2401 ( .A1(a[21]), .A2(net297244), .ZN(net294804) );
  NAND2_X2 U2402 ( .A1(n1467), .A2(net295387), .ZN(net295385) );
  NAND2_X2 U2403 ( .A1(a[19]), .A2(net297272), .ZN(n1467) );
  NAND3_X1 U2404 ( .A1(a[19]), .A2(n1466), .A3(net297274), .ZN(net295288) );
  INV_X4 U2405 ( .A(net295387), .ZN(n1466) );
  XNOR2_X2 U2406 ( .A(net298959), .B(net294840), .ZN(net294657) );
  NAND4_X2 U2407 ( .A1(b[24]), .A2(net297180), .A3(a[5]), .A4(net297640), .ZN(
        net297022) );
  AOI22_X4 U2408 ( .A1(b[27]), .A2(net294051), .B1(b[19]), .B2(net294053), 
        .ZN(net297100) );
  INV_X4 U2409 ( .A(n1469), .ZN(n1468) );
  XNOR2_X2 U2410 ( .A(n1269), .B(n1468), .ZN(net295756) );
  NAND2_X2 U2411 ( .A1(a[15]), .A2(net297485), .ZN(n1469) );
  AOI22_X4 U2412 ( .A1(net294052), .A2(net299241), .B1(net294054), .B2(
        net297196), .ZN(net299240) );
  INV_X4 U2413 ( .A(net297196), .ZN(net297190) );
  NAND2_X2 U2414 ( .A1(n1121), .A2(n1471), .ZN(n1470) );
  NAND2_X4 U2415 ( .A1(net294117), .A2(n1470), .ZN(net293924) );
  NAND2_X2 U2416 ( .A1(\set_product_in_sig/z1 [29]), .A2(net297190), .ZN(n1471) );
  NAND2_X4 U2417 ( .A1(\set_product_in_sig/z1 [29]), .A2(net294220), .ZN(
        net293935) );
  NOR2_X4 U2418 ( .A1(n1472), .A2(n1473), .ZN(net297071) );
  INV_X8 U2419 ( .A(n1474), .ZN(n1473) );
  NOR2_X2 U2420 ( .A1(n1472), .A2(n1473), .ZN(net298916) );
  NAND3_X4 U2421 ( .A1(net297182), .A2(b[9]), .A3(control[1]), .ZN(n1474) );
  INV_X32 U2422 ( .A(control[0]), .ZN(net297182) );
  INV_X4 U2423 ( .A(n1475), .ZN(n1472) );
  NAND3_X4 U2424 ( .A1(control[0]), .A2(control[1]), .A3(b[1]), .ZN(n1475) );
  XNOR2_X2 U2425 ( .A(net294369), .B(net299300), .ZN(net298730) );
  OAI21_X4 U2426 ( .B1(n1477), .B2(n1478), .A(net298969), .ZN(net294372) );
  NAND3_X2 U2427 ( .A1(net294372), .A2(net294371), .A3(net294370), .ZN(
        net299300) );
  INV_X16 U2428 ( .A(net294042), .ZN(net298969) );
  INV_X8 U2429 ( .A(net294314), .ZN(net294042) );
  NAND2_X4 U2430 ( .A1(n1479), .A2(net298969), .ZN(net294371) );
  INV_X2 U2431 ( .A(net294333), .ZN(n1479) );
  NAND2_X2 U2432 ( .A1(n1476), .A2(net298969), .ZN(net294370) );
  NAND2_X4 U2434 ( .A1(net294314), .A2(net294330), .ZN(n1476) );
  NAND4_X4 U2435 ( .A1(net294333), .A2(net294331), .A3(net294332), .A4(
        net294330), .ZN(net294045) );
  XNOR2_X2 U2436 ( .A(net294360), .B(n1476), .ZN(net294359) );
  INV_X4 U2437 ( .A(n1476), .ZN(net294303) );
  NOR2_X2 U2438 ( .A1(n1364), .A2(n1480), .ZN(net295743) );
  NAND3_X1 U2439 ( .A1(net295748), .A2(net295749), .A3(net295750), .ZN(n1480)
         );
  NAND2_X2 U2440 ( .A1(a[11]), .A2(net294188), .ZN(n1483) );
  NAND2_X4 U2441 ( .A1(n1481), .A2(n1482), .ZN(net295745) );
  NAND3_X2 U2442 ( .A1(net298937), .A2(net295745), .A3(net296417), .ZN(
        net296337) );
  INV_X8 U2443 ( .A(net296418), .ZN(n1482) );
  NAND2_X2 U2444 ( .A1(n1481), .A2(n1482), .ZN(net296104) );
  AOI211_X4 U2445 ( .C1(n1481), .C2(n1482), .A(net295995), .B(net295996), .ZN(
        net295982) );
  INV_X8 U2446 ( .A(net296419), .ZN(n1481) );
  NAND2_X2 U2447 ( .A1(net294911), .A2(net294913), .ZN(net294653) );
  INV_X4 U2448 ( .A(net294543), .ZN(n1485) );
  NAND2_X4 U2449 ( .A1(net294543), .A2(n1484), .ZN(net294406) );
  INV_X4 U2450 ( .A(net294544), .ZN(n1484) );
  NAND2_X2 U2451 ( .A1(n1486), .A2(net295020), .ZN(net295019) );
  NAND2_X2 U2452 ( .A1(n1487), .A2(net295168), .ZN(n1486) );
  NAND2_X2 U2453 ( .A1(a[21]), .A2(net297272), .ZN(n1487) );
  INV_X4 U2454 ( .A(net295168), .ZN(net295167) );
  NAND2_X2 U2455 ( .A1(n1489), .A2(net294810), .ZN(n1488) );
  INV_X2 U2456 ( .A(net294809), .ZN(n1489) );
  NAND3_X2 U2457 ( .A1(a[18]), .A2(net295380), .A3(net297260), .ZN(net295030)
         );
  NAND2_X4 U2458 ( .A1(net295275), .A2(n1490), .ZN(net295031) );
  NAND2_X4 U2459 ( .A1(net295291), .A2(n1267), .ZN(net295032) );
  XNOR2_X2 U2460 ( .A(net295291), .B(n1267), .ZN(net298655) );
  NAND2_X2 U2461 ( .A1(n1491), .A2(net295379), .ZN(net295377) );
  INV_X4 U2462 ( .A(net295380), .ZN(net295379) );
  NAND2_X2 U2463 ( .A1(a[18]), .A2(net297260), .ZN(n1491) );
  INV_X2 U2464 ( .A(n2339), .ZN(n1666) );
  INV_X2 U2465 ( .A(net294577), .ZN(net294576) );
  OAI21_X4 U2466 ( .B1(n1846), .B2(n1845), .A(n1847), .ZN(n1492) );
  NOR2_X4 U2467 ( .A1(n2653), .A2(n2652), .ZN(n2524) );
  XNOR2_X2 U2469 ( .A(n2602), .B(n2868), .ZN(n1494) );
  INV_X8 U2470 ( .A(n2764), .ZN(n2868) );
  XNOR2_X2 U2471 ( .A(net294526), .B(n1257), .ZN(n1495) );
  XNOR2_X2 U2472 ( .A(n2016), .B(n2017), .ZN(n1496) );
  OAI211_X4 U2473 ( .C1(n3388), .C2(n3387), .A(n1507), .B(n1543), .ZN(n3389)
         );
  NAND2_X4 U2474 ( .A1(n3500), .A2(n3501), .ZN(n3536) );
  INV_X4 U2475 ( .A(net298392), .ZN(net299331) );
  NAND2_X4 U2476 ( .A1(n2136), .A2(n2230), .ZN(n2316) );
  NAND2_X1 U2477 ( .A1(n2136), .A2(n2230), .ZN(n2292) );
  NAND2_X4 U2480 ( .A1(n1743), .A2(n4249), .ZN(n2186) );
  XNOR2_X2 U2481 ( .A(n3077), .B(n1500), .ZN(n1497) );
  XNOR2_X2 U2482 ( .A(n2873), .B(n1585), .ZN(n1641) );
  XNOR2_X2 U2483 ( .A(n1243), .B(n2981), .ZN(n1498) );
  NAND2_X4 U2484 ( .A1(n3661), .A2(n3662), .ZN(net294840) );
  NAND2_X4 U2485 ( .A1(n3663), .A2(n3662), .ZN(n3758) );
  NAND3_X2 U2486 ( .A1(a[22]), .A2(n3594), .A3(net297260), .ZN(n3662) );
  XNOR2_X2 U2487 ( .A(n3077), .B(n1500), .ZN(n1499) );
  NAND2_X4 U2488 ( .A1(n2830), .A2(n2906), .ZN(n2812) );
  XNOR2_X2 U2489 ( .A(n3995), .B(n1285), .ZN(n1501) );
  OAI21_X2 U2490 ( .B1(net295585), .B2(n3186), .A(n3213), .ZN(n3086) );
  INV_X4 U2492 ( .A(n1799), .ZN(n1510) );
  INV_X1 U2496 ( .A(n4250), .ZN(n2554) );
  INV_X4 U2497 ( .A(n3341), .ZN(n1506) );
  INV_X4 U2498 ( .A(n1506), .ZN(n1507) );
  NAND2_X4 U2499 ( .A1(n3660), .A2(n3759), .ZN(n3760) );
  NOR2_X2 U2500 ( .A1(n1774), .A2(net294995), .ZN(n3504) );
  NAND2_X4 U2501 ( .A1(n3341), .A2(n1543), .ZN(net294995) );
  AOI21_X4 U2502 ( .B1(n3750), .B2(n1281), .A(n1509), .ZN(n1508) );
  INV_X4 U2503 ( .A(n3750), .ZN(n3806) );
  NAND2_X4 U2504 ( .A1(n4067), .A2(net299044), .ZN(n4176) );
  NAND2_X2 U2505 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  NAND2_X4 U2507 ( .A1(n3822), .A2(n3821), .ZN(n3939) );
  OAI21_X4 U2509 ( .B1(n2829), .B2(n2828), .A(n2814), .ZN(n2894) );
  INV_X4 U2510 ( .A(n2826), .ZN(n2829) );
  NAND2_X4 U2511 ( .A1(net294303), .A2(n3935), .ZN(n3936) );
  OAI21_X2 U2512 ( .B1(net294305), .B2(n3934), .A(n1344), .ZN(n3935) );
  INV_X4 U2514 ( .A(n1513), .ZN(n1514) );
  INV_X1 U2515 ( .A(n4292), .ZN(n1515) );
  INV_X2 U2516 ( .A(n1515), .ZN(n1516) );
  NAND2_X4 U2517 ( .A1(n3853), .A2(n4061), .ZN(n3715) );
  AOI21_X2 U2518 ( .B1(n3673), .B2(net294779), .A(n1774), .ZN(n3505) );
  NAND2_X2 U2520 ( .A1(n4045), .A2(n1512), .ZN(n4046) );
  INV_X4 U2521 ( .A(n2005), .ZN(n2007) );
  NAND3_X2 U2522 ( .A1(a[4]), .A2(n2005), .A3(net297260), .ZN(n2234) );
  NAND2_X4 U2523 ( .A1(n3902), .A2(net294394), .ZN(n1517) );
  XNOR2_X2 U2524 ( .A(n3678), .B(n3679), .ZN(n1519) );
  XNOR2_X1 U2525 ( .A(n2722), .B(n4253), .ZN(n1520) );
  NAND2_X2 U2526 ( .A1(n3382), .A2(n1108), .ZN(n3170) );
  INV_X4 U2527 ( .A(n2835), .ZN(n2706) );
  OAI22_X2 U2528 ( .A1(n3112), .A2(n3111), .B1(n3110), .B2(n3109), .ZN(n1521)
         );
  NOR2_X2 U2529 ( .A1(n3108), .A2(n3107), .ZN(n3109) );
  INV_X1 U2530 ( .A(n3118), .ZN(n2983) );
  XNOR2_X1 U2531 ( .A(n1242), .B(n3394), .ZN(n1522) );
  INV_X1 U2532 ( .A(net299073), .ZN(net294252) );
  XNOR2_X2 U2533 ( .A(n3770), .B(n3769), .ZN(n1523) );
  AOI22_X4 U2534 ( .A1(n3741), .A2(n3740), .B1(n3739), .B2(n3905), .ZN(n3770)
         );
  INV_X1 U2535 ( .A(n2278), .ZN(n2281) );
  OAI22_X2 U2536 ( .A1(n2697), .A2(n2757), .B1(n2757), .B2(n2766), .ZN(n2698)
         );
  INV_X2 U2538 ( .A(n3556), .ZN(n3550) );
  OAI221_X2 U2539 ( .B1(net294092), .B2(net294093), .C1(n4072), .C2(n4071), 
        .A(n4070), .ZN(n1525) );
  NAND2_X2 U2540 ( .A1(n2242), .A2(n1607), .ZN(n2483) );
  NAND2_X4 U2541 ( .A1(n3347), .A2(n3346), .ZN(n3560) );
  NAND2_X4 U2542 ( .A1(n4104), .A2(n4075), .ZN(n4076) );
  INV_X8 U2543 ( .A(n1526), .ZN(n1527) );
  INV_X4 U2544 ( .A(net296781), .ZN(net299191) );
  NAND2_X4 U2545 ( .A1(n1796), .A2(net299191), .ZN(n2220) );
  INV_X2 U2546 ( .A(n2114), .ZN(n1529) );
  NAND2_X4 U2547 ( .A1(n3745), .A2(n3744), .ZN(n3678) );
  AOI21_X2 U2548 ( .B1(n2297), .B2(n2292), .A(n2296), .ZN(n2294) );
  OAI21_X4 U2549 ( .B1(n3384), .B2(n3383), .A(n1595), .ZN(n1530) );
  NAND3_X2 U2550 ( .A1(n3715), .A2(n3870), .A3(n1623), .ZN(n1531) );
  NAND2_X2 U2551 ( .A1(net294040), .A2(n4085), .ZN(n4087) );
  INV_X4 U2552 ( .A(net297009), .ZN(net297615) );
  NAND2_X4 U2553 ( .A1(n2720), .A2(n2721), .ZN(n2722) );
  NAND2_X4 U2554 ( .A1(n2892), .A2(n2891), .ZN(n1532) );
  NAND2_X2 U2555 ( .A1(n2892), .A2(n2891), .ZN(n3368) );
  NAND2_X4 U2556 ( .A1(n1150), .A2(n3073), .ZN(n3106) );
  INV_X8 U2557 ( .A(n3906), .ZN(n3902) );
  INV_X2 U2558 ( .A(n3393), .ZN(n1534) );
  INV_X8 U2559 ( .A(n1534), .ZN(n1535) );
  NAND2_X4 U2560 ( .A1(n2867), .A2(n2866), .ZN(n2766) );
  NAND2_X1 U2561 ( .A1(n1687), .A2(n1332), .ZN(n1536) );
  INV_X1 U2562 ( .A(n1778), .ZN(n1537) );
  NOR2_X2 U2563 ( .A1(n2217), .A2(n2216), .ZN(n2219) );
  XNOR2_X2 U2564 ( .A(n1538), .B(n3648), .ZN(n3594) );
  XNOR2_X2 U2565 ( .A(n3542), .B(n1161), .ZN(n3700) );
  NOR2_X4 U2566 ( .A1(n1636), .A2(n2980), .ZN(n1551) );
  NAND2_X4 U2567 ( .A1(n3790), .A2(n4054), .ZN(n4060) );
  NAND2_X4 U2568 ( .A1(n1560), .A2(n2889), .ZN(n3099) );
  XOR2_X1 U2569 ( .A(n4134), .B(n4010), .Z(n1541) );
  INV_X8 U2570 ( .A(n3703), .ZN(n3707) );
  INV_X8 U2571 ( .A(n3502), .ZN(n3311) );
  INV_X2 U2572 ( .A(n2751), .ZN(n1775) );
  CLKBUF_X3 U2573 ( .A(n2730), .Z(n1545) );
  NOR2_X4 U2574 ( .A1(n2742), .A2(n2741), .ZN(n2745) );
  INV_X4 U2575 ( .A(n2798), .ZN(n1546) );
  NAND2_X2 U2576 ( .A1(n2934), .A2(n2933), .ZN(n2941) );
  NAND2_X4 U2577 ( .A1(n2102), .A2(n2301), .ZN(n2103) );
  INV_X4 U2578 ( .A(net294175), .ZN(net297268) );
  INV_X4 U2579 ( .A(net297268), .ZN(net297262) );
  NAND2_X2 U2580 ( .A1(n1924), .A2(n1586), .ZN(n1870) );
  XNOR2_X2 U2581 ( .A(net294800), .B(net294801), .ZN(n1547) );
  XNOR2_X2 U2582 ( .A(net294154), .B(net294153), .ZN(net299073) );
  INV_X1 U2583 ( .A(n1930), .ZN(n2067) );
  INV_X2 U2584 ( .A(n2323), .ZN(n2071) );
  OAI21_X4 U2585 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n1548) );
  OAI21_X2 U2586 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(net299066) );
  INV_X4 U2587 ( .A(n1549), .ZN(n1550) );
  INV_X8 U2588 ( .A(n1551), .ZN(n3257) );
  INV_X2 U2589 ( .A(n2980), .ZN(n3022) );
  NAND2_X4 U2590 ( .A1(a[13]), .A2(net297244), .ZN(n2980) );
  INV_X2 U2591 ( .A(n1950), .ZN(n1552) );
  INV_X2 U2592 ( .A(n1553), .ZN(n1950) );
  NOR2_X4 U2593 ( .A1(n1644), .A2(n1259), .ZN(n2909) );
  AOI211_X2 U2594 ( .C1(n2418), .C2(n1168), .A(net296672), .B(n2211), .ZN(
        n2217) );
  NOR2_X2 U2595 ( .A1(n3433), .A2(n4043), .ZN(n3428) );
  INV_X1 U2596 ( .A(net294326), .ZN(net299046) );
  INV_X2 U2597 ( .A(net299046), .ZN(net299047) );
  NAND2_X2 U2598 ( .A1(n2855), .A2(n2949), .ZN(n2835) );
  NOR2_X4 U2599 ( .A1(n1852), .A2(n1554), .ZN(n1553) );
  OAI21_X4 U2600 ( .B1(n3926), .B2(net297278), .A(n3925), .ZN(n3995) );
  INV_X1 U2601 ( .A(n3637), .ZN(n3638) );
  BUF_X4 U2602 ( .A(n2324), .Z(n1556) );
  OAI21_X1 U2603 ( .B1(n3221), .B2(net297278), .A(n3220), .ZN(n3353) );
  AOI22_X1 U2604 ( .A1(n3353), .A2(n3352), .B1(n3448), .B2(n3287), .ZN(n3288)
         );
  INV_X2 U2605 ( .A(n3353), .ZN(n3448) );
  NAND2_X4 U2606 ( .A1(n2451), .A2(n2625), .ZN(n2452) );
  OAI21_X4 U2607 ( .B1(n3101), .B2(n3100), .A(n3099), .ZN(n3102) );
  NAND2_X2 U2608 ( .A1(n3100), .A2(n3101), .ZN(n3018) );
  XNOR2_X2 U2609 ( .A(n4063), .B(n3623), .ZN(n1557) );
  NAND2_X2 U2610 ( .A1(n1524), .A2(n1155), .ZN(n1692) );
  XNOR2_X2 U2611 ( .A(n2888), .B(n2887), .ZN(n1560) );
  NAND2_X2 U2612 ( .A1(n3127), .A2(n3116), .ZN(n2888) );
  INV_X2 U2613 ( .A(n2065), .ZN(n2106) );
  INV_X2 U2614 ( .A(net298730), .ZN(net299020) );
  NAND2_X2 U2615 ( .A1(n4034), .A2(n4274), .ZN(n4035) );
  NAND2_X1 U2616 ( .A1(a[23]), .A2(net297272), .ZN(n3585) );
  NAND3_X2 U2617 ( .A1(a[21]), .A2(net295167), .A3(net297272), .ZN(net295020)
         );
  NAND3_X2 U2618 ( .A1(n3587), .A2(a[23]), .A3(net297272), .ZN(n3646) );
  NAND3_X2 U2619 ( .A1(n2734), .A2(n2718), .A3(n1545), .ZN(n2721) );
  NOR2_X1 U2620 ( .A1(net294308), .A2(net294309), .ZN(n3934) );
  XNOR2_X2 U2621 ( .A(n3544), .B(n1563), .ZN(n1562) );
  INV_X8 U2622 ( .A(n3725), .ZN(n1763) );
  INV_X8 U2623 ( .A(net296932), .ZN(net296771) );
  XNOR2_X2 U2624 ( .A(n1565), .B(n1566), .ZN(n3628) );
  AND3_X4 U2625 ( .A1(n3563), .A2(n3562), .A3(n3564), .ZN(n1565) );
  AND3_X2 U2626 ( .A1(n3565), .A2(n1593), .A3(n3564), .ZN(n1566) );
  INV_X1 U2627 ( .A(n3911), .ZN(n3775) );
  NAND2_X2 U2628 ( .A1(n2084), .A2(n1634), .ZN(n2090) );
  NAND3_X4 U2629 ( .A1(n1244), .A2(n1798), .A3(n3425), .ZN(n3300) );
  INV_X8 U2630 ( .A(n1981), .ZN(n2111) );
  INV_X2 U2631 ( .A(n2116), .ZN(n1568) );
  INV_X4 U2632 ( .A(n1568), .ZN(n1569) );
  INV_X2 U2633 ( .A(net294299), .ZN(net294155) );
  NAND2_X4 U2634 ( .A1(n2957), .A2(n1132), .ZN(n3054) );
  AND2_X2 U2637 ( .A1(n3835), .A2(n3774), .ZN(n1571) );
  AND2_X2 U2638 ( .A1(n3121), .A2(n1192), .ZN(n3115) );
  NAND2_X4 U2639 ( .A1(n2723), .A2(n2724), .ZN(n2727) );
  INV_X4 U2640 ( .A(net298912), .ZN(net294016) );
  NAND2_X4 U2641 ( .A1(n2885), .A2(n2886), .ZN(n2887) );
  XNOR2_X2 U2642 ( .A(n1120), .B(n3106), .ZN(n1575) );
  NAND2_X1 U2643 ( .A1(n1828), .A2(n1849), .ZN(net296472) );
  INV_X4 U2644 ( .A(n3603), .ZN(n3605) );
  XNOR2_X2 U2645 ( .A(n2973), .B(n2972), .ZN(n1576) );
  NAND3_X2 U2646 ( .A1(n2072), .A2(n2233), .A3(n2232), .ZN(n2235) );
  NAND2_X1 U2647 ( .A1(n2206), .A2(n1796), .ZN(n2233) );
  NAND2_X4 U2648 ( .A1(n3967), .A2(n3999), .ZN(n4000) );
  NAND2_X2 U2650 ( .A1(n2336), .A2(n2489), .ZN(n2415) );
  OAI21_X4 U2651 ( .B1(n1212), .B2(n1936), .A(n1941), .ZN(n1578) );
  NAND2_X4 U2652 ( .A1(a[3]), .A2(net294175), .ZN(n1941) );
  XNOR2_X2 U2653 ( .A(n3891), .B(n3890), .ZN(n1579) );
  NAND3_X2 U2654 ( .A1(net294787), .A2(net294786), .A3(net294788), .ZN(n3668)
         );
  XOR2_X2 U2655 ( .A(n3964), .B(n3963), .Z(n1580) );
  XNOR2_X2 U2656 ( .A(n4134), .B(n4010), .ZN(n4115) );
  NAND2_X4 U2657 ( .A1(n4121), .A2(n4006), .ZN(n4134) );
  INV_X2 U2658 ( .A(n4010), .ZN(n4135) );
  NAND2_X4 U2659 ( .A1(n4009), .A2(n4008), .ZN(n4010) );
  NAND2_X4 U2660 ( .A1(n2634), .A2(n2730), .ZN(n2545) );
  INV_X1 U2661 ( .A(n1696), .ZN(n1581) );
  XNOR2_X2 U2662 ( .A(n3539), .B(n3606), .ZN(n1583) );
  XNOR2_X2 U2663 ( .A(net294918), .B(net294840), .ZN(n1584) );
  NOR2_X2 U2664 ( .A1(n3912), .A2(net294309), .ZN(n3688) );
  INV_X1 U2665 ( .A(net295991), .ZN(net298937) );
  NAND2_X2 U2666 ( .A1(n3543), .A2(n1365), .ZN(n3633) );
  INV_X2 U2667 ( .A(n1920), .ZN(n1921) );
  INV_X8 U2668 ( .A(n3950), .ZN(n3953) );
  NAND2_X4 U2669 ( .A1(n3426), .A2(n3300), .ZN(n4045) );
  XNOR2_X2 U2671 ( .A(n3896), .B(n3895), .ZN(n1610) );
  INV_X1 U2672 ( .A(net295008), .ZN(net295010) );
  INV_X4 U2674 ( .A(n2890), .ZN(n2891) );
  INV_X2 U2675 ( .A(n2260), .ZN(n2258) );
  OAI21_X4 U2676 ( .B1(n3696), .B2(n3695), .A(n3694), .ZN(n3711) );
  NAND4_X4 U2677 ( .A1(b[0]), .A2(net297166), .A3(a[3]), .A4(control[0]), .ZN(
        n1586) );
  NAND2_X4 U2678 ( .A1(net297515), .A2(a[3]), .ZN(n1650) );
  INV_X1 U2679 ( .A(net296910), .ZN(net298912) );
  INV_X4 U2680 ( .A(net297481), .ZN(net296910) );
  NAND3_X2 U2681 ( .A1(n3517), .A2(n3400), .A3(n3401), .ZN(n3318) );
  XNOR2_X2 U2683 ( .A(net295621), .B(net298907), .ZN(n1617) );
  NAND2_X4 U2684 ( .A1(n2610), .A2(n2609), .ZN(n2612) );
  NOR2_X2 U2685 ( .A1(n2297), .A2(n2298), .ZN(n2299) );
  XNOR2_X2 U2686 ( .A(n1587), .B(n3953), .ZN(net294426) );
  XNOR2_X2 U2687 ( .A(n3414), .B(n3413), .ZN(n1588) );
  XNOR2_X2 U2688 ( .A(n2876), .B(n2875), .ZN(n1589) );
  NAND2_X4 U2689 ( .A1(n2859), .A2(n2860), .ZN(n2876) );
  NAND2_X4 U2691 ( .A1(n1299), .A2(n2810), .ZN(n2913) );
  NAND2_X4 U2692 ( .A1(n1352), .A2(n3484), .ZN(n3565) );
  NAND2_X4 U2693 ( .A1(n2906), .A2(n2902), .ZN(n2713) );
  NAND2_X4 U2694 ( .A1(n1644), .A2(n1259), .ZN(n2906) );
  XNOR2_X2 U2695 ( .A(n2682), .B(n2774), .ZN(n1591) );
  XNOR2_X1 U2696 ( .A(n3156), .B(n3155), .ZN(n1592) );
  NAND3_X1 U2697 ( .A1(n1857), .A2(n1858), .A3(n1859), .ZN(n1848) );
  NAND2_X2 U2698 ( .A1(n1492), .A2(n1848), .ZN(n1850) );
  NAND2_X4 U2699 ( .A1(n2901), .A2(n2900), .ZN(n3369) );
  NAND2_X2 U2700 ( .A1(n2719), .A2(n2718), .ZN(n2720) );
  NAND2_X4 U2701 ( .A1(n3418), .A2(n3419), .ZN(n1593) );
  NAND2_X4 U2702 ( .A1(n2468), .A2(n2467), .ZN(n2442) );
  NOR2_X4 U2703 ( .A1(n2618), .A2(n1283), .ZN(n1594) );
  INV_X8 U2704 ( .A(n1594), .ZN(n2917) );
  AND2_X4 U2705 ( .A1(n3623), .A2(n1611), .ZN(n1596) );
  INV_X1 U2706 ( .A(n4063), .ZN(n1611) );
  INV_X8 U2707 ( .A(n3829), .ZN(n1597) );
  NAND3_X2 U2709 ( .A1(n3438), .A2(n3437), .A3(n3436), .ZN(n1598) );
  XNOR2_X2 U2710 ( .A(n2381), .B(n2462), .ZN(net298860) );
  XNOR2_X2 U2711 ( .A(n1890), .B(n1552), .ZN(n1599) );
  XNOR2_X2 U2712 ( .A(n2894), .B(n1621), .ZN(n1600) );
  AOI21_X2 U2713 ( .B1(n2669), .B2(n2797), .A(n2563), .ZN(n2514) );
  NAND2_X4 U2714 ( .A1(n3573), .A2(n3540), .ZN(n3574) );
  NAND3_X2 U2715 ( .A1(n2938), .A2(n1133), .A3(n2939), .ZN(n2940) );
  NAND2_X2 U2716 ( .A1(n3444), .A2(n1598), .ZN(n4058) );
  INV_X4 U2717 ( .A(n2479), .ZN(n1601) );
  NAND3_X1 U2718 ( .A1(net294100), .A2(n4175), .A3(net293935), .ZN(n4071) );
  NAND2_X2 U2719 ( .A1(n1593), .A2(n3734), .ZN(n3575) );
  XNOR2_X2 U2720 ( .A(n3602), .B(net294901), .ZN(n3603) );
  INV_X4 U2721 ( .A(n3582), .ZN(n1603) );
  INV_X8 U2722 ( .A(n1603), .ZN(n1604) );
  INV_X1 U2723 ( .A(n4248), .ZN(n1605) );
  INV_X2 U2724 ( .A(net298389), .ZN(net298829) );
  OAI21_X4 U2725 ( .B1(n2848), .B2(n1215), .A(n3031), .ZN(n3033) );
  NAND3_X2 U2726 ( .A1(net296222), .A2(n2589), .A3(n1637), .ZN(n2596) );
  INV_X2 U2729 ( .A(n2607), .ZN(n2608) );
  XNOR2_X2 U2730 ( .A(n2587), .B(n2588), .ZN(n2771) );
  INV_X4 U2731 ( .A(n3624), .ZN(n1608) );
  INV_X4 U2732 ( .A(n3788), .ZN(n3624) );
  XNOR2_X2 U2733 ( .A(net296424), .B(n1483), .ZN(net296221) );
  NAND3_X2 U2735 ( .A1(n1621), .A2(n4254), .A3(n3013), .ZN(n2996) );
  AOI21_X2 U2736 ( .B1(n2552), .B2(n2641), .A(n1272), .ZN(n2553) );
  INV_X2 U2737 ( .A(n2641), .ZN(n2466) );
  INV_X4 U2738 ( .A(n1575), .ZN(n2985) );
  NAND2_X4 U2740 ( .A1(n4197), .A2(n1260), .ZN(n3341) );
  INV_X8 U2741 ( .A(n3905), .ZN(n3913) );
  XNOR2_X2 U2742 ( .A(n2637), .B(n2647), .ZN(n1612) );
  XNOR2_X2 U2743 ( .A(n4076), .B(n1261), .ZN(n1613) );
  NOR2_X2 U2744 ( .A1(n3430), .A2(n3446), .ZN(n3431) );
  AOI21_X1 U2745 ( .B1(net294053), .B2(n4051), .A(n4050), .ZN(n4052) );
  NOR2_X4 U2746 ( .A1(n3726), .A2(n3680), .ZN(n1614) );
  INV_X8 U2747 ( .A(n1614), .ZN(n3905) );
  INV_X2 U2748 ( .A(n3680), .ZN(n3727) );
  NAND2_X4 U2749 ( .A1(a[19]), .A2(net297204), .ZN(n3680) );
  NAND2_X4 U2750 ( .A1(n1280), .A2(n3083), .ZN(n1615) );
  NAND2_X4 U2752 ( .A1(n2995), .A2(n3010), .ZN(n3280) );
  INV_X4 U2753 ( .A(n3012), .ZN(n1620) );
  INV_X4 U2754 ( .A(n2624), .ZN(n1622) );
  NAND2_X4 U2756 ( .A1(n3489), .A2(n3490), .ZN(n3307) );
  NAND3_X2 U2757 ( .A1(n3488), .A2(n3489), .A3(n3490), .ZN(n3491) );
  INV_X1 U2758 ( .A(net294087), .ZN(net294367) );
  AOI21_X4 U2759 ( .B1(n3781), .B2(n1656), .A(net294102), .ZN(n3782) );
  INV_X4 U2760 ( .A(n2760), .ZN(n1624) );
  INV_X8 U2761 ( .A(n1624), .ZN(n1625) );
  NAND2_X4 U2764 ( .A1(net296529), .A2(n1345), .ZN(n2407) );
  NAND2_X1 U2765 ( .A1(a[7]), .A2(net297230), .ZN(n2337) );
  XNOR2_X2 U2766 ( .A(n1225), .B(n1884), .ZN(n1627) );
  XNOR2_X2 U2767 ( .A(n3270), .B(n3577), .ZN(n1628) );
  NAND2_X4 U2768 ( .A1(n1156), .A2(n2827), .ZN(n2814) );
  NAND2_X4 U2769 ( .A1(n4201), .A2(net296524), .ZN(n1629) );
  INV_X4 U2770 ( .A(n1583), .ZN(n3682) );
  OAI21_X2 U2772 ( .B1(n3313), .B2(n3076), .A(n3386), .ZN(n3314) );
  INV_X4 U2773 ( .A(n1931), .ZN(n1817) );
  INV_X4 U2774 ( .A(n2236), .ZN(n2335) );
  XOR2_X2 U2775 ( .A(n2507), .B(n2506), .Z(n1631) );
  XNOR2_X2 U2776 ( .A(n2073), .B(n2076), .ZN(n1632) );
  NOR2_X4 U2777 ( .A1(n3416), .A2(n3415), .ZN(net298731) );
  INV_X2 U2778 ( .A(n3415), .ZN(n3501) );
  NAND3_X2 U2780 ( .A1(n2992), .A2(n2814), .A3(n1148), .ZN(n3013) );
  NAND3_X2 U2781 ( .A1(n2116), .A2(n2115), .A3(n2114), .ZN(n2117) );
  XNOR2_X2 U2782 ( .A(net294642), .B(net294643), .ZN(net298716) );
  XNOR2_X2 U2783 ( .A(n2979), .B(n1239), .ZN(n1636) );
  XNOR2_X2 U2784 ( .A(n2678), .B(n2677), .ZN(n1637) );
  XNOR2_X2 U2785 ( .A(n1639), .B(n3817), .ZN(n3764) );
  AND2_X4 U2786 ( .A1(n3814), .A2(n3816), .ZN(n1639) );
  NAND2_X2 U2787 ( .A1(n2467), .A2(n2405), .ZN(n2347) );
  INV_X1 U2788 ( .A(net295176), .ZN(net295175) );
  XNOR2_X2 U2789 ( .A(n2631), .B(n2632), .ZN(n1640) );
  BUF_X2 U2790 ( .A(n2118), .Z(n1643) );
  XNOR2_X2 U2791 ( .A(n2712), .B(n2711), .ZN(n1644) );
  NAND2_X4 U2792 ( .A1(net294087), .A2(net294088), .ZN(net294326) );
  NAND2_X2 U2793 ( .A1(n4089), .A2(n4040), .ZN(n1648) );
  NAND2_X2 U2794 ( .A1(n1646), .A2(n1647), .ZN(n1649) );
  NAND2_X4 U2795 ( .A1(n1648), .A2(n1649), .ZN(n4090) );
  INV_X4 U2796 ( .A(n4041), .ZN(n1646) );
  INV_X4 U2797 ( .A(n4040), .ZN(n1647) );
  NAND2_X4 U2798 ( .A1(n3766), .A2(n4275), .ZN(n3773) );
  NAND2_X4 U2799 ( .A1(n2194), .A2(n2107), .ZN(n2109) );
  INV_X4 U2800 ( .A(n3671), .ZN(n3677) );
  NAND2_X1 U2801 ( .A1(n3066), .A2(n3137), .ZN(n1654) );
  NAND2_X4 U2802 ( .A1(n1654), .A2(n1655), .ZN(n3259) );
  INV_X2 U2803 ( .A(n3066), .ZN(n1652) );
  NAND2_X1 U2804 ( .A1(n4107), .A2(n4207), .ZN(n4149) );
  NAND3_X2 U2806 ( .A1(n2488), .A2(n2487), .A3(n2486), .ZN(n2507) );
  NAND2_X4 U2807 ( .A1(n3371), .A2(n3103), .ZN(n3227) );
  NAND2_X4 U2808 ( .A1(net294188), .A2(a[8]), .ZN(n2120) );
  INV_X8 U2809 ( .A(n2120), .ZN(n2202) );
  XNOR2_X2 U2810 ( .A(n1980), .B(n2305), .ZN(n2024) );
  INV_X4 U2811 ( .A(n1980), .ZN(n2306) );
  INV_X4 U2812 ( .A(net298655), .ZN(net295372) );
  NAND3_X2 U2815 ( .A1(net294786), .A2(net294788), .A3(net294879), .ZN(n3732)
         );
  NAND3_X2 U2816 ( .A1(n3595), .A2(net294913), .A3(n3596), .ZN(net294656) );
  NAND2_X4 U2817 ( .A1(n3121), .A2(n3122), .ZN(n3123) );
  NAND2_X4 U2818 ( .A1(n2878), .A2(n2877), .ZN(n2939) );
  INV_X4 U2820 ( .A(n1157), .ZN(n2967) );
  AOI21_X2 U2821 ( .B1(n2757), .B2(n1691), .A(n2862), .ZN(n2769) );
  XNOR2_X2 U2822 ( .A(n4108), .B(n4025), .ZN(n1657) );
  NAND2_X4 U2823 ( .A1(n3803), .A2(n3802), .ZN(n3938) );
  NOR2_X4 U2824 ( .A1(n1597), .A2(n1769), .ZN(n1768) );
  AOI21_X4 U2825 ( .B1(n1630), .B2(n1713), .A(n1880), .ZN(n1882) );
  NOR2_X2 U2826 ( .A1(n1871), .A2(n1870), .ZN(n1872) );
  NAND2_X4 U2827 ( .A1(n3801), .A2(n3800), .ZN(net294450) );
  INV_X1 U2828 ( .A(n1557), .ZN(n4056) );
  AOI21_X2 U2829 ( .B1(n3619), .B2(n3692), .A(n1557), .ZN(n3620) );
  NAND2_X2 U2830 ( .A1(n2250), .A2(n2251), .ZN(n2404) );
  NAND2_X4 U2831 ( .A1(n3257), .A2(n3327), .ZN(n1662) );
  OAI21_X4 U2832 ( .B1(net297196), .B2(net294485), .A(n1548), .ZN(n4069) );
  NAND3_X2 U2833 ( .A1(n3827), .A2(n3842), .A3(n3843), .ZN(net294485) );
  INV_X2 U2834 ( .A(n2279), .ZN(n2280) );
  OAI21_X2 U2835 ( .B1(n1676), .B2(n1951), .A(n1492), .ZN(n1886) );
  NAND2_X2 U2836 ( .A1(n3312), .A2(n3231), .ZN(n3385) );
  INV_X4 U2837 ( .A(net296842), .ZN(net296788) );
  NAND2_X4 U2838 ( .A1(n3331), .A2(n1663), .ZN(n3069) );
  INV_X4 U2839 ( .A(n1662), .ZN(n1663) );
  AND2_X4 U2840 ( .A1(n1692), .A2(n2699), .ZN(n1664) );
  NAND2_X2 U2841 ( .A1(n2791), .A2(n2949), .ZN(n2792) );
  NAND2_X1 U2842 ( .A1(n2340), .A2(n2339), .ZN(n1667) );
  NAND2_X2 U2843 ( .A1(n1666), .A2(n1665), .ZN(n1668) );
  NAND2_X2 U2844 ( .A1(n1667), .A2(n1668), .ZN(n2341) );
  INV_X4 U2845 ( .A(n2340), .ZN(n1665) );
  INV_X2 U2846 ( .A(n2585), .ZN(n2203) );
  NAND2_X2 U2848 ( .A1(n3278), .A2(n1616), .ZN(n3084) );
  INV_X4 U2849 ( .A(n3142), .ZN(n3145) );
  INV_X4 U2850 ( .A(n2100), .ZN(n1959) );
  NAND2_X1 U2851 ( .A1(n2007), .A2(n2006), .ZN(n1669) );
  NOR2_X1 U2852 ( .A1(net294016), .A2(n1810), .ZN(n1808) );
  INV_X1 U2853 ( .A(n2317), .ZN(n1670) );
  OAI21_X2 U2854 ( .B1(n1989), .B2(n1988), .A(n2118), .ZN(n1990) );
  NAND2_X1 U2855 ( .A1(n4005), .A2(n4004), .ZN(n4006) );
  INV_X2 U2856 ( .A(n4005), .ZN(n4002) );
  INV_X4 U2858 ( .A(n2578), .ZN(n2581) );
  NAND2_X4 U2859 ( .A1(n3406), .A2(net295158), .ZN(n3520) );
  INV_X2 U2860 ( .A(net295156), .ZN(net295158) );
  NAND2_X4 U2861 ( .A1(n3275), .A2(n3464), .ZN(n3425) );
  INV_X8 U2862 ( .A(n2759), .ZN(n2493) );
  NAND2_X2 U2863 ( .A1(n3673), .A2(net294779), .ZN(n3675) );
  NAND2_X2 U2864 ( .A1(n1331), .A2(n1525), .ZN(n1761) );
  INV_X4 U2865 ( .A(n2617), .ZN(n1672) );
  NOR2_X4 U2866 ( .A1(n1827), .A2(n1826), .ZN(n1676) );
  INV_X4 U2867 ( .A(n3853), .ZN(n1677) );
  NAND2_X2 U2868 ( .A1(n2706), .A2(n2705), .ZN(n1681) );
  NAND2_X4 U2869 ( .A1(n1679), .A2(n1680), .ZN(n1682) );
  NAND2_X4 U2870 ( .A1(n1681), .A2(n1682), .ZN(n2799) );
  INV_X4 U2871 ( .A(n2706), .ZN(n1679) );
  INV_X4 U2872 ( .A(n2705), .ZN(n1680) );
  INV_X4 U2873 ( .A(n2842), .ZN(n2843) );
  INV_X4 U2874 ( .A(net296326), .ZN(net296781) );
  INV_X8 U2875 ( .A(n2108), .ZN(n2110) );
  NAND2_X1 U2876 ( .A1(n3478), .A2(n1240), .ZN(n3481) );
  INV_X1 U2877 ( .A(n1637), .ZN(n2590) );
  INV_X2 U2878 ( .A(n3929), .ZN(n1708) );
  AOI21_X2 U2879 ( .B1(n3919), .B2(net298149), .A(n3918), .ZN(n3928) );
  OAI21_X2 U2880 ( .B1(n3917), .B2(net294353), .A(net297196), .ZN(n3918) );
  NAND2_X2 U2881 ( .A1(a[2]), .A2(net297281), .ZN(n1811) );
  NAND2_X2 U2882 ( .A1(n2944), .A2(n2942), .ZN(n1685) );
  NAND2_X4 U2883 ( .A1(n1684), .A2(n2865), .ZN(n1686) );
  NAND2_X4 U2884 ( .A1(n1685), .A2(n1686), .ZN(n2785) );
  INV_X8 U2885 ( .A(n2944), .ZN(n1684) );
  OAI21_X2 U2886 ( .B1(n2763), .B2(n2762), .A(n2761), .ZN(n2767) );
  NAND2_X4 U2887 ( .A1(n3223), .A2(n3224), .ZN(n1687) );
  NAND2_X2 U2888 ( .A1(n2342), .A2(n1537), .ZN(n1779) );
  OAI21_X4 U2889 ( .B1(n1306), .B2(n3793), .A(n3792), .ZN(n3794) );
  NOR2_X4 U2890 ( .A1(n1640), .A2(n1262), .ZN(n1688) );
  NAND2_X2 U2891 ( .A1(n3916), .A2(n3874), .ZN(n3839) );
  NOR3_X2 U2892 ( .A1(n2652), .A2(n2653), .A3(n2654), .ZN(n2658) );
  NAND2_X4 U2893 ( .A1(n3715), .A2(n3716), .ZN(n3718) );
  NAND2_X2 U2895 ( .A1(n1517), .A2(n4267), .ZN(n3904) );
  NOR2_X1 U2896 ( .A1(n2296), .A2(n4204), .ZN(n2293) );
  NAND2_X1 U2897 ( .A1(n2296), .A2(n4204), .ZN(n2300) );
  NAND2_X4 U2898 ( .A1(net296326), .A2(n2107), .ZN(n2108) );
  NOR2_X4 U2899 ( .A1(net298483), .A2(net297276), .ZN(net298482) );
  INV_X4 U2900 ( .A(n1923), .ZN(n1926) );
  NOR2_X4 U2901 ( .A1(n1870), .A2(n1871), .ZN(n1840) );
  INV_X4 U2902 ( .A(n1840), .ZN(n1750) );
  NAND4_X4 U2903 ( .A1(b[16]), .A2(control[0]), .A3(a[3]), .A4(net297172), 
        .ZN(n1923) );
  INV_X2 U2904 ( .A(n1711), .ZN(n1960) );
  NAND3_X4 U2905 ( .A1(n2177), .A2(n4258), .A3(n4249), .ZN(n2188) );
  NAND2_X4 U2906 ( .A1(net295754), .A2(net297526), .ZN(n2770) );
  OAI22_X4 U2907 ( .A1(n3778), .A2(n3779), .B1(n1768), .B2(n3779), .ZN(n3780)
         );
  NAND2_X1 U2908 ( .A1(n2199), .A2(n2229), .ZN(n2127) );
  AOI21_X2 U2910 ( .B1(n4275), .B2(net294448), .A(n3680), .ZN(n3670) );
  NAND2_X4 U2911 ( .A1(n2483), .A2(n1590), .ZN(n2312) );
  INV_X4 U2912 ( .A(n2197), .ZN(n1755) );
  NOR2_X4 U2913 ( .A1(n2370), .A2(n2369), .ZN(n2380) );
  INV_X2 U2914 ( .A(n2174), .ZN(n2148) );
  OAI21_X2 U2916 ( .B1(n3474), .B2(n3473), .A(n4044), .ZN(n3475) );
  NOR2_X2 U2918 ( .A1(net297166), .A2(net296909), .ZN(n1903) );
  NAND3_X4 U2919 ( .A1(net297166), .A2(net298225), .A3(b[10]), .ZN(n1820) );
  INV_X1 U2920 ( .A(n2496), .ZN(n2429) );
  NOR2_X4 U2921 ( .A1(n1277), .A2(n2205), .ZN(n2208) );
  NAND2_X4 U2922 ( .A1(net295273), .A2(n3319), .ZN(n3321) );
  INV_X4 U2923 ( .A(n1755), .ZN(n1756) );
  NAND2_X4 U2924 ( .A1(n3154), .A2(n3400), .ZN(n3246) );
  INV_X8 U2925 ( .A(n3246), .ZN(n3248) );
  NOR2_X2 U2926 ( .A1(n3402), .A2(n3515), .ZN(n3405) );
  NAND2_X4 U2927 ( .A1(n2413), .A2(n2412), .ZN(n2490) );
  NAND2_X4 U2928 ( .A1(n3299), .A2(n3300), .ZN(n3349) );
  NAND2_X4 U2930 ( .A1(a[6]), .A2(net297202), .ZN(n2654) );
  NAND2_X4 U2931 ( .A1(n3563), .A2(n3562), .ZN(n3421) );
  NAND2_X2 U2932 ( .A1(n3849), .A2(net294484), .ZN(n3850) );
  INV_X4 U2933 ( .A(n2989), .ZN(n2991) );
  NAND2_X2 U2935 ( .A1(n1691), .A2(n1246), .ZN(n1693) );
  NAND2_X2 U2936 ( .A1(net294792), .A2(net298829), .ZN(n1694) );
  NAND2_X4 U2937 ( .A1(net298388), .A2(net298389), .ZN(n1695) );
  NAND2_X4 U2938 ( .A1(n1694), .A2(n1695), .ZN(n3671) );
  INV_X4 U2939 ( .A(net294792), .ZN(net298388) );
  NAND2_X2 U2940 ( .A1(net299331), .A2(n3773), .ZN(n1697) );
  NAND2_X4 U2941 ( .A1(net298392), .A2(n1696), .ZN(n1698) );
  NAND2_X4 U2942 ( .A1(n1697), .A2(n1698), .ZN(n3906) );
  INV_X4 U2943 ( .A(n3773), .ZN(n1696) );
  NAND2_X4 U2944 ( .A1(n3671), .A2(net294791), .ZN(n3800) );
  NAND2_X4 U2945 ( .A1(n3906), .A2(net294388), .ZN(net294322) );
  NAND3_X2 U2946 ( .A1(n3175), .A2(net297254), .A3(a[12]), .ZN(n3458) );
  NAND2_X2 U2947 ( .A1(n1699), .A2(n1700), .ZN(n1702) );
  INV_X2 U2948 ( .A(n3670), .ZN(n1699) );
  INV_X4 U2949 ( .A(n3669), .ZN(n1700) );
  NAND2_X1 U2950 ( .A1(n3514), .A2(n3511), .ZN(n3340) );
  NAND2_X4 U2951 ( .A1(n3948), .A2(n3947), .ZN(n4014) );
  NAND3_X2 U2953 ( .A1(net298051), .A2(n1284), .A3(net298605), .ZN(n1988) );
  NAND2_X4 U2955 ( .A1(n3125), .A2(n2884), .ZN(n2711) );
  OAI21_X2 U2956 ( .B1(n2071), .B2(n2215), .A(n2214), .ZN(n2216) );
  XNOR2_X2 U2957 ( .A(n3714), .B(n1188), .ZN(product_out[25]) );
  NAND3_X2 U2958 ( .A1(n2315), .A2(n2314), .A3(n2313), .ZN(n1704) );
  NAND3_X2 U2959 ( .A1(n1163), .A2(n1602), .A3(n2311), .ZN(n2314) );
  NAND2_X4 U2960 ( .A1(n3229), .A2(n3228), .ZN(n3230) );
  INV_X2 U2961 ( .A(n2801), .ZN(n2803) );
  NOR3_X4 U2962 ( .A1(n1715), .A2(n3045), .A3(n2936), .ZN(n2849) );
  INV_X4 U2963 ( .A(n3871), .ZN(n3786) );
  INV_X4 U2964 ( .A(n3303), .ZN(n1705) );
  INV_X4 U2965 ( .A(n1959), .ZN(n1706) );
  NAND2_X4 U2966 ( .A1(n2969), .A2(n2970), .ZN(n3135) );
  NOR2_X1 U2967 ( .A1(n2227), .A2(n2226), .ZN(n2240) );
  NAND2_X1 U2968 ( .A1(n2227), .A2(n2226), .ZN(n2239) );
  NAND2_X2 U2969 ( .A1(n3930), .A2(n3929), .ZN(n1709) );
  NAND2_X2 U2970 ( .A1(n1710), .A2(n1709), .ZN(product_out[28]) );
  INV_X4 U2971 ( .A(n3930), .ZN(n1707) );
  NAND2_X2 U2972 ( .A1(n2493), .A2(n1625), .ZN(n2762) );
  INV_X2 U2973 ( .A(n3138), .ZN(n3058) );
  NAND2_X1 U2974 ( .A1(n2212), .A2(net296554), .ZN(n2215) );
  NAND2_X4 U2976 ( .A1(n1650), .A2(n1878), .ZN(n1981) );
  NAND2_X4 U2977 ( .A1(n3565), .A2(n1276), .ZN(n3684) );
  NAND3_X1 U2978 ( .A1(n3483), .A2(n3480), .A3(n3479), .ZN(n3487) );
  NOR2_X2 U2979 ( .A1(net296771), .A2(n2121), .ZN(n2123) );
  OAI22_X4 U2980 ( .A1(n1533), .A2(n3913), .B1(n3913), .B2(net294388), .ZN(
        n3908) );
  INV_X4 U2982 ( .A(net294448), .ZN(net294575) );
  NAND2_X4 U2983 ( .A1(n1867), .A2(n1932), .ZN(n1879) );
  AOI22_X4 U2984 ( .A1(n1713), .A2(n1931), .B1(n1873), .B2(n1872), .ZN(n1877)
         );
  NAND2_X4 U2986 ( .A1(n3251), .A2(n3252), .ZN(n3507) );
  NAND2_X2 U2988 ( .A1(n2452), .A2(n2534), .ZN(n1718) );
  NAND2_X4 U2989 ( .A1(n1716), .A2(n1717), .ZN(n1719) );
  NAND2_X4 U2990 ( .A1(n1718), .A2(n1719), .ZN(n2455) );
  INV_X4 U2991 ( .A(n2452), .ZN(n1716) );
  INV_X4 U2992 ( .A(n2534), .ZN(n1717) );
  NAND2_X1 U2994 ( .A1(n2368), .A2(n2367), .ZN(n2266) );
  NAND2_X4 U2995 ( .A1(net294301), .A2(n3936), .ZN(n3987) );
  NAND2_X4 U2996 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  NAND2_X2 U2997 ( .A1(net296324), .A2(net296326), .ZN(n2211) );
  OAI21_X2 U2998 ( .B1(n1511), .B2(n2608), .A(n2703), .ZN(n2610) );
  NAND2_X2 U2999 ( .A1(n2517), .A2(n2555), .ZN(n2352) );
  OAI211_X2 U3000 ( .C1(n4038), .C2(n4037), .A(n4036), .B(n4035), .ZN(n4104)
         );
  NAND3_X1 U3002 ( .A1(n3981), .A2(net294194), .A3(net294241), .ZN(n3978) );
  NOR2_X4 U3003 ( .A1(n4037), .A2(net294194), .ZN(n3982) );
  NAND2_X4 U3004 ( .A1(n3310), .A2(n3309), .ZN(n3345) );
  NAND2_X4 U3005 ( .A1(n2364), .A2(n2363), .ZN(n2459) );
  INV_X2 U3006 ( .A(n2477), .ZN(n2480) );
  NAND2_X2 U3007 ( .A1(n2009), .A2(n2008), .ZN(n2010) );
  NOR2_X1 U3008 ( .A1(n4109), .A2(n4280), .ZN(n4147) );
  NAND2_X1 U3009 ( .A1(n4020), .A2(n4021), .ZN(n4024) );
  INV_X2 U3010 ( .A(n3955), .ZN(n3957) );
  NAND2_X4 U3011 ( .A1(n3954), .A2(n3955), .ZN(n4008) );
  INV_X1 U3012 ( .A(n3653), .ZN(n3651) );
  NAND2_X4 U3013 ( .A1(n1887), .A2(n1952), .ZN(n1949) );
  NAND2_X4 U3014 ( .A1(n1945), .A2(n1944), .ZN(n1947) );
  NAND3_X2 U3015 ( .A1(n1939), .A2(n1564), .A3(n1940), .ZN(n1945) );
  NAND3_X2 U3016 ( .A1(n1940), .A2(n1564), .A3(n1937), .ZN(n1933) );
  NAND2_X4 U3017 ( .A1(net294578), .A2(net294446), .ZN(net294573) );
  INV_X2 U3018 ( .A(n2033), .ZN(n2031) );
  NAND2_X2 U3019 ( .A1(n2049), .A2(n2046), .ZN(n2030) );
  AOI21_X4 U3020 ( .B1(n3828), .B2(n1722), .A(n3724), .ZN(n3783) );
  NAND2_X4 U3021 ( .A1(n2193), .A2(n2192), .ZN(n2254) );
  NAND3_X2 U3022 ( .A1(n2285), .A2(n1721), .A3(n2191), .ZN(n2192) );
  INV_X4 U3023 ( .A(n3684), .ZN(n3686) );
  OAI22_X4 U3024 ( .A1(b[16]), .A2(net297182), .B1(b[24]), .B2(control[0]), 
        .ZN(n1860) );
  NAND2_X1 U3025 ( .A1(net294053), .A2(net294054), .ZN(n4096) );
  NAND2_X4 U3026 ( .A1(n2386), .A2(n2392), .ZN(n2393) );
  NAND2_X4 U3027 ( .A1(n2384), .A2(n2385), .ZN(n2392) );
  NAND2_X4 U3028 ( .A1(n2382), .A2(n2383), .ZN(n2386) );
  NOR2_X1 U3029 ( .A1(n3743), .A2(n1126), .ZN(n3611) );
  INV_X2 U3030 ( .A(n2974), .ZN(n2977) );
  INV_X1 U3031 ( .A(net296325), .ZN(net296547) );
  NAND2_X4 U3032 ( .A1(n2110), .A2(n2111), .ZN(n2223) );
  INV_X2 U3033 ( .A(net295732), .ZN(net295734) );
  NAND2_X4 U3034 ( .A1(n1900), .A2(n2013), .ZN(n1953) );
  NOR2_X4 U3035 ( .A1(net296554), .A2(n2321), .ZN(n2326) );
  NOR2_X4 U3036 ( .A1(n3119), .A2(n3120), .ZN(n3122) );
  NAND3_X2 U3037 ( .A1(n2871), .A2(n2782), .A3(n2781), .ZN(n2863) );
  NAND2_X4 U3038 ( .A1(n2861), .A2(n2863), .ZN(n2942) );
  AOI21_X1 U3039 ( .B1(n4014), .B2(n4271), .A(n4013), .ZN(n4016) );
  INV_X32 U3040 ( .A(control[0]), .ZN(net298225) );
  INV_X32 U3041 ( .A(control[0]), .ZN(net298226) );
  INV_X4 U3042 ( .A(n3158), .ZN(n3329) );
  OAI221_X4 U3043 ( .B1(n2197), .B2(n1527), .C1(n1756), .C2(n1219), .A(n2324), 
        .ZN(n2419) );
  INV_X1 U3044 ( .A(n1763), .ZN(n1722) );
  NAND2_X2 U3045 ( .A1(n2794), .A2(n2854), .ZN(n1725) );
  NAND2_X4 U3046 ( .A1(n1723), .A2(n1724), .ZN(n1726) );
  NAND2_X4 U3047 ( .A1(n1725), .A2(n1726), .ZN(n2842) );
  INV_X4 U3048 ( .A(n2794), .ZN(n1723) );
  INV_X1 U3049 ( .A(n2854), .ZN(n1724) );
  NAND2_X2 U3050 ( .A1(n2879), .A2(n2921), .ZN(n1729) );
  NAND2_X4 U3051 ( .A1(n1727), .A2(n1728), .ZN(n1730) );
  INV_X4 U3052 ( .A(n2879), .ZN(n1727) );
  INV_X1 U3053 ( .A(n2921), .ZN(n1728) );
  NAND2_X2 U3054 ( .A1(n2424), .A2(n1302), .ZN(n1733) );
  NAND2_X4 U3055 ( .A1(n1731), .A2(n1732), .ZN(n1734) );
  NAND2_X4 U3056 ( .A1(n1734), .A2(n1733), .ZN(n2568) );
  INV_X4 U3057 ( .A(n2424), .ZN(n1731) );
  NAND2_X4 U3058 ( .A1(n1736), .A2(n1737), .ZN(n2227) );
  NAND2_X2 U3059 ( .A1(n1915), .A2(n1914), .ZN(n1740) );
  NAND2_X4 U3060 ( .A1(n1738), .A2(n1739), .ZN(n1741) );
  NAND2_X4 U3061 ( .A1(n1741), .A2(n1740), .ZN(n1989) );
  INV_X8 U3062 ( .A(n1915), .ZN(n1738) );
  NAND2_X4 U3063 ( .A1(n2880), .A2(n2922), .ZN(n3127) );
  INV_X8 U3064 ( .A(n1989), .ZN(n2114) );
  NAND3_X4 U3065 ( .A1(n2329), .A2(n1757), .A3(net296524), .ZN(n2330) );
  NAND2_X4 U3066 ( .A1(n1642), .A2(n2008), .ZN(n1954) );
  INV_X4 U3067 ( .A(n2056), .ZN(n1900) );
  XNOR2_X1 U3069 ( .A(n2375), .B(n2373), .ZN(n2262) );
  NAND2_X4 U3070 ( .A1(n3091), .A2(n3090), .ZN(n3093) );
  NAND2_X4 U3071 ( .A1(n2496), .A2(n2687), .ZN(n2579) );
  INV_X8 U3072 ( .A(n3859), .ZN(n3441) );
  INV_X2 U3073 ( .A(n2331), .ZN(n2329) );
  INV_X8 U3074 ( .A(n2752), .ZN(n2788) );
  NAND2_X2 U3076 ( .A1(n3855), .A2(n3856), .ZN(n3857) );
  NAND4_X4 U3077 ( .A1(b[1]), .A2(net297166), .A3(a[2]), .A4(control[0]), .ZN(
        n1918) );
  NOR2_X2 U3078 ( .A1(n1869), .A2(n1868), .ZN(n1873) );
  INV_X8 U3079 ( .A(n3092), .ZN(n3011) );
  NAND2_X1 U3080 ( .A1(a[29]), .A2(net297272), .ZN(n4005) );
  NAND2_X4 U3081 ( .A1(n3938), .A2(n3937), .ZN(n3878) );
  NAND2_X4 U3082 ( .A1(n2158), .A2(n2157), .ZN(n2173) );
  NAND2_X4 U3083 ( .A1(n1742), .A2(n2570), .ZN(n2471) );
  OAI211_X2 U3084 ( .C1(n1134), .C2(n2701), .A(n2576), .B(n2575), .ZN(n2609)
         );
  NAND2_X4 U3085 ( .A1(n3493), .A2(n3494), .ZN(n3495) );
  NAND3_X2 U3086 ( .A1(n2428), .A2(n2427), .A3(n2470), .ZN(n2431) );
  OAI21_X4 U3087 ( .B1(n2583), .B2(n2584), .A(n2582), .ZN(n2602) );
  NAND2_X1 U3088 ( .A1(n3854), .A2(n4054), .ZN(n3869) );
  NOR2_X2 U3089 ( .A1(n4100), .A2(n4091), .ZN(n4077) );
  NAND2_X2 U3090 ( .A1(n4081), .A2(n4080), .ZN(n4082) );
  INV_X4 U3091 ( .A(net294908), .ZN(net294910) );
  NAND2_X4 U3092 ( .A1(n3591), .A2(n3590), .ZN(n3645) );
  NAND2_X4 U3093 ( .A1(n3945), .A2(n3944), .ZN(n3998) );
  NAND2_X4 U3094 ( .A1(n3889), .A2(n3888), .ZN(n3948) );
  NAND4_X4 U3095 ( .A1(n1909), .A2(net297022), .A3(n1908), .A4(n1907), .ZN(
        n1915) );
  AOI21_X2 U3096 ( .B1(n1782), .B2(n1556), .A(n1796), .ZN(n2069) );
  NAND2_X4 U3097 ( .A1(n2316), .A2(n2131), .ZN(n2076) );
  INV_X8 U3098 ( .A(n3622), .ZN(n4063) );
  INV_X4 U3099 ( .A(n3857), .ZN(n3861) );
  INV_X1 U3100 ( .A(n1772), .ZN(n3279) );
  INV_X2 U3101 ( .A(n2332), .ZN(n1757) );
  NAND2_X4 U3102 ( .A1(n1687), .A2(n1332), .ZN(n3378) );
  NAND2_X4 U3103 ( .A1(n3079), .A2(n3078), .ZN(n3305) );
  OAI211_X2 U3104 ( .C1(n3308), .C2(n3307), .A(n1361), .B(n3492), .ZN(n3309)
         );
  NAND2_X4 U3105 ( .A1(a[10]), .A2(net297272), .ZN(net296424) );
  OAI22_X4 U3106 ( .A1(net295864), .A2(n2872), .B1(net299089), .B2(n2963), 
        .ZN(n2959) );
  NAND4_X4 U3107 ( .A1(b[8]), .A2(net297166), .A3(a[3]), .A4(net297184), .ZN(
        n1924) );
  NAND2_X4 U3108 ( .A1(n3067), .A2(n3256), .ZN(n3163) );
  NAND3_X4 U3109 ( .A1(n2495), .A2(net298909), .A3(n2494), .ZN(n2687) );
  OAI21_X4 U3110 ( .B1(n2420), .B2(net295995), .A(net295991), .ZN(n2495) );
  NAND2_X4 U3111 ( .A1(n1882), .A2(n1940), .ZN(n1883) );
  NAND2_X4 U3112 ( .A1(n3749), .A2(n3748), .ZN(n3750) );
  NAND2_X4 U3113 ( .A1(n1765), .A2(net297862), .ZN(n1767) );
  NAND2_X4 U3114 ( .A1(n2718), .A2(n2733), .ZN(n2719) );
  NAND2_X4 U3115 ( .A1(n2681), .A2(n2680), .ZN(n2682) );
  NAND2_X4 U3116 ( .A1(n2679), .A2(net295749), .ZN(n2680) );
  NAND2_X4 U3117 ( .A1(n2865), .A2(n1691), .ZN(n2958) );
  NAND2_X2 U3118 ( .A1(n4161), .A2(n4159), .ZN(n4157) );
  OAI211_X4 U3119 ( .C1(n1562), .C2(net297279), .A(n4096), .B(n4095), .ZN(
        n4165) );
  NAND3_X1 U3121 ( .A1(net296324), .A2(net296325), .A3(net296326), .ZN(n2586)
         );
  NAND4_X2 U3122 ( .A1(a[2]), .A2(n1981), .A3(net294175), .A4(n2196), .ZN(
        n1884) );
  NAND2_X2 U3123 ( .A1(n3721), .A2(n3709), .ZN(n3828) );
  NAND2_X4 U3124 ( .A1(n2956), .A2(n2601), .ZN(n2764) );
  NAND2_X2 U3125 ( .A1(n2939), .A2(n3043), .ZN(n2921) );
  NOR2_X4 U3126 ( .A1(n2910), .A2(n2911), .ZN(n2912) );
  INV_X8 U3127 ( .A(n2797), .ZN(n2848) );
  NAND2_X4 U3128 ( .A1(n2924), .A2(n2925), .ZN(n2879) );
  NAND2_X2 U3129 ( .A1(n2790), .A2(n2855), .ZN(n2791) );
  OAI21_X4 U3130 ( .B1(n2581), .B2(n2580), .A(n2866), .ZN(n2582) );
  NAND2_X4 U3131 ( .A1(n1641), .A2(n2951), .ZN(n3048) );
  NAND2_X4 U3132 ( .A1(net294196), .A2(net294044), .ZN(n4078) );
  NAND2_X4 U3133 ( .A1(n2469), .A2(n2470), .ZN(n1742) );
  INV_X4 U3134 ( .A(n2083), .ZN(n1743) );
  AND2_X2 U3135 ( .A1(n3194), .A2(n3195), .ZN(n1744) );
  NOR2_X2 U3136 ( .A1(n1744), .A2(net299240), .ZN(n3197) );
  AND2_X2 U3137 ( .A1(n3777), .A2(n1162), .ZN(n1769) );
  INV_X2 U3138 ( .A(n2871), .ZN(n2778) );
  NAND2_X4 U3139 ( .A1(n2871), .A2(net295750), .ZN(net295866) );
  AOI21_X4 U3140 ( .B1(net294575), .B2(net294446), .A(net294576), .ZN(
        net294574) );
  NAND2_X1 U3141 ( .A1(n3632), .A2(n4293), .ZN(n3635) );
  NAND2_X4 U3142 ( .A1(n3456), .A2(n3552), .ZN(n3859) );
  INV_X4 U3143 ( .A(n2505), .ZN(n2573) );
  NAND2_X4 U3144 ( .A1(n2505), .A2(n2504), .ZN(n2607) );
  NAND2_X4 U3145 ( .A1(n1199), .A2(n3135), .ZN(n2978) );
  INV_X1 U3146 ( .A(n3885), .ZN(n3810) );
  NAND2_X4 U3147 ( .A1(n2195), .A2(n1527), .ZN(n1930) );
  AOI21_X4 U3148 ( .B1(n2101), .B2(n1706), .A(n1770), .ZN(n2102) );
  NAND2_X2 U3149 ( .A1(n2282), .A2(n2283), .ZN(n2284) );
  OAI211_X2 U3150 ( .C1(n1174), .C2(n4090), .A(n4042), .B(net297196), .ZN(
        n4074) );
  INV_X4 U3151 ( .A(n1340), .ZN(n2882) );
  INV_X1 U3152 ( .A(n2758), .ZN(n2763) );
  NAND2_X1 U3153 ( .A1(n4185), .A2(n4184), .ZN(n1747) );
  NAND2_X4 U3154 ( .A1(n1745), .A2(n1746), .ZN(n1748) );
  NAND2_X2 U3155 ( .A1(n1747), .A2(n1748), .ZN(product_out[31]) );
  INV_X4 U3156 ( .A(n4185), .ZN(n1745) );
  INV_X4 U3157 ( .A(n4184), .ZN(n1746) );
  NAND2_X4 U3158 ( .A1(net297281), .A2(a[4]), .ZN(n1878) );
  NAND2_X2 U3159 ( .A1(n1841), .A2(n1840), .ZN(n1751) );
  NAND2_X4 U3160 ( .A1(n1749), .A2(n1750), .ZN(n1752) );
  NAND2_X4 U3161 ( .A1(n1751), .A2(n1752), .ZN(n1881) );
  INV_X2 U3162 ( .A(n1841), .ZN(n1749) );
  NAND2_X4 U3163 ( .A1(n1842), .A2(n1881), .ZN(n1858) );
  INV_X4 U3164 ( .A(n1881), .ZN(n1843) );
  NAND2_X1 U3165 ( .A1(n2957), .A2(n2958), .ZN(n2870) );
  INV_X8 U3166 ( .A(n2976), .ZN(n2952) );
  OAI21_X4 U3167 ( .B1(n2947), .B2(n3051), .A(n3050), .ZN(n2975) );
  NAND2_X2 U3168 ( .A1(n3050), .A2(n3048), .ZN(n2875) );
  NAND2_X4 U3169 ( .A1(n2874), .A2(n1266), .ZN(n3050) );
  INV_X1 U3170 ( .A(n2949), .ZN(n2746) );
  NOR2_X1 U3171 ( .A1(n2746), .A2(n2795), .ZN(n2754) );
  INV_X4 U3173 ( .A(n2204), .ZN(n1782) );
  NOR2_X2 U3174 ( .A1(n3130), .A2(n3071), .ZN(n2930) );
  NAND2_X2 U3175 ( .A1(n2055), .A2(n1567), .ZN(n1753) );
  NAND2_X4 U3176 ( .A1(n1754), .A2(n2054), .ZN(n2135) );
  INV_X4 U3177 ( .A(n1753), .ZN(n1754) );
  NAND2_X4 U3178 ( .A1(n1599), .A2(n1896), .ZN(n2026) );
  INV_X8 U3179 ( .A(n2295), .ZN(n2317) );
  NAND2_X4 U3180 ( .A1(n2202), .A2(n2201), .ZN(net296324) );
  OAI21_X4 U3181 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3868) );
  NAND2_X2 U3182 ( .A1(n1761), .A2(n1762), .ZN(n4073) );
  INV_X1 U3183 ( .A(n1350), .ZN(n1760) );
  NAND3_X1 U3185 ( .A1(n4098), .A2(n4085), .A3(n4079), .ZN(n4080) );
  INV_X8 U3186 ( .A(n4085), .ZN(n4100) );
  NOR2_X1 U3187 ( .A1(net297276), .A2(n1807), .ZN(n1809) );
  NOR2_X1 U3188 ( .A1(net297276), .A2(n4118), .ZN(n4119) );
  INV_X4 U3189 ( .A(net299323), .ZN(net296672) );
  NAND2_X4 U3190 ( .A1(n2447), .A2(n2448), .ZN(n2660) );
  NAND2_X4 U3191 ( .A1(n1957), .A2(n1553), .ZN(n2097) );
  NAND2_X4 U3192 ( .A1(n1263), .A2(n3713), .ZN(n4061) );
  NAND2_X4 U3193 ( .A1(n3785), .A2(net297190), .ZN(n3713) );
  NOR3_X4 U3194 ( .A1(n3861), .A2(n1226), .A3(n3860), .ZN(n3864) );
  NOR2_X4 U3195 ( .A1(n2414), .A2(n1803), .ZN(n2416) );
  NAND2_X4 U3196 ( .A1(n1244), .A2(n1798), .ZN(n3920) );
  OAI21_X4 U3197 ( .B1(n3993), .B2(net297188), .A(n3351), .ZN(n3456) );
  NAND2_X4 U3198 ( .A1(n2751), .A2(n1573), .ZN(n2790) );
  NAND2_X4 U3199 ( .A1(n2750), .A2(n2703), .ZN(n2752) );
  INV_X4 U3200 ( .A(n2344), .ZN(n2346) );
  NAND2_X4 U3201 ( .A1(a[2]), .A2(net294175), .ZN(n1880) );
  INV_X2 U3202 ( .A(n1782), .ZN(n1764) );
  INV_X4 U3203 ( .A(net294322), .ZN(net294364) );
  NOR2_X2 U3204 ( .A1(net294367), .A2(net299020), .ZN(n3919) );
  NOR2_X1 U3205 ( .A1(n3290), .A2(n3298), .ZN(n3289) );
  INV_X2 U3206 ( .A(n3298), .ZN(n3921) );
  XNOR2_X1 U3207 ( .A(n2728), .B(n1147), .ZN(product_out[14]) );
  NAND2_X4 U3208 ( .A1(n3362), .A2(n3363), .ZN(n3365) );
  INV_X2 U3209 ( .A(n3828), .ZN(n3841) );
  INV_X4 U3210 ( .A(n3037), .ZN(n3042) );
  AOI21_X1 U3211 ( .B1(net294053), .B2(n1605), .A(n3923), .ZN(n3925) );
  INV_X2 U3212 ( .A(n2449), .ZN(n2447) );
  NOR2_X4 U3213 ( .A1(n3175), .A2(n1773), .ZN(n1772) );
  INV_X4 U3214 ( .A(n1530), .ZN(n3388) );
  NAND2_X4 U3215 ( .A1(n2717), .A2(n2993), .ZN(n2729) );
  OAI221_X4 U3216 ( .B1(n1763), .B2(n3877), .C1(n3876), .C2(n1763), .A(n3875), 
        .ZN(net294087) );
  NAND2_X2 U3217 ( .A1(n3131), .A2(n3230), .ZN(n3171) );
  NAND2_X1 U3218 ( .A1(n3852), .A2(n1232), .ZN(n1766) );
  NAND2_X2 U3219 ( .A1(n1766), .A2(n1767), .ZN(product_out[27]) );
  INV_X4 U3220 ( .A(n3852), .ZN(n1765) );
  NAND3_X4 U3221 ( .A1(n3025), .A2(n3034), .A3(n1576), .ZN(n3327) );
  NAND2_X4 U3222 ( .A1(n3034), .A2(n3035), .ZN(n3159) );
  NAND2_X2 U3224 ( .A1(n3905), .A2(n3799), .ZN(net294310) );
  NAND4_X4 U3225 ( .A1(b[17]), .A2(control[0]), .A3(a[2]), .A4(net297170), 
        .ZN(n1928) );
  NAND2_X4 U3226 ( .A1(n2660), .A2(n2651), .ZN(n2534) );
  NAND2_X4 U3227 ( .A1(n3973), .A2(n3974), .ZN(n4033) );
  NAND2_X4 U3229 ( .A1(n2156), .A2(n2155), .ZN(n2276) );
  NAND3_X1 U3230 ( .A1(a[25]), .A2(n3753), .A3(net297274), .ZN(n3805) );
  NAND2_X1 U3231 ( .A1(a[26]), .A2(net297274), .ZN(n3804) );
  NAND2_X1 U3232 ( .A1(a[25]), .A2(net297274), .ZN(n3751) );
  NAND2_X1 U3233 ( .A1(a[24]), .A2(net297274), .ZN(n3649) );
  NAND2_X1 U3234 ( .A1(a[22]), .A2(net297274), .ZN(n3522) );
  NAND3_X2 U3235 ( .A1(n4069), .A2(n4175), .A3(net293935), .ZN(n4070) );
  NAND3_X1 U3237 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n3632) );
  NAND2_X2 U3238 ( .A1(n3469), .A2(n3470), .ZN(n3471) );
  INV_X4 U3239 ( .A(n1770), .ZN(n1771) );
  NAND2_X4 U3240 ( .A1(n3886), .A2(n3885), .ZN(n3950) );
  NAND2_X4 U3241 ( .A1(n3826), .A2(net294515), .ZN(n3842) );
  NAND2_X4 U3242 ( .A1(n3394), .A2(n1535), .ZN(n3508) );
  NAND2_X4 U3243 ( .A1(n3907), .A2(n3908), .ZN(net294331) );
  OAI221_X4 U3244 ( .B1(net294126), .B2(n3618), .C1(n3617), .C2(net294048), 
        .A(n3616), .ZN(n3622) );
  INV_X2 U3245 ( .A(n1523), .ZN(n3834) );
  AND2_X4 U3246 ( .A1(a[12]), .A2(net297254), .ZN(n1773) );
  NAND3_X4 U3247 ( .A1(n3496), .A2(n3495), .A3(n1360), .ZN(n3569) );
  NAND2_X4 U3249 ( .A1(n2317), .A2(n2316), .ZN(n2491) );
  OAI21_X4 U3251 ( .B1(n3868), .B2(n3869), .A(n3867), .ZN(n3870) );
  XNOR2_X1 U3252 ( .A(n1290), .B(n1539), .ZN(product_out[13]) );
  AOI21_X2 U3253 ( .B1(n2291), .B2(n2334), .A(n2137), .ZN(n2138) );
  OAI22_X4 U3254 ( .A1(net294048), .A2(net296472), .B1(net298860), .B2(
        net297190), .ZN(n2384) );
  NAND2_X1 U3255 ( .A1(n2854), .A2(n2844), .ZN(n2786) );
  NAND2_X1 U3257 ( .A1(n4196), .A2(n1851), .ZN(n1854) );
  NAND2_X4 U3258 ( .A1(n3305), .A2(n3490), .ZN(n3225) );
  INV_X4 U3259 ( .A(n1589), .ZN(n3024) );
  INV_X1 U3260 ( .A(n2950), .ZN(n2851) );
  NAND2_X4 U3261 ( .A1(n2179), .A2(n2180), .ZN(n2183) );
  OAI21_X4 U3262 ( .B1(n2977), .B2(n1542), .A(n2975), .ZN(n2979) );
  INV_X4 U3263 ( .A(n2438), .ZN(n2439) );
  INV_X8 U3264 ( .A(n2200), .ZN(n2418) );
  NAND2_X4 U3265 ( .A1(n1795), .A2(n2199), .ZN(n2200) );
  NAND2_X4 U3266 ( .A1(n3013), .A2(n3012), .ZN(n3281) );
  NAND2_X4 U3267 ( .A1(n3605), .A2(n3531), .ZN(net297774) );
  NAND2_X4 U3268 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  OAI21_X2 U3269 ( .B1(n3731), .B2(n3730), .A(net294701), .ZN(n3740) );
  INV_X8 U3272 ( .A(net294321), .ZN(net294510) );
  INV_X4 U3273 ( .A(n2195), .ZN(n1876) );
  NAND2_X1 U3274 ( .A1(n2425), .A2(n1625), .ZN(n2426) );
  OAI21_X4 U3275 ( .B1(n1274), .B2(n2198), .A(n2232), .ZN(n2136) );
  NAND3_X2 U3276 ( .A1(n4183), .A2(n4182), .A3(n4181), .ZN(n4184) );
  NAND2_X4 U3277 ( .A1(n2453), .A2(n2454), .ZN(n2457) );
  NAND2_X4 U3278 ( .A1(n1495), .A2(net294525), .ZN(net294330) );
  INV_X8 U3279 ( .A(n2537), .ZN(n2630) );
  NAND2_X4 U3280 ( .A1(n2275), .A2(n2276), .ZN(n2375) );
  NAND3_X4 U3281 ( .A1(a[17]), .A2(net295372), .A3(net297226), .ZN(n3401) );
  XNOR2_X2 U3283 ( .A(n2149), .B(n1721), .ZN(n2150) );
  NAND2_X1 U3284 ( .A1(n3134), .A2(n4200), .ZN(n3066) );
  NAND4_X2 U3285 ( .A1(n3128), .A2(n1328), .A3(n2884), .A4(n2917), .ZN(n2885)
         );
  NAND2_X4 U3286 ( .A1(n1777), .A2(n1778), .ZN(n1780) );
  NAND2_X4 U3287 ( .A1(n1780), .A2(n1779), .ZN(n2344) );
  INV_X4 U3288 ( .A(n2342), .ZN(n1777) );
  NAND2_X4 U3289 ( .A1(n1781), .A2(n1782), .ZN(n1784) );
  NAND2_X4 U3290 ( .A1(n1783), .A2(n1784), .ZN(n2005) );
  INV_X4 U3291 ( .A(n2004), .ZN(n1781) );
  INV_X4 U3292 ( .A(n2975), .ZN(n2948) );
  NAND2_X4 U3293 ( .A1(n2591), .A2(n2590), .ZN(n2679) );
  NAND2_X4 U3294 ( .A1(n2864), .A2(n1105), .ZN(n2960) );
  NAND2_X4 U3295 ( .A1(n2862), .A2(n2861), .ZN(n2864) );
  NAND2_X4 U3296 ( .A1(n2868), .A2(n2766), .ZN(n2954) );
  INV_X8 U3297 ( .A(n2960), .ZN(n2957) );
  NAND2_X4 U3298 ( .A1(n1496), .A2(n2020), .ZN(n2104) );
  NAND2_X2 U3299 ( .A1(n2841), .A2(n3037), .ZN(n2933) );
  INV_X16 U3300 ( .A(n1795), .ZN(n1796) );
  NAND3_X2 U3301 ( .A1(n2119), .A2(n2117), .A3(n1643), .ZN(n2221) );
  NAND2_X4 U3302 ( .A1(net299240), .A2(n3195), .ZN(n3191) );
  NAND2_X4 U3303 ( .A1(n2093), .A2(n1106), .ZN(n2282) );
  NAND2_X4 U3304 ( .A1(n2419), .A2(n1168), .ZN(net296419) );
  NOR2_X1 U3305 ( .A1(n3830), .A2(n4270), .ZN(n3832) );
  OAI21_X2 U3306 ( .B1(n3775), .B2(n3910), .A(n4215), .ZN(n3778) );
  NOR2_X2 U3307 ( .A1(n3045), .A2(n2932), .ZN(n2934) );
  NAND2_X4 U3308 ( .A1(n2777), .A2(net295978), .ZN(n2871) );
  NAND4_X4 U3309 ( .A1(b[9]), .A2(control[1]), .A3(a[2]), .A4(net297180), .ZN(
        n1919) );
  NAND3_X2 U3310 ( .A1(n3236), .A2(n3058), .A3(n3239), .ZN(n3059) );
  NAND2_X4 U3311 ( .A1(n2756), .A2(n2765), .ZN(n2755) );
  NAND3_X1 U3312 ( .A1(n1573), .A2(n2672), .A3(n2611), .ZN(n2605) );
  NAND3_X2 U3313 ( .A1(n2315), .A2(n2313), .A3(n2314), .ZN(n2433) );
  NAND2_X4 U3314 ( .A1(n2222), .A2(n2223), .ZN(n2112) );
  AOI21_X2 U3315 ( .B1(n2338), .B2(n2415), .A(n2337), .ZN(n2339) );
  NOR2_X4 U3316 ( .A1(n3572), .A2(n4268), .ZN(n3576) );
  NAND2_X4 U3317 ( .A1(net297481), .A2(a[7]), .ZN(n2065) );
  NOR2_X2 U3318 ( .A1(n3146), .A2(n3235), .ZN(n3149) );
  NAND2_X1 U3319 ( .A1(n2817), .A2(n2816), .ZN(n2728) );
  NAND2_X4 U3320 ( .A1(n3798), .A2(n4215), .ZN(n3722) );
  NAND2_X4 U3321 ( .A1(n2540), .A2(n2539), .ZN(n2634) );
  OAI21_X4 U3322 ( .B1(n2530), .B2(n2661), .A(n2529), .ZN(n2533) );
  NAND3_X2 U3323 ( .A1(n2651), .A2(n2625), .A3(n2626), .ZN(n2529) );
  NAND2_X4 U3324 ( .A1(n1917), .A2(n1916), .ZN(n1867) );
  NOR2_X2 U3325 ( .A1(n1951), .A2(n1952), .ZN(n1956) );
  OAI21_X4 U3326 ( .B1(n1275), .B2(n3915), .A(n3914), .ZN(net294332) );
  NOR2_X2 U3327 ( .A1(n3912), .A2(n3911), .ZN(n3915) );
  NAND3_X4 U3328 ( .A1(n3629), .A2(n3630), .A3(n3628), .ZN(n3566) );
  OAI211_X4 U3329 ( .C1(n2240), .C2(n2292), .A(n2238), .B(n2239), .ZN(n2241)
         );
  NOR3_X4 U3330 ( .A1(n1821), .A2(control[0]), .A3(net297168), .ZN(n1824) );
  NAND2_X4 U3331 ( .A1(a[1]), .A2(net297230), .ZN(n1952) );
  INV_X16 U3332 ( .A(n1426), .ZN(net297230) );
  NAND2_X4 U3333 ( .A1(n1310), .A2(n2351), .ZN(n2555) );
  NAND3_X2 U3335 ( .A1(control[0]), .A2(net297168), .A3(n1792), .ZN(n1910) );
  INV_X2 U3336 ( .A(n1791), .ZN(n1792) );
  OAI21_X4 U3337 ( .B1(n3575), .B2(n3576), .A(n4261), .ZN(n3612) );
  NAND2_X4 U3338 ( .A1(n3142), .A2(n4272), .ZN(n3139) );
  INV_X32 U3339 ( .A(a[5]), .ZN(net296909) );
  NAND2_X4 U3340 ( .A1(n2255), .A2(n2398), .ZN(n2515) );
  AOI21_X2 U3341 ( .B1(n2334), .B2(n1505), .A(n2094), .ZN(n2078) );
  NAND2_X4 U3342 ( .A1(n1881), .A2(n1982), .ZN(n1940) );
  INV_X4 U3343 ( .A(n4170), .ZN(n4158) );
  NAND2_X4 U3344 ( .A1(n1844), .A2(n1843), .ZN(n1859) );
  NAND2_X4 U3345 ( .A1(n3024), .A2(n3023), .ZN(n3043) );
  NAND2_X4 U3346 ( .A1(n2852), .A2(n2950), .ZN(n2854) );
  NAND2_X4 U3348 ( .A1(n3723), .A2(n3831), .ZN(n3725) );
  NAND2_X4 U3349 ( .A1(net295017), .A2(n3524), .ZN(n3590) );
  OAI21_X2 U3350 ( .B1(n3524), .B2(n4264), .A(n3590), .ZN(net295013) );
  NAND2_X4 U3351 ( .A1(n3807), .A2(n3808), .ZN(n3885) );
  INV_X32 U3353 ( .A(b[8]), .ZN(n1786) );
  NAND2_X4 U3354 ( .A1(n2434), .A2(n2435), .ZN(n2436) );
  NAND3_X2 U3355 ( .A1(n2116), .A2(n2114), .A3(n2115), .ZN(n2066) );
  NAND4_X4 U3356 ( .A1(b[25]), .A2(net299325), .A3(a[4]), .A4(net298226), .ZN(
        n1913) );
  NAND4_X4 U3357 ( .A1(b[9]), .A2(control[1]), .A3(a[4]), .A4(net298225), .ZN(
        n1911) );
  NAND2_X4 U3358 ( .A1(n1911), .A2(n1913), .ZN(n1789) );
  NAND2_X4 U3359 ( .A1(n2814), .A2(n3007), .ZN(n2828) );
  NAND2_X4 U3360 ( .A1(n1366), .A2(n2813), .ZN(n3007) );
  INV_X4 U3361 ( .A(n2906), .ZN(n2911) );
  NAND2_X4 U3362 ( .A1(n3259), .A2(n3068), .ZN(n3334) );
  NAND3_X4 U3363 ( .A1(net297168), .A2(control[0]), .A3(b[2]), .ZN(n1822) );
  NAND2_X2 U3364 ( .A1(n2402), .A2(n2403), .ZN(n2406) );
  NAND3_X2 U3365 ( .A1(n1924), .A2(n1586), .A3(net297002), .ZN(n1925) );
  INV_X4 U3366 ( .A(n3712), .ZN(n1787) );
  INV_X1 U3367 ( .A(n3712), .ZN(n4067) );
  OAI22_X4 U3368 ( .A1(n1832), .A2(n1831), .B1(n1829), .B2(n1830), .ZN(n1838)
         );
  NAND3_X1 U3369 ( .A1(net297182), .A2(n1906), .A3(a[6]), .ZN(n2002) );
  NAND2_X1 U3370 ( .A1(n1919), .A2(n1918), .ZN(n1922) );
  NAND2_X2 U3372 ( .A1(a[7]), .A2(net296932), .ZN(n2122) );
  INV_X4 U3373 ( .A(n3191), .ZN(n3193) );
  INV_X4 U3374 ( .A(n1742), .ZN(n2571) );
  OAI21_X2 U3375 ( .B1(n3332), .B2(n3333), .A(n3507), .ZN(n3338) );
  NAND2_X1 U3376 ( .A1(n2570), .A2(n2472), .ZN(n2435) );
  NOR2_X4 U3377 ( .A1(n2907), .A2(n1259), .ZN(n1788) );
  INV_X4 U3378 ( .A(n1788), .ZN(n2902) );
  NAND2_X4 U3379 ( .A1(n2176), .A2(n2177), .ZN(n2084) );
  NAND2_X4 U3380 ( .A1(n2164), .A2(n2165), .ZN(n2264) );
  NOR2_X2 U3381 ( .A1(n3373), .A2(n3372), .ZN(n3379) );
  NAND2_X4 U3382 ( .A1(n2531), .A2(n2532), .ZN(n2730) );
  OAI211_X4 U3383 ( .C1(n1641), .C2(n2951), .A(n2950), .B(n2949), .ZN(n2976)
         );
  INV_X4 U3384 ( .A(n3667), .ZN(n3664) );
  NAND2_X4 U3385 ( .A1(n2734), .A2(n1545), .ZN(n2635) );
  NAND2_X4 U3386 ( .A1(n2265), .A2(n2264), .ZN(n2368) );
  NAND3_X2 U3387 ( .A1(n1790), .A2(n1910), .A3(n1912), .ZN(n1914) );
  INV_X4 U3388 ( .A(n1789), .ZN(n1790) );
  NAND2_X2 U3389 ( .A1(b[1]), .A2(a[4]), .ZN(n1791) );
  NAND3_X1 U3390 ( .A1(n2925), .A2(n2924), .A3(n2923), .ZN(n2926) );
  NAND2_X4 U3391 ( .A1(n1800), .A2(n2850), .ZN(n2855) );
  NAND2_X4 U3392 ( .A1(n2573), .A2(n2574), .ZN(n2703) );
  NAND2_X4 U3393 ( .A1(n2473), .A2(n1794), .ZN(n2474) );
  NAND3_X2 U3394 ( .A1(n1377), .A2(n2309), .A3(n2310), .ZN(n2473) );
  NAND2_X4 U3395 ( .A1(n3627), .A2(n3626), .ZN(n3703) );
  NAND2_X4 U3396 ( .A1(n3380), .A2(n3497), .ZN(n3562) );
  INV_X8 U3398 ( .A(n2845), .ZN(n2937) );
  NAND2_X4 U3399 ( .A1(n2633), .A2(n2634), .ZN(n2734) );
  NAND2_X2 U3401 ( .A1(n1949), .A2(n2096), .ZN(n1890) );
  NAND2_X4 U3402 ( .A1(n1888), .A2(n1889), .ZN(n2096) );
  NAND2_X4 U3403 ( .A1(n3425), .A2(n3561), .ZN(n3298) );
  NAND2_X4 U3404 ( .A1(n3277), .A2(n3276), .ZN(n3561) );
  NAND2_X4 U3405 ( .A1(n2173), .A2(n2172), .ZN(n2275) );
  NAND2_X2 U3406 ( .A1(n3504), .A2(n1112), .ZN(n3608) );
  INV_X8 U3407 ( .A(n1796), .ZN(n2198) );
  NAND2_X4 U3408 ( .A1(n3823), .A2(n3939), .ZN(n3940) );
  NAND3_X2 U3409 ( .A1(n3661), .A2(net294815), .A3(net294816), .ZN(n3663) );
  INV_X2 U3410 ( .A(n3594), .ZN(n3592) );
  NAND2_X4 U3411 ( .A1(n2053), .A2(n1771), .ZN(n1980) );
  NAND2_X4 U3412 ( .A1(n2457), .A2(n2542), .ZN(n2543) );
  NAND2_X4 U3413 ( .A1(n2456), .A2(n2455), .ZN(n2542) );
  NAND2_X4 U3414 ( .A1(n2614), .A2(n1373), .ZN(n2441) );
  NOR2_X4 U3415 ( .A1(n4177), .A2(n4176), .ZN(n4072) );
  NAND4_X2 U3416 ( .A1(n2126), .A2(n1370), .A3(n2220), .A4(n2226), .ZN(n2125)
         );
  NAND2_X4 U3417 ( .A1(n2018), .A2(n2019), .ZN(n2301) );
  NAND2_X2 U3418 ( .A1(n2663), .A2(n2651), .ZN(n2629) );
  NAND2_X4 U3419 ( .A1(net294359), .A2(net294358), .ZN(net294349) );
  NAND3_X2 U3420 ( .A1(n2433), .A2(n1314), .A3(n2570), .ZN(n2434) );
  OAI22_X4 U3421 ( .A1(n1835), .A2(n1836), .B1(n1833), .B2(n1834), .ZN(n1837)
         );
  NAND2_X1 U3422 ( .A1(n1897), .A2(n2026), .ZN(n3922) );
  NAND2_X1 U3423 ( .A1(n1894), .A2(n1895), .ZN(n1897) );
  INV_X1 U3424 ( .A(n1332), .ZN(n3222) );
  XNOR2_X1 U3425 ( .A(n1966), .B(n2026), .ZN(n1971) );
  NAND2_X4 U3426 ( .A1(net295737), .A2(net295738), .ZN(net295626) );
  NAND3_X2 U3427 ( .A1(net295757), .A2(net295755), .A3(net295750), .ZN(
        net295506) );
  NAND2_X4 U3428 ( .A1(n2060), .A2(n2057), .ZN(n1976) );
  NOR2_X4 U3429 ( .A1(n3036), .A2(n3159), .ZN(n3047) );
  NAND3_X2 U3430 ( .A1(n2495), .A2(net298909), .A3(n2494), .ZN(n2423) );
  INV_X8 U3431 ( .A(n2061), .ZN(n2133) );
  NAND4_X2 U3432 ( .A1(net296932), .A2(net294188), .A3(a[5]), .A4(a[4]), .ZN(
        n2118) );
  NAND2_X4 U3433 ( .A1(n3654), .A2(n3653), .ZN(n3748) );
  NAND2_X4 U3434 ( .A1(n3743), .A2(n3742), .ZN(net294770) );
  NAND2_X4 U3435 ( .A1(n2666), .A2(n2665), .ZN(n2903) );
  NAND2_X4 U3437 ( .A1(n1676), .A2(n1898), .ZN(n2055) );
  NAND2_X4 U3438 ( .A1(n3093), .A2(n3092), .ZN(n3282) );
  NAND2_X4 U3439 ( .A1(n2991), .A2(n2990), .ZN(n3092) );
  NAND2_X2 U3440 ( .A1(n3026), .A2(n1373), .ZN(n2511) );
  OAI21_X2 U3441 ( .B1(n2470), .B2(n2469), .A(n2567), .ZN(n2476) );
  NAND2_X1 U3442 ( .A1(n2226), .A2(n1561), .ZN(n2124) );
  NAND2_X4 U3443 ( .A1(n2694), .A2(n2423), .ZN(n2496) );
  NAND3_X2 U3444 ( .A1(n3452), .A2(n3451), .A3(n3450), .ZN(n3453) );
  NOR2_X2 U3447 ( .A1(n4036), .A2(n4038), .ZN(n4031) );
  NAND2_X2 U3448 ( .A1(n2953), .A2(n3052), .ZN(n2973) );
  NAND2_X4 U3449 ( .A1(n3022), .A2(n2971), .ZN(n2972) );
  NAND2_X4 U3450 ( .A1(n3328), .A2(n3327), .ZN(n3333) );
  NAND2_X4 U3451 ( .A1(n1958), .A2(n2100), .ZN(n2053) );
  NAND2_X4 U3452 ( .A1(n2768), .A2(n2769), .ZN(n2944) );
  NAND2_X4 U3453 ( .A1(net294241), .A2(n3981), .ZN(n4037) );
  NAND2_X4 U3454 ( .A1(n2202), .A2(n2201), .ZN(n2322) );
  XNOR2_X1 U3455 ( .A(n4107), .B(n4106), .ZN(n4102) );
  OAI211_X4 U3456 ( .C1(n2255), .C2(n2398), .A(n2396), .B(n2397), .ZN(n2516)
         );
  NAND2_X4 U3457 ( .A1(n1547), .A2(n3666), .ZN(net294448) );
  NAND2_X4 U3458 ( .A1(n2417), .A2(n2427), .ZN(n2424) );
  OAI221_X4 U3459 ( .B1(net294285), .B2(n3948), .C1(net294285), .C2(n3947), 
        .A(n3946), .ZN(n3964) );
  INV_X8 U3460 ( .A(net294171), .ZN(net294285) );
  NAND2_X4 U3461 ( .A1(n3901), .A2(net294299), .ZN(net294156) );
  NAND2_X4 U3462 ( .A1(n3899), .A2(n3900), .ZN(net294299) );
  NAND2_X1 U3464 ( .A1(n3483), .A2(n3343), .ZN(n3344) );
  NAND2_X4 U3465 ( .A1(n3492), .A2(n3491), .ZN(n3496) );
  INV_X4 U3466 ( .A(n3458), .ZN(n1797) );
  INV_X8 U3467 ( .A(n1797), .ZN(n1798) );
  NAND2_X4 U3468 ( .A1(n3980), .A2(n4033), .ZN(n4034) );
  NAND3_X2 U3469 ( .A1(n2327), .A2(n2069), .A3(n2068), .ZN(n2232) );
  NAND2_X4 U3470 ( .A1(n2066), .A2(n1268), .ZN(n2327) );
  NAND2_X4 U3471 ( .A1(n3021), .A2(n2980), .ZN(n3034) );
  OAI221_X4 U3472 ( .B1(n3677), .B2(net294772), .C1(n3676), .C2(n3675), .A(
        n3674), .ZN(n3745) );
  OAI22_X4 U3473 ( .A1(net297276), .A2(net296909), .B1(net296910), .B2(
        net296911), .ZN(n2194) );
  NAND2_X4 U3474 ( .A1(n2358), .A2(n2359), .ZN(n2661) );
  NOR2_X2 U3475 ( .A1(n1989), .A2(n2111), .ZN(n1992) );
  NAND2_X4 U3476 ( .A1(n2063), .A2(n2062), .ZN(n2324) );
  AOI21_X4 U3477 ( .B1(n2567), .B2(n2470), .A(n1191), .ZN(n1799) );
  NAND2_X1 U3478 ( .A1(a[8]), .A2(net297230), .ZN(n2569) );
  OAI21_X2 U3479 ( .B1(n3605), .B2(n3604), .A(n3532), .ZN(n3742) );
  NAND2_X4 U3480 ( .A1(n1591), .A2(n2683), .ZN(n2756) );
  NOR2_X2 U3481 ( .A1(n2948), .A2(n2980), .ZN(n2953) );
  AOI21_X2 U3482 ( .B1(n2672), .B2(n2671), .A(n1374), .ZN(n2674) );
  INV_X4 U3484 ( .A(n2338), .ZN(n1803) );
  NAND2_X4 U3485 ( .A1(n3063), .A2(n3064), .ZN(n3249) );
  XNOR2_X2 U3486 ( .A(n3062), .B(n3139), .ZN(n3132) );
  NOR3_X2 U3487 ( .A1(n3130), .A2(n3071), .A3(n3072), .ZN(n3075) );
  NAND2_X4 U3488 ( .A1(n2252), .A2(n2253), .ZN(n2400) );
  INV_X4 U3489 ( .A(n2693), .ZN(n2955) );
  INV_X8 U3490 ( .A(n2800), .ZN(n2936) );
  NAND2_X4 U3491 ( .A1(n3336), .A2(n3393), .ZN(n3394) );
  NAND3_X2 U3492 ( .A1(n3127), .A2(n3312), .A3(n3128), .ZN(n3074) );
  NAND2_X4 U3493 ( .A1(n3245), .A2(n3401), .ZN(n3317) );
  OAI21_X2 U3494 ( .B1(n3405), .B2(n1254), .A(n4291), .ZN(n3408) );
  NAND2_X4 U3495 ( .A1(n2022), .A2(n2023), .ZN(n2046) );
  INV_X8 U3496 ( .A(n1540), .ZN(n3260) );
  INV_X1 U3497 ( .A(n3729), .ZN(n3730) );
  NAND2_X4 U3498 ( .A1(n2950), .A2(n2946), .ZN(n3049) );
  NAND2_X4 U3500 ( .A1(n2785), .A2(n2943), .ZN(n2950) );
  NAND2_X4 U3501 ( .A1(n2432), .A2(n1378), .ZN(n2570) );
  NAND2_X1 U3502 ( .A1(n3715), .A2(n1608), .ZN(n3719) );
  OAI211_X4 U3503 ( .C1(n3642), .C2(net294048), .A(n3641), .B(n3640), .ZN(
        n3710) );
  AOI21_X2 U3504 ( .B1(n2734), .B2(n2735), .A(n1688), .ZN(n2736) );
  NAND2_X2 U3505 ( .A1(n1294), .A2(n2498), .ZN(n1802) );
  NAND2_X4 U3506 ( .A1(n3265), .A2(n3266), .ZN(n3477) );
  NAND3_X2 U3507 ( .A1(n2413), .A2(n2237), .A3(n2335), .ZN(n2238) );
  NAND3_X2 U3508 ( .A1(n3334), .A2(n3257), .A3(n3327), .ZN(n3164) );
  NAND2_X4 U3509 ( .A1(n3163), .A2(n3334), .ZN(n3335) );
  NAND2_X4 U3510 ( .A1(n3329), .A2(n3330), .ZN(n3393) );
  NAND2_X4 U3511 ( .A1(n1532), .A2(n3099), .ZN(n3008) );
  NAND2_X4 U3512 ( .A1(n3664), .A2(n3665), .ZN(n3801) );
  NAND2_X4 U3513 ( .A1(n2727), .A2(n3194), .ZN(n2818) );
  NAND2_X4 U3514 ( .A1(n3736), .A2(n3737), .ZN(n3799) );
  NAND2_X4 U3515 ( .A1(n1617), .A2(n3060), .ZN(n3142) );
  NAND2_X4 U3516 ( .A1(n2130), .A2(n2129), .ZN(n2295) );
  NAND2_X4 U3517 ( .A1(n1254), .A2(n4291), .ZN(n3519) );
  NAND2_X4 U3518 ( .A1(n2965), .A2(n3144), .ZN(n3138) );
  NAND3_X2 U3519 ( .A1(n3459), .A2(n1550), .A3(n3460), .ZN(n3274) );
  NAND2_X4 U3521 ( .A1(n1271), .A2(n3070), .ZN(n3231) );
  NAND2_X4 U3522 ( .A1(n2444), .A2(n2443), .ZN(n2521) );
  NAND2_X4 U3523 ( .A1(n2346), .A2(n2345), .ZN(n2405) );
  NAND2_X4 U3524 ( .A1(n2646), .A2(n1612), .ZN(n2817) );
  AOI22_X4 U3526 ( .A1(n2636), .A2(n2648), .B1(n2648), .B2(net297188), .ZN(
        n2637) );
  INV_X2 U3527 ( .A(net294310), .ZN(net294305) );
  NAND2_X4 U3528 ( .A1(n2059), .A2(n1578), .ZN(n2061) );
  NAND2_X4 U3529 ( .A1(n3306), .A2(n3374), .ZN(n3493) );
  NAND2_X2 U3530 ( .A1(n1932), .A2(n1931), .ZN(n1844) );
  NAND2_X4 U3531 ( .A1(n2840), .A2(n2845), .ZN(n3037) );
  NAND2_X4 U3532 ( .A1(n3477), .A2(n3502), .ZN(n3503) );
  NAND2_X4 U3533 ( .A1(n3767), .A2(net294388), .ZN(net294307) );
  NAND2_X4 U3534 ( .A1(n3902), .A2(net294394), .ZN(net294393) );
  NAND2_X1 U3535 ( .A1(n2747), .A2(n2703), .ZN(n2577) );
  NAND2_X4 U3536 ( .A1(n2550), .A2(n2643), .ZN(n2644) );
  NAND2_X4 U3537 ( .A1(n2548), .A2(n2549), .ZN(n2643) );
  NAND2_X4 U3538 ( .A1(n2546), .A2(n2547), .ZN(n2550) );
  NAND2_X4 U3539 ( .A1(n2449), .A2(n2450), .ZN(n2651) );
  OAI22_X4 U3540 ( .A1(net297278), .A2(n3922), .B1(n3221), .B2(net297188), 
        .ZN(n2548) );
  NAND3_X2 U3541 ( .A1(n2058), .A2(n1567), .A3(n1558), .ZN(n2014) );
  NAND2_X1 U3542 ( .A1(n3604), .A2(n3603), .ZN(n3533) );
  NAND2_X4 U3543 ( .A1(net295271), .A2(n3320), .ZN(n3518) );
  NAND3_X2 U3544 ( .A1(n1629), .A2(n2408), .A3(n4263), .ZN(n2409) );
  NAND2_X4 U3545 ( .A1(n3834), .A2(n3835), .ZN(n3916) );
  OAI211_X4 U3546 ( .C1(n3841), .C2(n3840), .A(n3839), .B(n3838), .ZN(n3848)
         );
  INV_X8 U3547 ( .A(n2562), .ZN(n2742) );
  NAND2_X4 U3548 ( .A1(n2882), .A2(n2883), .ZN(n3125) );
  NAND2_X4 U3549 ( .A1(n2989), .A2(n2988), .ZN(n3283) );
  NAND3_X1 U3550 ( .A1(net297640), .A2(b[18]), .A3(control[0]), .ZN(n1819) );
  NAND4_X1 U3551 ( .A1(b[17]), .A2(control[0]), .A3(a[4]), .A4(net297172), 
        .ZN(n1912) );
  INV_X8 U3552 ( .A(net299325), .ZN(net297168) );
  NAND2_X1 U3553 ( .A1(n1826), .A2(n1107), .ZN(n1828) );
  NAND2_X4 U3554 ( .A1(n2611), .A2(n2750), .ZN(n2751) );
  NAND2_X4 U3555 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND3_X2 U3556 ( .A1(n2186), .A2(n2188), .A3(n2187), .ZN(n2396) );
  NAND2_X4 U3557 ( .A1(n1216), .A2(n2104), .ZN(n2305) );
  NAND2_X4 U3558 ( .A1(n2670), .A2(n3028), .ZN(n2615) );
  NAND2_X4 U3559 ( .A1(n2509), .A2(n2508), .ZN(n3028) );
  NAND2_X4 U3560 ( .A1(n3566), .A2(n4293), .ZN(n3702) );
  NAND2_X4 U3561 ( .A1(n1631), .A2(n2510), .ZN(n2670) );
  NOR3_X2 U3562 ( .A1(n2203), .A2(net296672), .A3(n2211), .ZN(n2210) );
  NAND2_X4 U3563 ( .A1(n2349), .A2(n2350), .ZN(n2517) );
  NAND2_X4 U3564 ( .A1(n1351), .A2(n2143), .ZN(n2287) );
  NAND2_X4 U3565 ( .A1(n1497), .A2(n3080), .ZN(n3490) );
  NAND2_X4 U3566 ( .A1(n3997), .A2(net294194), .ZN(n4085) );
  NAND2_X4 U3567 ( .A1(n3985), .A2(n3984), .ZN(n4098) );
  NOR2_X4 U3568 ( .A1(n1801), .A2(n2954), .ZN(n3055) );
  NAND2_X4 U3569 ( .A1(n2598), .A2(n2597), .ZN(n2956) );
  INV_X8 U3570 ( .A(n2599), .ZN(n2598) );
  NAND3_X2 U3572 ( .A1(n2246), .A2(n1163), .A3(n1602), .ZN(n2247) );
  OAI211_X4 U3573 ( .C1(n2753), .C2(n1712), .A(n2790), .B(n2855), .ZN(n2974)
         );
  NOR2_X4 U3574 ( .A1(n1363), .A2(n3720), .ZN(n3709) );
  NAND2_X4 U3575 ( .A1(n2229), .A2(n2228), .ZN(n2413) );
  NAND2_X4 U3576 ( .A1(n2806), .A2(n1264), .ZN(n3124) );
  NAND3_X2 U3577 ( .A1(n2058), .A2(n1567), .A3(n1558), .ZN(n2134) );
  NAND2_X4 U3578 ( .A1(n3836), .A2(n1570), .ZN(n3874) );
  NAND2_X4 U3579 ( .A1(n3833), .A2(n3772), .ZN(n3836) );
  NAND2_X4 U3580 ( .A1(n1353), .A2(n3553), .ZN(n3554) );
  NAND2_X4 U3581 ( .A1(n2439), .A2(n2440), .ZN(n2669) );
  NAND2_X4 U3582 ( .A1(n2843), .A2(n2844), .ZN(n2935) );
  NAND2_X4 U3583 ( .A1(n1582), .A2(n3033), .ZN(n3161) );
  NAND2_X4 U3584 ( .A1(n2425), .A2(n2407), .ZN(n2759) );
  NAND3_X2 U3585 ( .A1(n3385), .A2(n1559), .A3(n3386), .ZN(n3232) );
  NAND2_X4 U3588 ( .A1(n1308), .A2(n2081), .ZN(n2278) );
  NAND3_X2 U3590 ( .A1(n2739), .A2(n2902), .A3(n2740), .ZN(n2830) );
  NAND2_X4 U3591 ( .A1(n1214), .A2(n1947), .ZN(n2057) );
  NAND3_X2 U3592 ( .A1(n3904), .A2(n1344), .A3(n3903), .ZN(net294333) );
  NAND2_X4 U3593 ( .A1(n1510), .A2(n2607), .ZN(n2747) );
  NAND2_X1 U3594 ( .A1(n2323), .A2(n1556), .ZN(n2064) );
  NAND2_X4 U3595 ( .A1(n3371), .A2(n3370), .ZN(n3488) );
  NAND2_X4 U3596 ( .A1(n2905), .A2(n2904), .ZN(n2914) );
  NAND2_X4 U3597 ( .A1(n2761), .A2(n1229), .ZN(n2693) );
  NAND2_X4 U3598 ( .A1(n2219), .A2(n2218), .ZN(n2412) );
  NAND2_X4 U3599 ( .A1(n2208), .A2(n2207), .ZN(n2218) );
  NAND3_X2 U3600 ( .A1(n3391), .A2(n1540), .A3(n3392), .ZN(n3510) );
  NAND2_X4 U3601 ( .A1(n3611), .A2(n3610), .ZN(net294696) );
  NAND2_X4 U3602 ( .A1(n2737), .A2(n2736), .ZN(n2992) );
  NAND2_X4 U3603 ( .A1(n2007), .A2(n2006), .ZN(n2059) );
  OAI21_X4 U3605 ( .B1(n2848), .B2(n1546), .A(n2847), .ZN(n2938) );
  OAI21_X4 U3606 ( .B1(n3261), .B2(n3262), .A(n1535), .ZN(n3263) );
  NAND2_X4 U3607 ( .A1(n4201), .A2(net296524), .ZN(n2688) );
  NAND2_X4 U3608 ( .A1(n2474), .A2(n2475), .ZN(n2702) );
  INV_X8 U3609 ( .A(n2471), .ZN(n2700) );
  XNOR2_X2 U3610 ( .A(n3722), .B(n4265), .ZN(n3723) );
  NAND2_X4 U3611 ( .A1(n1519), .A2(n3680), .ZN(n3737) );
  INV_X8 U3612 ( .A(n3247), .ZN(n3136) );
  NAND2_X4 U3613 ( .A1(n2145), .A2(n2146), .ZN(n2285) );
  NAND2_X4 U3614 ( .A1(n1544), .A2(n2672), .ZN(n2800) );
  NAND2_X4 U3615 ( .A1(n2416), .A2(n2415), .ZN(n2427) );
  OAI21_X4 U3616 ( .B1(n3398), .B2(n3399), .A(n3397), .ZN(n3414) );
  NAND2_X4 U3617 ( .A1(n3682), .A2(n3683), .ZN(n3734) );
  NAND2_X4 U3618 ( .A1(n3530), .A2(n3529), .ZN(net294844) );
  NAND2_X4 U3619 ( .A1(n3526), .A2(net294913), .ZN(net294911) );
  NAND2_X4 U3620 ( .A1(n2442), .A2(n2614), .ZN(n3026) );
  NAND2_X2 U3621 ( .A1(n2438), .A2(n2437), .ZN(n2614) );
  NAND2_X4 U3622 ( .A1(n1359), .A2(n2715), .ZN(n2993) );
  NAND2_X4 U3623 ( .A1(n3851), .A2(n3850), .ZN(net293933) );
  NAND2_X4 U3624 ( .A1(net294510), .A2(net298857), .ZN(n3798) );
  AOI21_X2 U3625 ( .B1(n3689), .B2(n4215), .A(n3688), .ZN(n3690) );
  NAND2_X1 U3626 ( .A1(n2335), .A2(n2334), .ZN(n2319) );
  NAND2_X1 U3627 ( .A1(n2291), .A2(n2334), .ZN(n2297) );
  NAND2_X4 U3628 ( .A1(n2334), .A2(n2335), .ZN(n2489) );
  NAND2_X1 U3629 ( .A1(n3453), .A2(n3439), .ZN(n3356) );
  INV_X8 U3630 ( .A(n3032), .ZN(n2798) );
  NAND2_X4 U3631 ( .A1(n2670), .A2(n2669), .ZN(n3032) );
  NAND2_X4 U3632 ( .A1(net294045), .A2(net298969), .ZN(net294196) );
  NAND2_X1 U3633 ( .A1(n3034), .A2(n3035), .ZN(n2981) );
  NAND3_X4 U3634 ( .A1(net297616), .A2(n1984), .A3(n1713), .ZN(n2116) );
  NAND2_X4 U3635 ( .A1(n1838), .A2(n1837), .ZN(n1932) );
  NAND2_X4 U3636 ( .A1(n3734), .A2(n1162), .ZN(net294309) );
  NAND2_X1 U3637 ( .A1(n3768), .A2(net294322), .ZN(n3932) );
  OAI22_X4 U3638 ( .A1(n1862), .A2(n1861), .B1(net297086), .B2(n1860), .ZN(
        n1917) );
  NAND2_X4 U3639 ( .A1(n2749), .A2(n2748), .ZN(n2789) );
  NAND2_X4 U3640 ( .A1(n1633), .A2(n3268), .ZN(n3502) );
  OAI22_X4 U3641 ( .A1(b[17]), .A2(net297180), .B1(b[25]), .B2(control[0]), 
        .ZN(n1863) );
  NAND2_X4 U3642 ( .A1(n3424), .A2(n3564), .ZN(n3631) );
  OAI22_X4 U3643 ( .A1(n1865), .A2(n1866), .B1(n1864), .B2(n1863), .ZN(n1916)
         );
  XNOR2_X2 U3644 ( .A(n3342), .B(n3482), .ZN(n3343) );
  OAI21_X2 U3645 ( .B1(n3786), .B2(n1678), .A(net294100), .ZN(n3787) );
  NAND3_X1 U3646 ( .A1(n2577), .A2(n2672), .A3(n2609), .ZN(n2606) );
  NAND3_X2 U3647 ( .A1(n3452), .A2(n3451), .A3(n3450), .ZN(n3855) );
  NAND2_X1 U3648 ( .A1(n2534), .A2(n2651), .ZN(n2535) );
  NAND2_X1 U3649 ( .A1(a[30]), .A2(net297485), .ZN(n4004) );
  NAND2_X1 U3650 ( .A1(a[28]), .A2(net297485), .ZN(n3881) );
  NAND2_X1 U3651 ( .A1(a[26]), .A2(net297485), .ZN(n3752) );
  NAND2_X1 U3652 ( .A1(a[24]), .A2(net297485), .ZN(n3586) );
  NAND2_X1 U3653 ( .A1(a[22]), .A2(net297485), .ZN(net295168) );
  NAND2_X1 U3654 ( .A1(a[20]), .A2(net297485), .ZN(net295387) );
  NAND2_X1 U3655 ( .A1(a[18]), .A2(net297485), .ZN(net295624) );
  NAND3_X2 U3656 ( .A1(n2054), .A2(n2055), .A3(n1567), .ZN(n2015) );
  AOI22_X4 U3658 ( .A1(n1531), .A2(n3872), .B1(net293933), .B2(n1548), .ZN(
        n3930) );
  INV_X8 U3659 ( .A(n3046), .ZN(n3160) );
  OAI22_X4 U3660 ( .A1(b[17]), .A2(net297184), .B1(b[25]), .B2(control[0]), 
        .ZN(n1833) );
  NAND2_X4 U3661 ( .A1(n1664), .A2(n1693), .ZN(n2949) );
  NAND2_X4 U3662 ( .A1(n1376), .A2(n3172), .ZN(n3374) );
  NAND2_X4 U3663 ( .A1(n2799), .A2(n2839), .ZN(n2845) );
  OAI22_X4 U3664 ( .A1(b[16]), .A2(net298225), .B1(b[24]), .B2(control[0]), 
        .ZN(n1829) );
  NAND2_X4 U3665 ( .A1(net296430), .A2(n2418), .ZN(net296418) );
  NAND3_X4 U3666 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3595) );
  NAND3_X2 U3667 ( .A1(n3517), .A2(n3518), .A3(n3516), .ZN(n3521) );
  NAND2_X4 U3669 ( .A1(n3905), .A2(n4215), .ZN(net294308) );
  NAND2_X1 U3671 ( .A1(n3464), .A2(n3459), .ZN(n3462) );
  NAND2_X4 U3672 ( .A1(n3118), .A2(n3117), .ZN(n3312) );
  NAND2_X4 U3673 ( .A1(n2442), .A2(n2614), .ZN(n2797) );
  NOR2_X2 U3674 ( .A1(n3787), .A2(n3795), .ZN(n3797) );
  NAND2_X4 U3675 ( .A1(n3321), .A2(n3518), .ZN(n3403) );
  NAND3_X2 U3676 ( .A1(n2418), .A2(n2327), .A3(n2419), .ZN(n2585) );
  NAND3_X2 U3677 ( .A1(n4057), .A2(n4058), .A3(n4059), .ZN(n4065) );
  INV_X2 U3678 ( .A(n1520), .ZN(n4051) );
  NAND2_X4 U3680 ( .A1(n2725), .A2(n2726), .ZN(n3194) );
  NAND3_X1 U3681 ( .A1(n1965), .A2(n1964), .A3(n2053), .ZN(n2047) );
  NAND2_X4 U3682 ( .A1(n1787), .A2(n4061), .ZN(n3853) );
  NAND2_X4 U3683 ( .A1(net294701), .A2(n3909), .ZN(n3910) );
  NAND2_X4 U3684 ( .A1(n2106), .A2(net296788), .ZN(net296326) );
  NAND2_X4 U3685 ( .A1(n2244), .A2(n2245), .ZN(n2482) );
  NAND2_X4 U3686 ( .A1(n3580), .A2(net294940), .ZN(n3672) );
  NAND2_X4 U3687 ( .A1(n3709), .A2(n3721), .ZN(n3873) );
  NAND3_X2 U3688 ( .A1(n2866), .A2(n2687), .A3(n1160), .ZN(n2583) );
  NAND2_X4 U3689 ( .A1(n2695), .A2(n2696), .ZN(n2866) );
  NAND2_X4 U3690 ( .A1(n3416), .A2(n3415), .ZN(n3538) );
  NAND2_X4 U3691 ( .A1(n3911), .A2(net294701), .ZN(net294321) );
  NAND3_X2 U3692 ( .A1(n1514), .A2(n3578), .A3(n3577), .ZN(net294994) );
  NAND3_X2 U3693 ( .A1(n3385), .A2(n1108), .A3(n3386), .ZN(n3579) );
  NAND2_X1 U3694 ( .A1(n2426), .A2(n1160), .ZN(n2428) );
  NAND2_X1 U3695 ( .A1(n2687), .A2(n1629), .ZN(n2497) );
  NAND2_X4 U3696 ( .A1(n3728), .A2(n3729), .ZN(n3911) );
  NAND3_X1 U3697 ( .A1(n3483), .A2(n1124), .A3(n3481), .ZN(n3486) );
  NAND2_X4 U3698 ( .A1(n3341), .A2(net294779), .ZN(n3482) );
  NAND3_X2 U3699 ( .A1(n3335), .A2(n1154), .A3(n3392), .ZN(n3509) );
  NAND2_X1 U3700 ( .A1(n2754), .A2(n2974), .ZN(n2787) );
  NAND2_X4 U3701 ( .A1(n2952), .A2(n2974), .ZN(n3052) );
  NAND2_X1 U3702 ( .A1(n2578), .A2(n2866), .ZN(n2502) );
  NAND2_X1 U3703 ( .A1(n2686), .A2(n2689), .ZN(n2578) );
  NAND2_X4 U3704 ( .A1(control[1]), .A2(net298225), .ZN(net294048) );
  INV_X32 U3705 ( .A(control[0]), .ZN(net297180) );
  NAND3_X4 U3707 ( .A1(control[0]), .A2(control[1]), .A3(b[0]), .ZN(n1804) );
  INV_X4 U3708 ( .A(n1804), .ZN(n1805) );
  NOR2_X4 U3709 ( .A1(n1805), .A2(n1785), .ZN(net297061) );
  INV_X4 U3710 ( .A(n3618), .ZN(n1806) );
  MUX2_X2 U3711 ( .A(\set_product_in_sig/z1 [0]), .B(n1806), .S(net297196), 
        .Z(product_out[0]) );
  INV_X4 U3712 ( .A(a[0]), .ZN(n1807) );
  INV_X4 U3713 ( .A(a[1]), .ZN(n1810) );
  XNOR2_X2 U3714 ( .A(n1809), .B(n1808), .ZN(n2268) );
  INV_X4 U3715 ( .A(n2268), .ZN(n3639) );
  MUX2_X2 U3716 ( .A(\set_product_in_sig/z1 [1]), .B(n3639), .S(net297196), 
        .Z(product_out[1]) );
  NOR2_X4 U3717 ( .A1(net296771), .A2(n1810), .ZN(n1812) );
  NAND2_X2 U3719 ( .A1(a[0]), .A2(control[1]), .ZN(n1816) );
  NAND2_X2 U3720 ( .A1(a[0]), .A2(net297172), .ZN(n1814) );
  OAI22_X2 U3721 ( .A1(n1816), .A2(n1815), .B1(n1814), .B2(n1813), .ZN(n1839)
         );
  NAND3_X2 U3722 ( .A1(net297281), .A2(a[1]), .A3(n1839), .ZN(n1931) );
  XNOR2_X2 U3723 ( .A(n1818), .B(n1817), .ZN(n1827) );
  INV_X4 U3724 ( .A(b[26]), .ZN(n1821) );
  INV_X4 U3725 ( .A(n1822), .ZN(n1823) );
  NOR3_X4 U3726 ( .A1(n1825), .A2(n1824), .A3(n1823), .ZN(net297128) );
  NAND2_X2 U3727 ( .A1(a[0]), .A2(net297262), .ZN(n1826) );
  INV_X4 U3728 ( .A(n1826), .ZN(n1856) );
  NAND2_X2 U3729 ( .A1(a[1]), .A2(control[1]), .ZN(n1832) );
  NAND2_X2 U3730 ( .A1(a[1]), .A2(n1380), .ZN(n1830) );
  NAND2_X2 U3731 ( .A1(a[2]), .A2(control[1]), .ZN(n1836) );
  NAND3_X2 U3732 ( .A1(net297481), .A2(a[1]), .A3(n1839), .ZN(n1984) );
  INV_X4 U3733 ( .A(n1844), .ZN(n1842) );
  INV_X4 U3734 ( .A(n1859), .ZN(n1845) );
  NAND2_X2 U3735 ( .A1(a[1]), .A2(net294175), .ZN(n1847) );
  OAI21_X4 U3736 ( .B1(n1846), .B2(n1845), .A(n1847), .ZN(n1898) );
  INV_X4 U3737 ( .A(n1847), .ZN(n1857) );
  XNOR2_X2 U3738 ( .A(n1849), .B(n1850), .ZN(n1852) );
  NAND2_X2 U3739 ( .A1(a[0]), .A2(net297226), .ZN(n1851) );
  INV_X4 U3740 ( .A(n1851), .ZN(n1853) );
  NAND2_X2 U3741 ( .A1(n1854), .A2(n1950), .ZN(n3825) );
  INV_X4 U3742 ( .A(n3825), .ZN(n2464) );
  MUX2_X2 U3743 ( .A(\set_product_in_sig/z1 [3]), .B(n2464), .S(net297196), 
        .Z(product_out[3]) );
  NAND2_X2 U3744 ( .A1(a[3]), .A2(control[1]), .ZN(n1862) );
  OAI22_X2 U3745 ( .A1(b[0]), .A2(net297180), .B1(b[8]), .B2(control[0]), .ZN(
        n1861) );
  NAND2_X2 U3746 ( .A1(a[2]), .A2(control[1]), .ZN(n1866) );
  OAI22_X2 U3747 ( .A1(b[1]), .A2(net298226), .B1(b[9]), .B2(control[0]), .ZN(
        n1865) );
  NAND2_X2 U3748 ( .A1(a[2]), .A2(net297640), .ZN(n1864) );
  INV_X4 U3749 ( .A(n1878), .ZN(n1875) );
  XNOR2_X2 U3750 ( .A(n1877), .B(n1876), .ZN(n2056) );
  NAND2_X2 U3751 ( .A1(a[2]), .A2(net297262), .ZN(n2008) );
  NAND3_X2 U3752 ( .A1(net294188), .A2(net296932), .A3(n1284), .ZN(n2196) );
  XNOR2_X2 U3754 ( .A(n1883), .B(n1884), .ZN(n2012) );
  XNOR2_X2 U3755 ( .A(n1886), .B(n1182), .ZN(n1887) );
  INV_X4 U3756 ( .A(n1952), .ZN(n1889) );
  NAND2_X2 U3757 ( .A1(b[12]), .A2(net294515), .ZN(n1893) );
  NAND2_X2 U3758 ( .A1(b[4]), .A2(net297196), .ZN(n1892) );
  AOI22_X2 U3759 ( .A1(b[28]), .A2(net294051), .B1(b[20]), .B2(net294053), 
        .ZN(n1891) );
  NAND2_X2 U3760 ( .A1(a[0]), .A2(net297244), .ZN(n1894) );
  INV_X4 U3761 ( .A(n1894), .ZN(n1896) );
  INV_X4 U3762 ( .A(n3922), .ZN(n3219) );
  MUX2_X2 U3763 ( .A(\set_product_in_sig/z1 [4]), .B(n3219), .S(net297196), 
        .Z(product_out[4]) );
  INV_X4 U3764 ( .A(n2055), .ZN(n1899) );
  NOR2_X4 U3765 ( .A1(n1899), .A2(n1951), .ZN(n1901) );
  INV_X4 U3766 ( .A(n2008), .ZN(n2013) );
  OAI21_X4 U3767 ( .B1(n1901), .B2(n1182), .A(n1953), .ZN(n1977) );
  NAND2_X2 U3768 ( .A1(b[16]), .A2(control[0]), .ZN(n1902) );
  INV_X4 U3769 ( .A(n1902), .ZN(n1998) );
  NAND2_X2 U3770 ( .A1(n1998), .A2(n1903), .ZN(n1909) );
  NAND2_X2 U3771 ( .A1(b[0]), .A2(control[1]), .ZN(n1994) );
  NOR2_X4 U3772 ( .A1(net297182), .A2(net296909), .ZN(n1904) );
  NAND2_X2 U3773 ( .A1(n1995), .A2(n1904), .ZN(n1908) );
  NAND2_X2 U3774 ( .A1(b[8]), .A2(control[1]), .ZN(n1996) );
  INV_X4 U3775 ( .A(n1996), .ZN(n1906) );
  NOR2_X4 U3776 ( .A1(control[0]), .A2(net296909), .ZN(n1905) );
  NAND2_X2 U3777 ( .A1(n1906), .A2(n1905), .ZN(n1907) );
  NOR2_X4 U3778 ( .A1(n1922), .A2(n1921), .ZN(n1929) );
  NOR2_X4 U3779 ( .A1(n1926), .A2(n1925), .ZN(n1927) );
  NAND3_X4 U3780 ( .A1(n1929), .A2(n4213), .A3(n1927), .ZN(n2115) );
  OAI21_X4 U3781 ( .B1(n1936), .B2(n1935), .A(n1941), .ZN(n2060) );
  INV_X4 U3782 ( .A(n1941), .ZN(n1943) );
  XNOR2_X2 U3784 ( .A(n1976), .B(n1975), .ZN(n1948) );
  XNOR2_X2 U3785 ( .A(n1948), .B(n1977), .ZN(n2100) );
  XNOR2_X2 U3786 ( .A(n1955), .B(n1956), .ZN(n1957) );
  OAI21_X4 U3787 ( .B1(n2097), .B2(n2098), .A(n2096), .ZN(n1958) );
  INV_X4 U3788 ( .A(n1965), .ZN(n1961) );
  NAND2_X2 U3789 ( .A1(a[1]), .A2(net297246), .ZN(n1963) );
  OAI21_X4 U3790 ( .B1(n1962), .B2(n1961), .A(n1963), .ZN(n2027) );
  INV_X4 U3791 ( .A(n1963), .ZN(n1964) );
  NAND2_X2 U3792 ( .A1(n1574), .A2(n2047), .ZN(n1966) );
  NAND2_X2 U3793 ( .A1(b[13]), .A2(net294515), .ZN(n1969) );
  NAND2_X2 U3794 ( .A1(b[5]), .A2(net297196), .ZN(n1968) );
  AOI22_X2 U3795 ( .A1(b[29]), .A2(net294051), .B1(b[21]), .B2(net294053), 
        .ZN(n1967) );
  NAND2_X2 U3796 ( .A1(a[0]), .A2(net297216), .ZN(n1970) );
  NAND2_X2 U3797 ( .A1(n1971), .A2(n1970), .ZN(n1974) );
  INV_X4 U3798 ( .A(n1970), .ZN(n1973) );
  INV_X4 U3799 ( .A(n1971), .ZN(n1972) );
  NAND2_X2 U3800 ( .A1(n1973), .A2(n1972), .ZN(n2043) );
  INV_X4 U3801 ( .A(n3994), .ZN(n3295) );
  MUX2_X2 U3802 ( .A(\set_product_in_sig/z1 [5]), .B(n3295), .S(net297196), 
        .Z(product_out[5]) );
  NAND2_X2 U3803 ( .A1(a[1]), .A2(net297218), .ZN(n2032) );
  NAND2_X2 U3804 ( .A1(a[2]), .A2(net297246), .ZN(n2023) );
  INV_X4 U3805 ( .A(n1975), .ZN(n1979) );
  INV_X4 U3806 ( .A(n2020), .ZN(n2019) );
  AOI21_X4 U3809 ( .B1(n1991), .B2(n1992), .A(n1990), .ZN(n2004) );
  NAND2_X2 U3810 ( .A1(a[5]), .A2(net297515), .ZN(n1993) );
  INV_X4 U3811 ( .A(n1993), .ZN(n2063) );
  INV_X4 U3812 ( .A(n1994), .ZN(n1995) );
  NAND2_X2 U3813 ( .A1(a[6]), .A2(net299325), .ZN(n1997) );
  INV_X4 U3814 ( .A(n1997), .ZN(n1999) );
  NAND2_X2 U3815 ( .A1(n1999), .A2(n1998), .ZN(n2000) );
  NAND4_X2 U3816 ( .A1(n2003), .A2(n2002), .A3(n2001), .A4(n2000), .ZN(n2062)
         );
  NAND2_X2 U3817 ( .A1(n2063), .A2(n2062), .ZN(n2107) );
  INV_X4 U3818 ( .A(a[6]), .ZN(net296911) );
  NAND2_X2 U3819 ( .A1(a[4]), .A2(net297260), .ZN(n2006) );
  NAND3_X4 U3820 ( .A1(n2015), .A2(n1759), .A3(n2014), .ZN(n2016) );
  XNOR2_X2 U3821 ( .A(n2016), .B(n2017), .ZN(n2021) );
  INV_X4 U3822 ( .A(n2024), .ZN(n2022) );
  INV_X4 U3823 ( .A(n2023), .ZN(n2025) );
  NAND2_X2 U3824 ( .A1(n2025), .A2(n2024), .ZN(n2049) );
  XNOR2_X2 U3825 ( .A(n2030), .B(n2029), .ZN(n2033) );
  NAND3_X2 U3826 ( .A1(a[1]), .A2(n2033), .A3(net297216), .ZN(n2177) );
  NAND2_X2 U3827 ( .A1(n2044), .A2(n2177), .ZN(n2034) );
  XNOR2_X2 U3828 ( .A(n2034), .B(n2043), .ZN(n2039) );
  NAND2_X2 U3829 ( .A1(b[14]), .A2(net294515), .ZN(n2037) );
  NAND2_X2 U3830 ( .A1(b[6]), .A2(net297196), .ZN(n2036) );
  AOI22_X2 U3831 ( .A1(b[30]), .A2(net294051), .B1(b[22]), .B2(net294053), 
        .ZN(n2035) );
  NAND2_X2 U3832 ( .A1(a[0]), .A2(net297202), .ZN(n2038) );
  NAND2_X2 U3833 ( .A1(n2039), .A2(n2038), .ZN(n2042) );
  INV_X4 U3834 ( .A(n2038), .ZN(n2041) );
  INV_X4 U3835 ( .A(n2039), .ZN(n2040) );
  NAND2_X2 U3836 ( .A1(n2042), .A2(n2161), .ZN(n4049) );
  INV_X4 U3837 ( .A(n4049), .ZN(n3359) );
  MUX2_X2 U3838 ( .A(\set_product_in_sig/z1 [6]), .B(n3359), .S(net297196), 
        .Z(product_out[6]) );
  INV_X4 U3839 ( .A(n2043), .ZN(n2045) );
  INV_X4 U3840 ( .A(n2084), .ZN(n2152) );
  INV_X4 U3841 ( .A(n2029), .ZN(n2050) );
  OAI21_X4 U3842 ( .B1(n2051), .B2(n2050), .A(n2049), .ZN(n2190) );
  NAND2_X2 U3843 ( .A1(a[2]), .A2(net297218), .ZN(n2052) );
  NAND2_X2 U3844 ( .A1(a[3]), .A2(net297246), .ZN(n2081) );
  INV_X4 U3845 ( .A(n2081), .ZN(n2093) );
  NAND3_X4 U3846 ( .A1(n2135), .A2(n2133), .A3(n2134), .ZN(n2334) );
  NAND2_X2 U3847 ( .A1(a[5]), .A2(net297260), .ZN(n2230) );
  INV_X4 U3848 ( .A(n2324), .ZN(n2113) );
  NOR3_X4 U3849 ( .A1(n2071), .A2(n2113), .A3(n2198), .ZN(n2231) );
  INV_X4 U3850 ( .A(n2327), .ZN(n2206) );
  NAND3_X2 U3851 ( .A1(n2072), .A2(n2233), .A3(n2232), .ZN(n2131) );
  XNOR2_X2 U3852 ( .A(n2073), .B(n2076), .ZN(n2304) );
  INV_X4 U3853 ( .A(n2304), .ZN(n2095) );
  NAND2_X2 U3854 ( .A1(a[4]), .A2(net297230), .ZN(n2094) );
  INV_X4 U3855 ( .A(n2094), .ZN(n2302) );
  XNOR2_X2 U3856 ( .A(n2074), .B(n2075), .ZN(n2279) );
  XNOR2_X2 U3857 ( .A(n2078), .B(n2077), .ZN(n2478) );
  INV_X4 U3859 ( .A(n2089), .ZN(n2086) );
  INV_X4 U3860 ( .A(n2090), .ZN(n2085) );
  NAND2_X2 U3861 ( .A1(a[1]), .A2(net297202), .ZN(n2087) );
  OAI21_X4 U3862 ( .B1(n2086), .B2(n2085), .A(n2087), .ZN(n2159) );
  INV_X4 U3863 ( .A(n2087), .ZN(n2088) );
  NAND3_X2 U3864 ( .A1(n2090), .A2(n2089), .A3(n2088), .ZN(n2160) );
  NAND2_X2 U3865 ( .A1(n2159), .A2(n2160), .ZN(n2091) );
  XNOR2_X2 U3866 ( .A(n2091), .B(n2161), .ZN(n2092) );
  INV_X4 U3867 ( .A(n2092), .ZN(n2168) );
  NAND2_X2 U3868 ( .A1(b[15]), .A2(net294515), .ZN(net296808) );
  INV_X4 U3869 ( .A(net294980), .ZN(net294052) );
  MUX2_X2 U3870 ( .A(\set_product_in_sig/z1 [7]), .B(net294052), .S(net297196), 
        .Z(product_out[7]) );
  NAND2_X2 U3871 ( .A1(a[2]), .A2(net297202), .ZN(n2158) );
  INV_X4 U3872 ( .A(n2158), .ZN(n2155) );
  INV_X4 U3873 ( .A(n2149), .ZN(n2191) );
  NAND2_X2 U3874 ( .A1(a[4]), .A2(net297246), .ZN(n2146) );
  INV_X4 U3875 ( .A(n2146), .ZN(n2143) );
  NAND2_X2 U3876 ( .A1(n2095), .A2(n2094), .ZN(n2105) );
  NAND2_X2 U3877 ( .A1(n2110), .A2(n2109), .ZN(n2222) );
  NOR2_X4 U3878 ( .A1(n2113), .A2(net296781), .ZN(n2119) );
  NAND2_X2 U3879 ( .A1(a[6]), .A2(net294175), .ZN(n2226) );
  INV_X4 U3880 ( .A(a[7]), .ZN(n2121) );
  INV_X4 U3881 ( .A(n2122), .ZN(n2201) );
  OAI21_X4 U3882 ( .B1(n2202), .B2(n2123), .A(n2322), .ZN(n2225) );
  XNOR2_X2 U3883 ( .A(n2125), .B(n2124), .ZN(n2130) );
  INV_X4 U3884 ( .A(n2226), .ZN(n2229) );
  XNOR2_X2 U3885 ( .A(n2128), .B(n2127), .ZN(n2129) );
  INV_X4 U3886 ( .A(n2132), .ZN(n2291) );
  INV_X4 U3887 ( .A(n2316), .ZN(n2137) );
  NAND2_X2 U3888 ( .A1(a[5]), .A2(net297230), .ZN(n2298) );
  INV_X4 U3889 ( .A(n2298), .ZN(n2296) );
  XNOR2_X2 U3890 ( .A(n2142), .B(n2141), .ZN(n2144) );
  INV_X4 U3891 ( .A(n2144), .ZN(n2145) );
  XNOR2_X2 U3892 ( .A(n2147), .B(n2178), .ZN(n2174) );
  INV_X4 U3893 ( .A(n2180), .ZN(n2175) );
  OAI22_X2 U3894 ( .A1(n2148), .A2(n2180), .B1(n2175), .B2(n2174), .ZN(n2154)
         );
  XNOR2_X2 U3895 ( .A(n2154), .B(n2153), .ZN(n2156) );
  INV_X4 U3896 ( .A(n2156), .ZN(n2157) );
  INV_X4 U3897 ( .A(n2159), .ZN(n2162) );
  OAI21_X4 U3898 ( .B1(n2162), .B2(n2161), .A(n2160), .ZN(n2172) );
  XNOR2_X2 U3899 ( .A(n2163), .B(n2172), .ZN(n2166) );
  INV_X4 U3900 ( .A(n2166), .ZN(n2164) );
  NAND2_X2 U3901 ( .A1(a[1]), .A2(net297254), .ZN(n2165) );
  INV_X4 U3902 ( .A(n2165), .ZN(n2167) );
  NAND2_X2 U3903 ( .A1(n1289), .A2(n2168), .ZN(n2263) );
  XNOR2_X2 U3904 ( .A(n2169), .B(n2263), .ZN(n2895) );
  OAI22_X2 U3905 ( .A1(net297279), .A2(n3618), .B1(n2895), .B2(net297188), 
        .ZN(n2171) );
  INV_X4 U3906 ( .A(n2171), .ZN(n2170) );
  XNOR2_X2 U3907 ( .A(n2170), .B(n1286), .ZN(product_out[8]) );
  NAND2_X2 U3908 ( .A1(n1286), .A2(n2171), .ZN(n2389) );
  INV_X4 U3909 ( .A(n2389), .ZN(n2274) );
  NAND2_X2 U3910 ( .A1(\set_product_in_sig/z1 [9]), .A2(net297188), .ZN(n2271)
         );
  INV_X4 U3911 ( .A(n2271), .ZN(n2269) );
  NAND2_X2 U3912 ( .A1(a[2]), .A2(net297254), .ZN(n2373) );
  NAND2_X2 U3913 ( .A1(n2175), .A2(n2174), .ZN(n2397) );
  INV_X4 U3914 ( .A(n2178), .ZN(n2179) );
  AOI21_X4 U3915 ( .B1(n2189), .B2(n1493), .A(n2401), .ZN(n2193) );
  INV_X4 U3916 ( .A(n2218), .ZN(n2209) );
  NAND2_X2 U3917 ( .A1(a[7]), .A2(net297260), .ZN(n2213) );
  OAI21_X4 U3918 ( .B1(n2210), .B2(n2209), .A(n2213), .ZN(n2760) );
  INV_X4 U3919 ( .A(n2211), .ZN(n2212) );
  INV_X4 U3920 ( .A(n2213), .ZN(n2214) );
  NAND4_X2 U3921 ( .A1(n2221), .A2(n2222), .A3(n2223), .A4(n2220), .ZN(n2224)
         );
  INV_X4 U3922 ( .A(n2227), .ZN(n2228) );
  XNOR2_X2 U3923 ( .A(n2241), .B(n2408), .ZN(n2243) );
  NAND2_X2 U3924 ( .A1(a[6]), .A2(net297230), .ZN(n2242) );
  INV_X4 U3925 ( .A(n2242), .ZN(n2245) );
  INV_X4 U3926 ( .A(n2243), .ZN(n2244) );
  NAND2_X2 U3928 ( .A1(a[5]), .A2(net297244), .ZN(n2250) );
  XNOR2_X2 U3929 ( .A(n2254), .B(n2288), .ZN(n2395) );
  INV_X4 U3931 ( .A(n2398), .ZN(n2256) );
  XNOR2_X2 U3932 ( .A(n2355), .B(n2257), .ZN(n2260) );
  NAND2_X2 U3933 ( .A1(a[3]), .A2(net297202), .ZN(n2259) );
  INV_X4 U3934 ( .A(n2259), .ZN(n2261) );
  NAND2_X2 U3935 ( .A1(n2261), .A2(n2260), .ZN(n2277) );
  NAND2_X2 U3936 ( .A1(n2527), .A2(n2277), .ZN(n2374) );
  XNOR2_X2 U3937 ( .A(n2262), .B(n2374), .ZN(n2267) );
  INV_X4 U3938 ( .A(n2263), .ZN(n2265) );
  XNOR2_X2 U3939 ( .A(n2267), .B(n2266), .ZN(n3637) );
  NAND2_X2 U3940 ( .A1(n2269), .A2(n2270), .ZN(n2388) );
  INV_X4 U3941 ( .A(n2270), .ZN(n2272) );
  NAND2_X2 U3942 ( .A1(n2272), .A2(n2271), .ZN(n2387) );
  NAND2_X2 U3943 ( .A1(n2388), .A2(n2387), .ZN(n2273) );
  XNOR2_X2 U3944 ( .A(n2274), .B(n2273), .ZN(product_out[9]) );
  NAND3_X4 U3945 ( .A1(n2277), .A2(n1296), .A3(n2275), .ZN(n2528) );
  NAND2_X2 U3946 ( .A1(a[5]), .A2(net297216), .ZN(n2351) );
  INV_X4 U3947 ( .A(n2351), .ZN(n2350) );
  NAND3_X2 U3948 ( .A1(n2286), .A2(n1493), .A3(n2284), .ZN(n2402) );
  NAND2_X2 U3949 ( .A1(a[6]), .A2(net297244), .ZN(n2345) );
  INV_X4 U3950 ( .A(n2345), .ZN(n2343) );
  XNOR2_X2 U3951 ( .A(n2294), .B(n2293), .ZN(n2310) );
  XOR2_X2 U3952 ( .A(n2299), .B(n2300), .Z(n2309) );
  NOR2_X4 U3953 ( .A1(n2302), .A2(n2303), .ZN(n2308) );
  INV_X4 U3954 ( .A(n2337), .ZN(n2432) );
  NAND2_X2 U3955 ( .A1(n2338), .A2(n2491), .ZN(n2318) );
  INV_X4 U3956 ( .A(n2320), .ZN(n2321) );
  NAND3_X4 U3957 ( .A1(n2323), .A2(n1556), .A3(net296544), .ZN(n2325) );
  OAI21_X4 U3958 ( .B1(n2326), .B2(net296547), .A(n2325), .ZN(n2331) );
  NAND2_X2 U3959 ( .A1(a[8]), .A2(net297260), .ZN(net296529) );
  INV_X4 U3960 ( .A(net296529), .ZN(net296524) );
  INV_X4 U3961 ( .A(net296536), .ZN(net296535) );
  XNOR2_X2 U3962 ( .A(n2330), .B(net296535), .ZN(n2425) );
  NOR2_X4 U3963 ( .A1(n2331), .A2(n2332), .ZN(net296530) );
  OAI21_X4 U3965 ( .B1(n2432), .B2(n1378), .A(n2341), .ZN(n2472) );
  NAND2_X2 U3966 ( .A1(n2343), .A2(n2344), .ZN(n2467) );
  INV_X4 U3967 ( .A(n1619), .ZN(n2349) );
  INV_X4 U3968 ( .A(n2352), .ZN(n2357) );
  INV_X4 U3969 ( .A(n2353), .ZN(n2354) );
  XNOR2_X2 U3970 ( .A(n2356), .B(n2357), .ZN(n2360) );
  INV_X4 U3971 ( .A(n2360), .ZN(n2358) );
  NAND2_X2 U3972 ( .A1(a[4]), .A2(net297202), .ZN(n2359) );
  INV_X4 U3973 ( .A(n2359), .ZN(n2361) );
  NAND2_X2 U3975 ( .A1(a[3]), .A2(net297254), .ZN(n2363) );
  INV_X4 U3976 ( .A(n2363), .ZN(n2366) );
  NAND2_X2 U3977 ( .A1(n2459), .A2(n2460), .ZN(n2381) );
  INV_X4 U3978 ( .A(n2368), .ZN(n2369) );
  INV_X4 U3979 ( .A(n2374), .ZN(n2372) );
  XNOR2_X2 U3980 ( .A(n2375), .B(n2373), .ZN(n2371) );
  XNOR2_X2 U3981 ( .A(n2371), .B(n2372), .ZN(n2379) );
  INV_X4 U3982 ( .A(n2373), .ZN(n2377) );
  XNOR2_X2 U3983 ( .A(n2375), .B(n2374), .ZN(n2376) );
  NAND2_X2 U3984 ( .A1(n2377), .A2(n2376), .ZN(n2378) );
  OAI21_X4 U3985 ( .B1(n2380), .B2(n2379), .A(n2378), .ZN(n2458) );
  INV_X4 U3986 ( .A(n2384), .ZN(n2382) );
  NAND2_X2 U3987 ( .A1(\set_product_in_sig/z1 [10]), .A2(net297188), .ZN(n2383) );
  INV_X4 U3988 ( .A(n2383), .ZN(n2385) );
  INV_X4 U3989 ( .A(n2387), .ZN(n2390) );
  OAI21_X4 U3990 ( .B1(n2390), .B2(n2389), .A(n2388), .ZN(n2391) );
  XNOR2_X2 U3991 ( .A(n2393), .B(n2391), .ZN(product_out[10]) );
  INV_X4 U3992 ( .A(n2391), .ZN(n2394) );
  OAI21_X4 U3993 ( .B1(n2394), .B2(n2393), .A(n2392), .ZN(n2641) );
  NAND2_X2 U3994 ( .A1(\set_product_in_sig/z1 [11]), .A2(net297188), .ZN(n2639) );
  NAND2_X2 U3995 ( .A1(a[6]), .A2(net297216), .ZN(n2443) );
  INV_X4 U3996 ( .A(n2443), .ZN(n2557) );
  NAND3_X2 U3997 ( .A1(n2406), .A2(n2405), .A3(n2404), .ZN(n2468) );
  INV_X4 U3998 ( .A(n2569), .ZN(n2470) );
  AOI21_X4 U3999 ( .B1(n2425), .B2(n2407), .A(n2414), .ZN(n2411) );
  INV_X4 U4000 ( .A(n2409), .ZN(n2410) );
  NOR2_X4 U4001 ( .A1(n2411), .A2(n2410), .ZN(n2417) );
  NAND2_X2 U4003 ( .A1(a[9]), .A2(net297260), .ZN(n2422) );
  OAI21_X4 U4004 ( .B1(n2421), .B2(net296416), .A(n2422), .ZN(n2694) );
  INV_X4 U4005 ( .A(n2422), .ZN(n2494) );
  NAND2_X2 U4006 ( .A1(n2429), .A2(n2470), .ZN(n2430) );
  XNOR2_X2 U4007 ( .A(n2431), .B(n2430), .ZN(n2567) );
  XNOR2_X2 U4008 ( .A(n2436), .B(n2476), .ZN(n2438) );
  NAND2_X2 U4009 ( .A1(a[7]), .A2(net297244), .ZN(n2437) );
  INV_X4 U4010 ( .A(n2437), .ZN(n2440) );
  NAND2_X2 U4011 ( .A1(n2521), .A2(n2558), .ZN(n2445) );
  XNOR2_X2 U4012 ( .A(n2445), .B(n2446), .ZN(n2449) );
  NAND2_X2 U4013 ( .A1(a[5]), .A2(net297202), .ZN(n2448) );
  INV_X4 U4014 ( .A(n2448), .ZN(n2450) );
  INV_X4 U4015 ( .A(n2455), .ZN(n2453) );
  NAND2_X2 U4016 ( .A1(a[4]), .A2(net297254), .ZN(n2454) );
  INV_X4 U4017 ( .A(n2454), .ZN(n2456) );
  INV_X4 U4018 ( .A(n2459), .ZN(n2461) );
  NAND2_X2 U4019 ( .A1(n2464), .A2(net294515), .ZN(n2465) );
  OAI21_X4 U4020 ( .B1(n3824), .B2(net297188), .A(n2465), .ZN(n2638) );
  XNOR2_X2 U4021 ( .A(n2639), .B(n2638), .ZN(n2552) );
  XNOR2_X2 U4022 ( .A(n2466), .B(n2552), .ZN(product_out[11]) );
  NAND2_X2 U4023 ( .A1(a[5]), .A2(net297254), .ZN(n2539) );
  INV_X4 U4024 ( .A(n2539), .ZN(n2532) );
  INV_X4 U4025 ( .A(n2654), .ZN(n2655) );
  NAND2_X2 U4026 ( .A1(a[7]), .A2(net297216), .ZN(n2563) );
  OAI21_X4 U4027 ( .B1(n2485), .B2(n2484), .A(n2483), .ZN(n2701) );
  NAND2_X2 U4028 ( .A1(a[9]), .A2(net297230), .ZN(n2504) );
  INV_X4 U4029 ( .A(n2504), .ZN(n2574) );
  INV_X4 U4030 ( .A(n2489), .ZN(n2492) );
  OAI21_X4 U4031 ( .B1(n2492), .B2(n4273), .A(n2338), .ZN(n2758) );
  NAND2_X2 U4032 ( .A1(a[11]), .A2(net297272), .ZN(net296334) );
  NAND2_X2 U4033 ( .A1(net295990), .A2(net295754), .ZN(n2593) );
  NAND2_X2 U4034 ( .A1(net296430), .A2(net295991), .ZN(n2498) );
  INV_X4 U4035 ( .A(n2586), .ZN(n2499) );
  XNOR2_X2 U4036 ( .A(n2593), .B(n2501), .ZN(n2686) );
  NAND2_X2 U4037 ( .A1(a[10]), .A2(net297260), .ZN(n2689) );
  INV_X4 U4038 ( .A(n2689), .ZN(n2696) );
  INV_X4 U4039 ( .A(n2686), .ZN(n2695) );
  XNOR2_X2 U4040 ( .A(n2503), .B(n2502), .ZN(n2505) );
  XNOR2_X2 U4041 ( .A(n2507), .B(n2506), .ZN(n2509) );
  NAND2_X2 U4042 ( .A1(a[8]), .A2(net297244), .ZN(n2508) );
  INV_X4 U4043 ( .A(n2508), .ZN(n2510) );
  XNOR2_X2 U4044 ( .A(n2511), .B(n2615), .ZN(n2564) );
  INV_X4 U4045 ( .A(n2564), .ZN(n2512) );
  XOR2_X2 U4047 ( .A(n2514), .B(n2513), .Z(n2652) );
  OAI21_X4 U4048 ( .B1(n2518), .B2(n4257), .A(n2517), .ZN(n2520) );
  OAI21_X4 U4049 ( .B1(n2522), .B2(n4259), .A(n2558), .ZN(n2656) );
  INV_X4 U4050 ( .A(n2656), .ZN(n2523) );
  XNOR2_X2 U4051 ( .A(n2524), .B(n2523), .ZN(n2525) );
  XNOR2_X2 U4053 ( .A(n2630), .B(n2533), .ZN(n2531) );
  XNOR2_X2 U4054 ( .A(n2538), .B(n1758), .ZN(n2540) );
  INV_X4 U4055 ( .A(n2541), .ZN(n2544) );
  OAI21_X4 U4056 ( .B1(n2544), .B2(n2543), .A(n2542), .ZN(n2633) );
  XNOR2_X2 U4057 ( .A(n2633), .B(n2545), .ZN(n3924) );
  INV_X4 U4058 ( .A(n3924), .ZN(n3221) );
  INV_X4 U4059 ( .A(n2548), .ZN(n2546) );
  NAND2_X2 U4060 ( .A1(\set_product_in_sig/z1 [12]), .A2(net297188), .ZN(n2547) );
  INV_X4 U4061 ( .A(n2547), .ZN(n2549) );
  INV_X4 U4062 ( .A(n2639), .ZN(n2551) );
  XNOR2_X2 U4063 ( .A(n2554), .B(n2553), .ZN(product_out[12]) );
  NAND2_X2 U4064 ( .A1(n3295), .A2(net294515), .ZN(n2648) );
  OAI21_X4 U4065 ( .B1(n1651), .B2(n2559), .A(n2558), .ZN(n2561) );
  INV_X4 U4066 ( .A(n2563), .ZN(n2565) );
  INV_X4 U4067 ( .A(n2566), .ZN(n2741) );
  NOR2_X4 U4068 ( .A1(n2742), .A2(n2741), .ZN(n2918) );
  INV_X4 U4069 ( .A(n2570), .ZN(n2572) );
  NAND2_X2 U4070 ( .A1(n2574), .A2(n2573), .ZN(n2575) );
  NAND2_X2 U4071 ( .A1(a[9]), .A2(net297244), .ZN(n2613) );
  INV_X4 U4072 ( .A(n2613), .ZN(n2672) );
  NAND3_X2 U4073 ( .A1(net295748), .A2(net297526), .A3(net295754), .ZN(
        net296230) );
  INV_X4 U4074 ( .A(net296230), .ZN(net296222) );
  NAND2_X2 U4075 ( .A1(a[12]), .A2(net297272), .ZN(n2587) );
  INV_X4 U4076 ( .A(n2587), .ZN(n2678) );
  INV_X4 U4077 ( .A(n2679), .ZN(n2592) );
  OAI21_X4 U4078 ( .B1(net296106), .B2(net296216), .A(n2592), .ZN(n2595) );
  NAND3_X4 U4079 ( .A1(n2596), .A2(n2595), .A3(n2594), .ZN(n2599) );
  NAND2_X2 U4080 ( .A1(a[11]), .A2(net297260), .ZN(n2600) );
  INV_X4 U4081 ( .A(n2600), .ZN(n2597) );
  NAND2_X2 U4082 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  NAND2_X2 U4083 ( .A1(a[10]), .A2(net297228), .ZN(n2603) );
  INV_X4 U4084 ( .A(n2603), .ZN(n2604) );
  XNOR2_X2 U4085 ( .A(n2606), .B(n2605), .ZN(n2671) );
  NOR2_X4 U4086 ( .A1(n1518), .A2(n2881), .ZN(n2619) );
  INV_X4 U4087 ( .A(n2621), .ZN(n2623) );
  NOR2_X4 U4088 ( .A1(n1295), .A2(n2624), .ZN(n2632) );
  NAND2_X2 U4089 ( .A1(n2626), .A2(n2625), .ZN(n2662) );
  INV_X4 U4090 ( .A(n2627), .ZN(n2628) );
  AOI21_X4 U4091 ( .B1(n2630), .B2(n2629), .A(n2628), .ZN(n2631) );
  XNOR2_X2 U4092 ( .A(n2631), .B(n2632), .ZN(n2732) );
  XNOR2_X2 U4093 ( .A(n2635), .B(n2719), .ZN(n3992) );
  INV_X4 U4094 ( .A(n3992), .ZN(n2636) );
  NAND2_X2 U4095 ( .A1(\set_product_in_sig/z1 [13]), .A2(net297188), .ZN(n2647) );
  INV_X4 U4096 ( .A(n2638), .ZN(n2640) );
  NAND2_X2 U4097 ( .A1(n2640), .A2(n2639), .ZN(n2642) );
  AOI21_X4 U4098 ( .B1(n2642), .B2(n2641), .A(n1272), .ZN(n2645) );
  OAI21_X4 U4099 ( .B1(n2645), .B2(n2644), .A(n4247), .ZN(n2646) );
  INV_X4 U4100 ( .A(n2647), .ZN(n2650) );
  INV_X4 U4101 ( .A(n2648), .ZN(n2649) );
  NAND2_X2 U4102 ( .A1(n2650), .A2(n2649), .ZN(n2816) );
  NAND2_X2 U4103 ( .A1(a[7]), .A2(net297254), .ZN(n2716) );
  INV_X4 U4104 ( .A(n2716), .ZN(n2715) );
  XNOR2_X2 U4105 ( .A(n2658), .B(n2657), .ZN(n2659) );
  NOR2_X4 U4106 ( .A1(n2936), .A2(n3028), .ZN(n2673) );
  OAI21_X4 U4107 ( .B1(n2848), .B2(n2676), .A(n2675), .ZN(n2710) );
  NAND2_X2 U4108 ( .A1(a[11]), .A2(net297228), .ZN(n2850) );
  INV_X4 U4109 ( .A(n2850), .ZN(n2699) );
  NAND2_X2 U4110 ( .A1(a[12]), .A2(net297260), .ZN(n2684) );
  INV_X4 U4111 ( .A(n2684), .ZN(n2683) );
  INV_X4 U4112 ( .A(net296106), .ZN(net296105) );
  NAND3_X2 U4113 ( .A1(net296104), .A2(net295749), .A3(net296105), .ZN(n2681)
         );
  NAND2_X2 U4114 ( .A1(a[13]), .A2(net297272), .ZN(net296098) );
  NAND2_X2 U4115 ( .A1(net295755), .A2(net296097), .ZN(n2773) );
  NOR2_X4 U4116 ( .A1(n2955), .A2(n2764), .ZN(n2697) );
  OAI21_X4 U4117 ( .B1(n2702), .B2(n2701), .A(n2700), .ZN(n2748) );
  INV_X4 U4118 ( .A(n2748), .ZN(n2704) );
  NAND2_X2 U4119 ( .A1(n2751), .A2(n1573), .ZN(n2857) );
  XNOR2_X2 U4121 ( .A(n1311), .B(n2709), .ZN(n2837) );
  OAI21_X4 U4122 ( .B1(n2839), .B2(n2799), .A(n2837), .ZN(n2801) );
  XNOR2_X2 U4123 ( .A(n4198), .B(n2801), .ZN(n2915) );
  NAND2_X2 U4124 ( .A1(a[9]), .A2(net297216), .ZN(n2916) );
  INV_X4 U4125 ( .A(n2916), .ZN(n2883) );
  XNOR2_X2 U4126 ( .A(n2712), .B(n2711), .ZN(n2907) );
  XNOR2_X2 U4127 ( .A(n2722), .B(n4253), .ZN(n4048) );
  NAND2_X2 U4128 ( .A1(\set_product_in_sig/z1 [14]), .A2(net297188), .ZN(n2724) );
  INV_X4 U4129 ( .A(n2724), .ZN(n2726) );
  NAND2_X2 U4130 ( .A1(\set_product_in_sig/z1 [15]), .A2(net297188), .ZN(n3195) );
  INV_X4 U4131 ( .A(n3195), .ZN(n2815) );
  INV_X4 U4132 ( .A(n2730), .ZN(n2731) );
  NAND2_X2 U4133 ( .A1(a[8]), .A2(net297254), .ZN(n2813) );
  INV_X4 U4134 ( .A(n2813), .ZN(n2827) );
  NAND2_X2 U4135 ( .A1(a[9]), .A2(net297202), .ZN(n2901) );
  OAI211_X2 U4136 ( .C1(n2745), .C2(n2744), .A(n3125), .B(n2743), .ZN(n2808)
         );
  NAND2_X2 U4137 ( .A1(a[11]), .A2(net297244), .ZN(n2795) );
  INV_X4 U4138 ( .A(n2756), .ZN(n2862) );
  NAND3_X2 U4139 ( .A1(net297526), .A2(net295749), .A3(net295754), .ZN(
        net295996) );
  INV_X4 U4140 ( .A(net295749), .ZN(net295983) );
  NOR2_X4 U4141 ( .A1(net295991), .A2(n2770), .ZN(n2772) );
  INV_X4 U4142 ( .A(net295990), .ZN(net295989) );
  NOR3_X4 U4143 ( .A1(n2772), .A2(n2771), .A3(net295989), .ZN(n2775) );
  INV_X4 U4144 ( .A(n2773), .ZN(n2774) );
  OAI21_X4 U4145 ( .B1(net295983), .B2(n2775), .A(n2774), .ZN(net295757) );
  OAI21_X4 U4146 ( .B1(net295982), .B2(net295757), .A(net295755), .ZN(n2777)
         );
  INV_X4 U4148 ( .A(net295756), .ZN(net295978) );
  NAND2_X2 U4149 ( .A1(a[13]), .A2(net297260), .ZN(n2780) );
  OAI21_X4 U4150 ( .B1(n2779), .B2(n2778), .A(n2780), .ZN(n2861) );
  INV_X4 U4151 ( .A(n2780), .ZN(n2781) );
  NAND2_X2 U4152 ( .A1(a[12]), .A2(net297228), .ZN(n2784) );
  INV_X4 U4153 ( .A(n2784), .ZN(n2943) );
  INV_X4 U4154 ( .A(n2795), .ZN(n2844) );
  XNOR2_X2 U4155 ( .A(n2787), .B(n2786), .ZN(n3039) );
  NAND2_X2 U4156 ( .A1(n2842), .A2(n2795), .ZN(n3038) );
  NAND2_X2 U4157 ( .A1(n3039), .A2(n3038), .ZN(n2796) );
  INV_X4 U4158 ( .A(n2796), .ZN(n2841) );
  NAND2_X2 U4159 ( .A1(n3028), .A2(n3027), .ZN(n2846) );
  AOI21_X4 U4160 ( .B1(n2804), .B2(n2803), .A(n2802), .ZN(n2805) );
  XNOR2_X2 U4161 ( .A(n2805), .B(n1776), .ZN(n2806) );
  XNOR2_X2 U4162 ( .A(n2808), .B(n2807), .ZN(n2809) );
  INV_X4 U4163 ( .A(n2809), .ZN(n2900) );
  NAND2_X2 U4164 ( .A1(n2901), .A2(n2900), .ZN(n2811) );
  INV_X4 U4165 ( .A(n2901), .ZN(n2810) );
  XNOR2_X2 U4166 ( .A(n2826), .B(n2828), .ZN(net294054) );
  INV_X4 U4167 ( .A(n2816), .ZN(n2821) );
  OAI21_X4 U4168 ( .B1(n2820), .B2(n2821), .A(n2819), .ZN(n3192) );
  OAI21_X4 U4169 ( .B1(n2832), .B2(n2831), .A(n2913), .ZN(n3009) );
  NAND2_X2 U4170 ( .A1(a[10]), .A2(net297202), .ZN(n2892) );
  INV_X4 U4171 ( .A(n2892), .ZN(n2889) );
  INV_X4 U4172 ( .A(n2857), .ZN(n2834) );
  XNOR2_X2 U4173 ( .A(n2836), .B(n1679), .ZN(n2838) );
  NAND2_X2 U4174 ( .A1(n2933), .A2(n1301), .ZN(n2925) );
  INV_X4 U4175 ( .A(n2846), .ZN(n2847) );
  NAND2_X2 U4176 ( .A1(a[12]), .A2(net297244), .ZN(n3023) );
  INV_X4 U4177 ( .A(n3023), .ZN(n2877) );
  AOI21_X4 U4178 ( .B1(n2853), .B2(n2852), .A(n2851), .ZN(n2860) );
  INV_X4 U4179 ( .A(n2854), .ZN(n2856) );
  NAND4_X2 U4180 ( .A1(n1338), .A2(n2857), .A3(n2856), .A4(n2855), .ZN(n2859)
         );
  INV_X4 U4181 ( .A(n2942), .ZN(n2865) );
  NAND2_X2 U4182 ( .A1(a[14]), .A2(net297260), .ZN(n2872) );
  INV_X4 U4183 ( .A(n2872), .ZN(n2963) );
  NAND2_X2 U4184 ( .A1(a[13]), .A2(net297228), .ZN(n2951) );
  INV_X4 U4185 ( .A(n2951), .ZN(n2874) );
  XNOR2_X2 U4186 ( .A(n2876), .B(n2875), .ZN(n2878) );
  NAND2_X2 U4187 ( .A1(a[11]), .A2(net297216), .ZN(n2922) );
  OAI21_X4 U4188 ( .B1(n2883), .B2(n2882), .A(n2881), .ZN(n3126) );
  XNOR2_X2 U4189 ( .A(n2888), .B(n2887), .ZN(n2890) );
  NAND2_X2 U4190 ( .A1(a[9]), .A2(net297254), .ZN(n2994) );
  XNOR2_X2 U4191 ( .A(n3008), .B(n2994), .ZN(n2893) );
  XNOR2_X2 U4192 ( .A(n2893), .B(n3009), .ZN(n3012) );
  XNOR2_X2 U4193 ( .A(n2894), .B(n1621), .ZN(n3617) );
  INV_X4 U4194 ( .A(n2895), .ZN(n3615) );
  OAI21_X4 U4195 ( .B1(n1600), .B2(net297188), .A(n2897), .ZN(n3200) );
  NAND2_X2 U4196 ( .A1(\set_product_in_sig/z1 [16]), .A2(net297188), .ZN(n3201) );
  XNOR2_X2 U4197 ( .A(n3200), .B(n3201), .ZN(n3002) );
  NAND2_X2 U4198 ( .A1(\set_product_in_sig/z1 [17]), .A2(net297188), .ZN(n3207) );
  INV_X4 U4199 ( .A(n3207), .ZN(n3005) );
  NAND2_X2 U4200 ( .A1(net294053), .A2(n3639), .ZN(n2899) );
  OAI21_X4 U4201 ( .B1(n3637), .B2(net297279), .A(n2899), .ZN(n3203) );
  NAND2_X2 U4202 ( .A1(n3005), .A2(n3203), .ZN(n3000) );
  NAND2_X2 U4203 ( .A1(a[10]), .A2(net297254), .ZN(n2990) );
  INV_X4 U4204 ( .A(n2990), .ZN(n2988) );
  INV_X4 U4205 ( .A(n2903), .ZN(n2904) );
  NAND3_X4 U4206 ( .A1(n2912), .A2(n2914), .A3(n2913), .ZN(n3367) );
  NAND3_X4 U4207 ( .A1(n1532), .A2(n3367), .A3(n3369), .ZN(n3103) );
  NAND2_X2 U4208 ( .A1(n2882), .A2(n2917), .ZN(n2920) );
  AOI21_X4 U4209 ( .B1(n2920), .B2(n2919), .A(n2918), .ZN(n3130) );
  XNOR2_X2 U4210 ( .A(n2927), .B(n2926), .ZN(n2928) );
  INV_X4 U4211 ( .A(n3127), .ZN(n2931) );
  INV_X4 U4212 ( .A(n2939), .ZN(n2932) );
  NAND3_X2 U4213 ( .A1(n2941), .A2(n2940), .A3(n3043), .ZN(n2982) );
  XNOR2_X2 U4214 ( .A(n2943), .B(n2942), .ZN(n2945) );
  XNOR2_X2 U4215 ( .A(n2945), .B(n2944), .ZN(n2946) );
  OAI21_X4 U4216 ( .B1(n2961), .B2(n2960), .A(n1238), .ZN(n3057) );
  INV_X4 U4217 ( .A(n3057), .ZN(n2962) );
  OAI21_X4 U4218 ( .B1(n3055), .B2(n3054), .A(n2962), .ZN(n3140) );
  NAND2_X2 U4219 ( .A1(n2963), .A2(net295759), .ZN(n3141) );
  NAND2_X2 U4220 ( .A1(a[15]), .A2(net297260), .ZN(n2964) );
  OAI21_X4 U4221 ( .B1(net295733), .B2(net295734), .A(n2964), .ZN(n2965) );
  XNOR2_X2 U4222 ( .A(n2966), .B(n3138), .ZN(n2969) );
  NAND2_X2 U4223 ( .A1(a[14]), .A2(net297228), .ZN(n2968) );
  INV_X4 U4224 ( .A(n2968), .ZN(n2970) );
  XNOR2_X2 U4225 ( .A(n2973), .B(n2972), .ZN(n3035) );
  XNOR2_X2 U4226 ( .A(n2979), .B(n2978), .ZN(n3021) );
  XNOR2_X2 U4227 ( .A(n2982), .B(n2981), .ZN(n3118) );
  INV_X4 U4228 ( .A(n3117), .ZN(n2984) );
  XNOR2_X2 U4229 ( .A(n1120), .B(n3106), .ZN(n3101) );
  NAND2_X2 U4230 ( .A1(a[11]), .A2(net297204), .ZN(n3100) );
  INV_X4 U4231 ( .A(n3100), .ZN(n3107) );
  INV_X4 U4233 ( .A(n2994), .ZN(n3010) );
  XNOR2_X2 U4234 ( .A(n3009), .B(n3008), .ZN(n2995) );
  NOR2_X4 U4235 ( .A1(n3005), .A2(n3203), .ZN(n2999) );
  NAND2_X2 U4236 ( .A1(n3000), .A2(n3215), .ZN(n3182) );
  INV_X4 U4237 ( .A(n3182), .ZN(n3004) );
  INV_X4 U4238 ( .A(n3201), .ZN(n3199) );
  NAND2_X2 U4239 ( .A1(n3199), .A2(n3200), .ZN(n3185) );
  NAND2_X2 U4241 ( .A1(n3005), .A2(n3203), .ZN(n3184) );
  OAI21_X4 U4242 ( .B1(n3006), .B2(n3182), .A(n3184), .ZN(n3087) );
  INV_X4 U4243 ( .A(n3007), .ZN(n3091) );
  NOR2_X4 U4244 ( .A1(n3011), .A2(n3091), .ZN(n3016) );
  NAND2_X2 U4245 ( .A1(n3010), .A2(n2995), .ZN(n3090) );
  OAI21_X4 U4246 ( .B1(n3011), .B2(n3280), .A(n3283), .ZN(n3015) );
  OAI21_X4 U4247 ( .B1(n3020), .B2(n3019), .A(n3018), .ZN(n3081) );
  NAND2_X2 U4248 ( .A1(a[12]), .A2(net297204), .ZN(n3080) );
  INV_X4 U4249 ( .A(n3080), .ZN(n3078) );
  INV_X4 U4250 ( .A(n3070), .ZN(n3114) );
  NOR2_X4 U4251 ( .A1(n3024), .A2(n3023), .ZN(n3025) );
  INV_X4 U4252 ( .A(n3027), .ZN(n3030) );
  NOR2_X4 U4253 ( .A1(n3030), .A2(n3029), .ZN(n3031) );
  NOR3_X4 U4254 ( .A1(n3042), .A2(n3040), .A3(n3041), .ZN(n3044) );
  OAI21_X4 U4255 ( .B1(n3044), .B2(n3045), .A(n3043), .ZN(n3046) );
  INV_X4 U4256 ( .A(n3049), .ZN(n3051) );
  OAI21_X4 U4257 ( .B1(n2947), .B2(n3051), .A(n3050), .ZN(n3053) );
  NAND3_X4 U4258 ( .A1(n3052), .A2(n1159), .A3(n3053), .ZN(n3134) );
  NOR2_X4 U4259 ( .A1(n3055), .A2(n3054), .ZN(n3056) );
  NAND2_X2 U4260 ( .A1(n3141), .A2(n3057), .ZN(n3239) );
  NAND2_X2 U4261 ( .A1(a[16]), .A2(net297260), .ZN(n3060) );
  INV_X4 U4262 ( .A(n3060), .ZN(n3061) );
  NAND2_X2 U4263 ( .A1(a[15]), .A2(net297228), .ZN(n3064) );
  INV_X4 U4264 ( .A(n3064), .ZN(n3133) );
  NAND2_X2 U4265 ( .A1(a[14]), .A2(net297244), .ZN(n3256) );
  INV_X4 U4266 ( .A(n3256), .ZN(n3068) );
  XNOR2_X2 U4267 ( .A(n3069), .B(n3335), .ZN(n3113) );
  NAND2_X2 U4268 ( .A1(n3114), .A2(n3113), .ZN(n3386) );
  XNOR2_X2 U4269 ( .A(n3085), .B(n3084), .ZN(net294611) );
  INV_X4 U4270 ( .A(n3186), .ZN(n3205) );
  NAND2_X2 U4271 ( .A1(n3205), .A2(net297188), .ZN(n3213) );
  NAND2_X2 U4272 ( .A1(\set_product_in_sig/z1 [18]), .A2(net297188), .ZN(n3204) );
  XNOR2_X2 U4273 ( .A(n3086), .B(n3204), .ZN(n3181) );
  XNOR2_X2 U4274 ( .A(n3087), .B(n1300), .ZN(product_out[18]) );
  OAI22_X2 U4275 ( .A1(net294519), .A2(n3825), .B1(n3824), .B2(net294048), 
        .ZN(n3178) );
  NAND2_X2 U4276 ( .A1(n1287), .A2(n3178), .ZN(n3439) );
  INV_X4 U4277 ( .A(n1117), .ZN(n3088) );
  INV_X4 U4279 ( .A(n3282), .ZN(n3094) );
  NAND2_X2 U4280 ( .A1(n3105), .A2(n3104), .ZN(n3111) );
  INV_X4 U4281 ( .A(n3111), .ZN(n3110) );
  OAI22_X2 U4282 ( .A1(n3112), .A2(n3111), .B1(n3110), .B2(n3109), .ZN(n3489)
         );
  OAI21_X4 U4283 ( .B1(n3308), .B2(n3307), .A(n1332), .ZN(n3174) );
  INV_X4 U4284 ( .A(n3231), .ZN(n3313) );
  INV_X4 U4285 ( .A(n3116), .ZN(n3120) );
  NAND3_X2 U4286 ( .A1(n3126), .A2(n3125), .A3(n3124), .ZN(n3129) );
  NAND3_X4 U4287 ( .A1(n3134), .A2(n3065), .A3(n4200), .ZN(n3247) );
  AOI21_X4 U4288 ( .B1(n3137), .B2(n3065), .A(n3136), .ZN(n3156) );
  OAI21_X4 U4289 ( .B1(n3145), .B2(n3144), .A(n4272), .ZN(n3235) );
  INV_X4 U4290 ( .A(net295494), .ZN(net295496) );
  NAND2_X2 U4291 ( .A1(a[17]), .A2(net297260), .ZN(n3147) );
  OAI21_X4 U4292 ( .B1(net295495), .B2(net295496), .A(n3147), .ZN(n3148) );
  NAND2_X2 U4293 ( .A1(n3148), .A2(net295393), .ZN(n3242) );
  NAND2_X2 U4294 ( .A1(a[16]), .A2(net297228), .ZN(n3151) );
  NAND2_X2 U4295 ( .A1(n3150), .A2(n3151), .ZN(n3154) );
  XNOR2_X2 U4297 ( .A(n3156), .B(n3155), .ZN(n3158) );
  NAND2_X2 U4298 ( .A1(a[15]), .A2(net297244), .ZN(n3157) );
  XNOR2_X2 U4300 ( .A(n3394), .B(n1242), .ZN(n3167) );
  NAND2_X2 U4301 ( .A1(a[14]), .A2(net297216), .ZN(n3166) );
  INV_X4 U4302 ( .A(n3166), .ZN(n3169) );
  XNOR2_X2 U4303 ( .A(n3171), .B(n3170), .ZN(n3173) );
  NAND2_X2 U4304 ( .A1(a[13]), .A2(net297204), .ZN(n3172) );
  INV_X4 U4305 ( .A(n3172), .ZN(n3224) );
  XNOR2_X2 U4306 ( .A(n3174), .B(n3493), .ZN(n3175) );
  XNOR2_X2 U4307 ( .A(n3177), .B(n3176), .ZN(n3826) );
  INV_X4 U4308 ( .A(n3204), .ZN(n3214) );
  NAND2_X2 U4309 ( .A1(n3214), .A2(n3186), .ZN(n3216) );
  INV_X4 U4310 ( .A(n3216), .ZN(n3187) );
  AOI21_X4 U4311 ( .B1(n3189), .B2(n3188), .A(n3187), .ZN(n3190) );
  XNOR2_X2 U4312 ( .A(n3190), .B(n1293), .ZN(product_out[19]) );
  NOR2_X4 U4313 ( .A1(n3192), .A2(n3193), .ZN(n3198) );
  NOR3_X4 U4314 ( .A1(n3198), .A2(n3197), .A3(n3196), .ZN(n3212) );
  INV_X4 U4316 ( .A(n3200), .ZN(n3202) );
  INV_X4 U4317 ( .A(n3203), .ZN(n3206) );
  OAI22_X2 U4318 ( .A1(n3207), .A2(n3206), .B1(n3205), .B2(n3204), .ZN(n3208)
         );
  NOR2_X4 U4319 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  OAI21_X4 U4320 ( .B1(n3212), .B2(n3211), .A(n3210), .ZN(n3452) );
  NOR2_X4 U4321 ( .A1(n3214), .A2(n3213), .ZN(n3218) );
  OAI21_X4 U4322 ( .B1(n3218), .B2(n3217), .A(n3216), .ZN(n3450) );
  NAND2_X2 U4323 ( .A1(n3219), .A2(net294053), .ZN(n3220) );
  NAND2_X2 U4324 ( .A1(\set_product_in_sig/z1 [20]), .A2(net297188), .ZN(n3352) );
  NAND2_X2 U4325 ( .A1(n3448), .A2(n3352), .ZN(n3290) );
  NAND2_X2 U4326 ( .A1(a[13]), .A2(net297254), .ZN(n3276) );
  INV_X4 U4327 ( .A(n3276), .ZN(n3464) );
  NAND2_X2 U4328 ( .A1(n3224), .A2(n3223), .ZN(n3494) );
  INV_X4 U4329 ( .A(n3232), .ZN(n3233) );
  NOR2_X4 U4330 ( .A1(n3234), .A2(n3233), .ZN(n3270) );
  NAND2_X2 U4331 ( .A1(a[17]), .A2(net297228), .ZN(n3244) );
  INV_X4 U4332 ( .A(n3242), .ZN(n3237) );
  NAND3_X4 U4333 ( .A1(n1241), .A2(n3248), .A3(n3249), .ZN(n3517) );
  XNOR2_X2 U4334 ( .A(n3250), .B(n3317), .ZN(n3253) );
  INV_X4 U4335 ( .A(n3253), .ZN(n3251) );
  NAND2_X2 U4336 ( .A1(a[16]), .A2(net297244), .ZN(n3252) );
  INV_X4 U4337 ( .A(n3252), .ZN(n3254) );
  NAND2_X2 U4338 ( .A1(n3254), .A2(n3253), .ZN(n3512) );
  NAND2_X2 U4339 ( .A1(n3507), .A2(n3512), .ZN(n3264) );
  INV_X4 U4340 ( .A(n3255), .ZN(n3262) );
  OAI21_X4 U4341 ( .B1(n3260), .B2(n3333), .A(n3336), .ZN(n3261) );
  XNOR2_X2 U4342 ( .A(n3263), .B(n3264), .ZN(n3267) );
  NAND2_X2 U4344 ( .A1(a[15]), .A2(net297216), .ZN(n3266) );
  INV_X4 U4345 ( .A(n3266), .ZN(n3268) );
  XNOR2_X2 U4346 ( .A(n3270), .B(n3577), .ZN(n3272) );
  NAND2_X2 U4347 ( .A1(a[14]), .A2(net297204), .ZN(n3271) );
  INV_X4 U4348 ( .A(n3271), .ZN(n3302) );
  XNOR2_X2 U4349 ( .A(n3274), .B(n3463), .ZN(n3275) );
  INV_X4 U4350 ( .A(n3275), .ZN(n3277) );
  NOR2_X4 U4351 ( .A1(n1772), .A2(n1504), .ZN(n3286) );
  NAND3_X4 U4352 ( .A1(n3283), .A2(n3282), .A3(n1118), .ZN(n3284) );
  NAND2_X2 U4353 ( .A1(n3352), .A2(net297190), .ZN(n3287) );
  AOI21_X2 U4354 ( .B1(n3289), .B2(n3920), .A(n3288), .ZN(n3294) );
  NAND2_X2 U4355 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  NAND2_X2 U4356 ( .A1(n3295), .A2(net294053), .ZN(n3296) );
  OAI21_X4 U4357 ( .B1(n3297), .B2(net297279), .A(n3296), .ZN(n3350) );
  NOR2_X4 U4359 ( .A1(n1255), .A2(n3311), .ZN(n3316) );
  NAND2_X2 U4360 ( .A1(a[19]), .A2(net297260), .ZN(net295277) );
  NAND2_X2 U4361 ( .A1(net295277), .A2(net295278), .ZN(net295274) );
  NAND2_X2 U4362 ( .A1(a[18]), .A2(net297228), .ZN(n3319) );
  INV_X4 U4363 ( .A(n3319), .ZN(n3320) );
  NAND2_X2 U4364 ( .A1(a[17]), .A2(net297244), .ZN(n3323) );
  NAND2_X2 U4369 ( .A1(a[15]), .A2(net297204), .ZN(n3483) );
  INV_X4 U4370 ( .A(n3483), .ZN(n3363) );
  INV_X4 U4371 ( .A(n3343), .ZN(n3362) );
  NAND2_X2 U4372 ( .A1(n3344), .A2(n3365), .ZN(n3364) );
  XNOR2_X2 U4373 ( .A(n3345), .B(n3364), .ZN(n3347) );
  NAND2_X2 U4374 ( .A1(a[14]), .A2(net297254), .ZN(n3346) );
  INV_X4 U4375 ( .A(n3346), .ZN(n3470) );
  XNOR2_X2 U4377 ( .A(n3349), .B(n3348), .ZN(n3993) );
  AOI21_X4 U4378 ( .B1(\set_product_in_sig/z1 [21]), .B2(net297188), .A(n3350), 
        .ZN(n3351) );
  INV_X4 U4379 ( .A(n3447), .ZN(n3357) );
  INV_X4 U4380 ( .A(n3352), .ZN(n3354) );
  NAND2_X2 U4381 ( .A1(n3354), .A2(n3353), .ZN(n3440) );
  INV_X4 U4382 ( .A(n3440), .ZN(n3355) );
  AOI21_X2 U4383 ( .B1(n3356), .B2(n3357), .A(n3355), .ZN(n3358) );
  XNOR2_X2 U4384 ( .A(n3358), .B(n1151), .ZN(product_out[21]) );
  NAND2_X2 U4385 ( .A1(\set_product_in_sig/z1 [22]), .A2(net297190), .ZN(n3429) );
  NAND2_X2 U4386 ( .A1(n3359), .A2(net294053), .ZN(n3360) );
  INV_X4 U4387 ( .A(n3361), .ZN(n3430) );
  NAND2_X2 U4388 ( .A1(n3430), .A2(net297190), .ZN(n3445) );
  NAND2_X2 U4389 ( .A1(n3429), .A2(n3445), .ZN(n3433) );
  NAND2_X2 U4391 ( .A1(n3364), .A2(n3571), .ZN(n3563) );
  INV_X4 U4392 ( .A(n3366), .ZN(n3497) );
  NAND3_X4 U4393 ( .A1(n3367), .A2(n3368), .A3(n3369), .ZN(n3370) );
  INV_X4 U4394 ( .A(n1360), .ZN(n3376) );
  NAND2_X2 U4395 ( .A1(n3482), .A2(n1507), .ZN(n3390) );
  OAI21_X4 U4396 ( .B1(n3384), .B2(n3383), .A(n1595), .ZN(n3578) );
  NAND3_X2 U4397 ( .A1(n4288), .A2(n3508), .A3(n3509), .ZN(n3398) );
  INV_X4 U4398 ( .A(n3512), .ZN(n3396) );
  NAND2_X2 U4401 ( .A1(n3401), .A2(n3400), .ZN(n3515) );
  NAND2_X2 U4402 ( .A1(a[19]), .A2(net297228), .ZN(n3406) );
  NAND3_X2 U4403 ( .A1(a[19]), .A2(net295156), .A3(net297226), .ZN(n3596) );
  XNOR2_X2 U4404 ( .A(n3408), .B(n3407), .ZN(n3411) );
  NAND2_X2 U4405 ( .A1(a[18]), .A2(net297244), .ZN(n3410) );
  INV_X4 U4406 ( .A(n3410), .ZN(n3412) );
  NAND2_X2 U4407 ( .A1(n3412), .A2(n3411), .ZN(n3582) );
  XNOR2_X2 U4408 ( .A(n3414), .B(n3413), .ZN(n3500) );
  XNOR2_X2 U4409 ( .A(n3417), .B(net299334), .ZN(n3485) );
  NAND2_X2 U4410 ( .A1(a[16]), .A2(net297204), .ZN(n3484) );
  INV_X4 U4411 ( .A(n3484), .ZN(n3419) );
  INV_X4 U4412 ( .A(n3485), .ZN(n3418) );
  XNOR2_X2 U4413 ( .A(n3421), .B(n3420), .ZN(n3423) );
  NAND2_X2 U4414 ( .A1(a[15]), .A2(net297254), .ZN(n3422) );
  INV_X4 U4415 ( .A(n3422), .ZN(n3564) );
  INV_X4 U4416 ( .A(n3423), .ZN(n3424) );
  NAND2_X2 U4417 ( .A1(n3631), .A2(n3630), .ZN(n4043) );
  INV_X4 U4418 ( .A(n3561), .ZN(n3473) );
  NOR2_X4 U4419 ( .A1(n3474), .A2(n3473), .ZN(n3426) );
  INV_X4 U4420 ( .A(n3429), .ZN(n3446) );
  INV_X4 U4421 ( .A(n3445), .ZN(n3432) );
  OAI22_X2 U4422 ( .A1(n3446), .A2(n3445), .B1(n3432), .B2(n3431), .ZN(n3437)
         );
  INV_X4 U4423 ( .A(n3433), .ZN(n3435) );
  NAND3_X2 U4424 ( .A1(n3435), .A2(n4043), .A3(n3434), .ZN(n3436) );
  NAND3_X2 U4425 ( .A1(n3436), .A2(n3437), .A3(n3438), .ZN(n3457) );
  INV_X4 U4426 ( .A(n3457), .ZN(n3555) );
  NAND2_X2 U4427 ( .A1(n3440), .A2(n3439), .ZN(n3449) );
  NAND2_X2 U4428 ( .A1(n3440), .A2(n3447), .ZN(n3858) );
  INV_X4 U4429 ( .A(n3552), .ZN(n3444) );
  NAND2_X2 U4430 ( .A1(n3446), .A2(n3445), .ZN(n4059) );
  NAND2_X2 U4431 ( .A1(n3448), .A2(n3447), .ZN(n3455) );
  INV_X4 U4432 ( .A(n3449), .ZN(n3856) );
  NAND4_X2 U4433 ( .A1(n3454), .A2(n1125), .A3(n3455), .A4(n1598), .ZN(n4057)
         );
  XNOR2_X2 U4434 ( .A(n3466), .B(n3465), .ZN(n3467) );
  NOR2_X4 U4435 ( .A1(n3468), .A2(n3467), .ZN(n3472) );
  NAND3_X4 U4436 ( .A1(n1512), .A2(n3472), .A3(n1244), .ZN(n3629) );
  NAND2_X2 U4437 ( .A1(a[16]), .A2(net297254), .ZN(n3699) );
  INV_X4 U4438 ( .A(n3699), .ZN(n3543) );
  INV_X4 U4440 ( .A(n3608), .ZN(n3506) );
  NAND2_X2 U4441 ( .A1(a[17]), .A2(net297204), .ZN(n3540) );
  NAND4_X2 U4442 ( .A1(n3508), .A2(n3510), .A3(n3509), .A4(n4288), .ZN(n3581)
         );
  NAND3_X2 U4443 ( .A1(n3581), .A2(n1604), .A3(n1273), .ZN(n3601) );
  NAND2_X2 U4444 ( .A1(a[19]), .A2(net297244), .ZN(n3530) );
  INV_X4 U4445 ( .A(n3530), .ZN(n3527) );
  INV_X4 U4446 ( .A(n3515), .ZN(n3516) );
  NAND2_X2 U4447 ( .A1(a[20]), .A2(net297226), .ZN(n3525) );
  INV_X4 U4448 ( .A(n3522), .ZN(n3589) );
  XNOR2_X2 U4449 ( .A(n3589), .B(n1170), .ZN(n3523) );
  INV_X4 U4450 ( .A(n3523), .ZN(n3524) );
  NAND2_X2 U4451 ( .A1(a[21]), .A2(net297260), .ZN(net295012) );
  NAND2_X2 U4452 ( .A1(n3525), .A2(net295010), .ZN(n3526) );
  XNOR2_X2 U4453 ( .A(n3597), .B(net294911), .ZN(n3528) );
  XNOR2_X2 U4454 ( .A(n3602), .B(net294901), .ZN(n3532) );
  NAND2_X2 U4455 ( .A1(n3606), .A2(n3683), .ZN(n3534) );
  NAND3_X4 U4458 ( .A1(net294993), .A2(n3537), .A3(n1683), .ZN(n3539) );
  XNOR2_X2 U4459 ( .A(n3606), .B(n3539), .ZN(n3573) );
  INV_X4 U4460 ( .A(n3547), .ZN(n3545) );
  NAND2_X2 U4461 ( .A1(\set_product_in_sig/z1 [23]), .A2(net297190), .ZN(n3546) );
  NAND2_X2 U4462 ( .A1(n3545), .A2(n3546), .ZN(n3549) );
  INV_X4 U4463 ( .A(n3546), .ZN(n3548) );
  OAI21_X4 U4464 ( .B1(n1562), .B2(net297188), .A(n4055), .ZN(n3556) );
  XNOR2_X2 U4465 ( .A(n3551), .B(n3550), .ZN(product_out[23]) );
  INV_X4 U4466 ( .A(n3863), .ZN(n3553) );
  NAND2_X2 U4467 ( .A1(n3556), .A2(n3862), .ZN(n3557) );
  OAI21_X4 U4468 ( .B1(n1689), .B2(n3557), .A(n3789), .ZN(n3558) );
  AOI21_X4 U4470 ( .B1(n3568), .B2(n3633), .A(n3567), .ZN(n3621) );
  NAND3_X4 U4471 ( .A1(n3569), .A2(n1705), .A3(n3571), .ZN(n3685) );
  NAND3_X2 U4472 ( .A1(n3578), .A2(n1514), .A3(n3577), .ZN(n3580) );
  NAND3_X2 U4473 ( .A1(n1604), .A2(n3581), .A3(n1273), .ZN(n3643) );
  OAI21_X4 U4474 ( .B1(n3584), .B2(n3583), .A(n1604), .ZN(n3644) );
  NAND2_X2 U4475 ( .A1(a[19]), .A2(net297216), .ZN(net294772) );
  NAND2_X2 U4476 ( .A1(a[22]), .A2(net297260), .ZN(n3593) );
  NAND2_X2 U4477 ( .A1(n3585), .A2(n3586), .ZN(n3588) );
  INV_X4 U4478 ( .A(n3586), .ZN(n3587) );
  NAND2_X2 U4479 ( .A1(n3588), .A2(n3646), .ZN(n3647) );
  NAND2_X2 U4480 ( .A1(n3589), .A2(n1170), .ZN(n3591) );
  NAND2_X2 U4481 ( .A1(n3593), .A2(n3592), .ZN(n3661) );
  INV_X4 U4483 ( .A(n1584), .ZN(n3598) );
  NOR2_X4 U4484 ( .A1(net294909), .A2(net294910), .ZN(net294907) );
  XNOR2_X2 U4485 ( .A(net294792), .B(net294905), .ZN(n3743) );
  NAND3_X2 U4487 ( .A1(n3609), .A2(n3608), .A3(net294888), .ZN(n3610) );
  NAND2_X2 U4488 ( .A1(a[18]), .A2(net297204), .ZN(net294881) );
  INV_X4 U4489 ( .A(net294882), .ZN(net294788) );
  INV_X4 U4490 ( .A(net294881), .ZN(net294879) );
  NAND2_X2 U4491 ( .A1(n3732), .A2(net294698), .ZN(n3687) );
  XNOR2_X2 U4492 ( .A(n3612), .B(n3910), .ZN(n3698) );
  NAND2_X2 U4493 ( .A1(a[17]), .A2(net297254), .ZN(n3697) );
  INV_X4 U4494 ( .A(n3697), .ZN(n3614) );
  NAND2_X2 U4496 ( .A1(net294053), .A2(n3615), .ZN(n3616) );
  NAND2_X2 U4497 ( .A1(\set_product_in_sig/z1 [24]), .A2(net297190), .ZN(n4062) );
  INV_X4 U4498 ( .A(n4062), .ZN(n3623) );
  XNOR2_X2 U4499 ( .A(n4063), .B(n3623), .ZN(n4054) );
  XNOR2_X2 U4500 ( .A(n3621), .B(n3620), .ZN(n3788) );
  INV_X4 U4501 ( .A(n3633), .ZN(n3634) );
  NAND2_X2 U4502 ( .A1(net294053), .A2(n3638), .ZN(n3641) );
  NAND2_X2 U4503 ( .A1(net294051), .A2(n3639), .ZN(n3640) );
  NAND2_X2 U4504 ( .A1(n3713), .A2(n3877), .ZN(n3695) );
  NAND2_X2 U4505 ( .A1(a[20]), .A2(net297216), .ZN(n3666) );
  INV_X4 U4506 ( .A(n3666), .ZN(n3665) );
  NAND3_X4 U4507 ( .A1(n3643), .A2(n3644), .A3(net294844), .ZN(net294843) );
  NAND2_X2 U4508 ( .A1(a[23]), .A2(net297260), .ZN(n3657) );
  INV_X4 U4511 ( .A(n3649), .ZN(n3747) );
  NAND2_X2 U4512 ( .A1(a[25]), .A2(net297485), .ZN(n3650) );
  INV_X4 U4513 ( .A(n3650), .ZN(n3746) );
  XNOR2_X2 U4514 ( .A(n3747), .B(n3746), .ZN(n3652) );
  NAND2_X2 U4515 ( .A1(n3651), .A2(n3652), .ZN(n3655) );
  INV_X4 U4516 ( .A(n3652), .ZN(n3654) );
  NAND2_X2 U4517 ( .A1(n3655), .A2(n3748), .ZN(n3656) );
  NAND2_X2 U4518 ( .A1(n3657), .A2(n3656), .ZN(n3660) );
  INV_X4 U4519 ( .A(n3656), .ZN(n3659) );
  INV_X4 U4520 ( .A(n3657), .ZN(n3658) );
  NAND2_X2 U4521 ( .A1(n3659), .A2(n3658), .ZN(n3759) );
  XNOR2_X2 U4522 ( .A(n3760), .B(n3758), .ZN(net294809) );
  NAND2_X2 U4523 ( .A1(a[22]), .A2(net297226), .ZN(net294810) );
  INV_X4 U4524 ( .A(net294810), .ZN(net294808) );
  NAND2_X2 U4525 ( .A1(net294808), .A2(net294809), .ZN(net294651) );
  XNOR2_X2 U4526 ( .A(net294800), .B(net294801), .ZN(n3667) );
  INV_X4 U4527 ( .A(net294772), .ZN(net294791) );
  INV_X4 U4529 ( .A(n3672), .ZN(n3676) );
  XNOR2_X2 U4530 ( .A(n3678), .B(n3679), .ZN(n3726) );
  INV_X4 U4531 ( .A(n3909), .ZN(n3912) );
  XNOR2_X2 U4532 ( .A(n3691), .B(n3690), .ZN(n3720) );
  NAND2_X2 U4533 ( .A1(n3713), .A2(n3693), .ZN(n3694) );
  OAI21_X4 U4535 ( .B1(n3708), .B2(n3707), .A(n3706), .ZN(n3721) );
  AOI21_X4 U4536 ( .B1(n3711), .B2(n1337), .A(n1263), .ZN(n3712) );
  INV_X4 U4537 ( .A(n3830), .ZN(n3831) );
  NAND3_X2 U4538 ( .A1(n3745), .A2(net294448), .A3(n3744), .ZN(n3766) );
  NAND2_X2 U4539 ( .A1(a[21]), .A2(net297216), .ZN(net294640) );
  NAND2_X2 U4540 ( .A1(a[23]), .A2(net297226), .ZN(n3763) );
  NAND2_X2 U4541 ( .A1(a[24]), .A2(net297260), .ZN(n3756) );
  NAND2_X2 U4542 ( .A1(n3747), .A2(n3746), .ZN(n3749) );
  NAND2_X2 U4543 ( .A1(n3751), .A2(n3752), .ZN(n3754) );
  INV_X4 U4544 ( .A(n3752), .ZN(n3753) );
  XNOR2_X2 U4545 ( .A(n3806), .B(n1281), .ZN(n3757) );
  INV_X4 U4546 ( .A(n3757), .ZN(n3755) );
  NAND2_X2 U4547 ( .A1(n3756), .A2(n3755), .ZN(n3814) );
  NAND3_X2 U4548 ( .A1(a[24]), .A2(n3757), .A3(net297260), .ZN(n3816) );
  INV_X4 U4549 ( .A(n3758), .ZN(n3761) );
  OAI21_X4 U4550 ( .B1(n3761), .B2(n3760), .A(n3759), .ZN(n3815) );
  NAND2_X2 U4552 ( .A1(n3763), .A2(n3762), .ZN(n3802) );
  NAND3_X2 U4553 ( .A1(n3764), .A2(net297226), .A3(a[23]), .ZN(n3937) );
  NAND2_X2 U4554 ( .A1(n3802), .A2(n3937), .ZN(n3765) );
  OAI21_X4 U4555 ( .B1(net294649), .B2(net294650), .A(net294651), .ZN(n3803)
         );
  XNOR2_X2 U4556 ( .A(n3803), .B(n3765), .ZN(net294645) );
  NAND2_X2 U4557 ( .A1(a[22]), .A2(net297244), .ZN(net294646) );
  XNOR2_X2 U4558 ( .A(net294642), .B(net294643), .ZN(net294580) );
  NAND2_X2 U4560 ( .A1(a[20]), .A2(net297204), .ZN(net294394) );
  INV_X4 U4561 ( .A(net294394), .ZN(net294388) );
  XNOR2_X2 U4562 ( .A(n3773), .B(n1256), .ZN(n3767) );
  NAND2_X2 U4563 ( .A1(a[19]), .A2(net297254), .ZN(n3772) );
  INV_X4 U4564 ( .A(n3772), .ZN(n3835) );
  XNOR2_X2 U4565 ( .A(net294628), .B(n1581), .ZN(n3774) );
  XNOR2_X2 U4567 ( .A(n3783), .B(n3782), .ZN(n3871) );
  XNOR2_X2 U4568 ( .A(n3784), .B(n1189), .ZN(product_out[26]) );
  INV_X4 U4569 ( .A(n4055), .ZN(n3854) );
  NAND3_X2 U4570 ( .A1(n3854), .A2(n3862), .A3(n3788), .ZN(n3793) );
  INV_X4 U4571 ( .A(n3789), .ZN(n3790) );
  INV_X4 U4572 ( .A(n4060), .ZN(n3865) );
  NOR3_X4 U4573 ( .A1(net293929), .A2(n3865), .A3(n1596), .ZN(n3792) );
  NOR2_X4 U4574 ( .A1(n3797), .A2(n3796), .ZN(n3852) );
  NAND2_X2 U4575 ( .A1(a[21]), .A2(net297204), .ZN(net294525) );
  INV_X4 U4576 ( .A(net294450), .ZN(net294578) );
  INV_X4 U4577 ( .A(n3804), .ZN(n3884) );
  XNOR2_X2 U4578 ( .A(n3884), .B(n1171), .ZN(n3809) );
  INV_X4 U4579 ( .A(n3809), .ZN(n3807) );
  NAND2_X2 U4580 ( .A1(a[25]), .A2(net297260), .ZN(n3811) );
  NOR2_X4 U4581 ( .A1(n1173), .A2(n3811), .ZN(n3812) );
  NAND2_X2 U4582 ( .A1(n3813), .A2(n3947), .ZN(n3887) );
  INV_X4 U4583 ( .A(n3814), .ZN(n3818) );
  INV_X4 U4584 ( .A(n3815), .ZN(n3817) );
  OAI21_X4 U4585 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(n3888) );
  XNOR2_X2 U4586 ( .A(n3887), .B(n3888), .ZN(n3821) );
  INV_X4 U4587 ( .A(n3821), .ZN(n3819) );
  NAND2_X2 U4588 ( .A1(a[24]), .A2(net297226), .ZN(n3820) );
  NAND2_X2 U4589 ( .A1(n3819), .A2(n3820), .ZN(n3823) );
  INV_X4 U4590 ( .A(n3820), .ZN(n3822) );
  XNOR2_X2 U4591 ( .A(n3878), .B(n3940), .ZN(net294543) );
  NAND2_X2 U4592 ( .A1(a[23]), .A2(net297244), .ZN(net294544) );
  NAND2_X2 U4593 ( .A1(a[20]), .A2(net297254), .ZN(net294366) );
  OAI22_X2 U4594 ( .A1(net294126), .A2(n3825), .B1(n3824), .B2(net294519), 
        .ZN(n3845) );
  INV_X4 U4595 ( .A(n3845), .ZN(n3827) );
  NAND2_X2 U4596 ( .A1(\set_product_in_sig/z1 [27]), .A2(net297190), .ZN(n3843) );
  XNOR2_X2 U4598 ( .A(n3832), .B(net294506), .ZN(n3837) );
  NAND2_X2 U4599 ( .A1(n3837), .A2(n3916), .ZN(n3840) );
  NAND3_X2 U4600 ( .A1(n3837), .A2(n3916), .A3(n1334), .ZN(n3838) );
  INV_X4 U4601 ( .A(n3842), .ZN(n3846) );
  INV_X4 U4602 ( .A(n3843), .ZN(n3844) );
  INV_X4 U4603 ( .A(n3848), .ZN(n3849) );
  INV_X4 U4604 ( .A(net299066), .ZN(net294479) );
  NOR2_X4 U4605 ( .A1(net293929), .A2(net294479), .ZN(n3872) );
  INV_X4 U4606 ( .A(n3858), .ZN(n3860) );
  NOR3_X4 U4607 ( .A1(n1596), .A2(n3866), .A3(n3865), .ZN(n3867) );
  NAND3_X2 U4608 ( .A1(n3715), .A2(n3870), .A3(n1623), .ZN(net294217) );
  NAND2_X2 U4610 ( .A1(a[23]), .A2(net297216), .ZN(net294253) );
  OAI21_X4 U4612 ( .B1(n3879), .B2(n3940), .A(n3939), .ZN(n3896) );
  NAND2_X2 U4613 ( .A1(a[25]), .A2(net297228), .ZN(n3893) );
  INV_X4 U4614 ( .A(n3893), .ZN(n3892) );
  NAND2_X2 U4615 ( .A1(a[27]), .A2(net297272), .ZN(n3880) );
  NAND2_X2 U4616 ( .A1(n3880), .A2(n3881), .ZN(n3883) );
  INV_X4 U4617 ( .A(n3881), .ZN(n3882) );
  NAND3_X4 U4618 ( .A1(a[27]), .A2(n3882), .A3(net297272), .ZN(n3951) );
  NAND2_X2 U4619 ( .A1(n3883), .A2(n3951), .ZN(n3952) );
  NAND2_X2 U4620 ( .A1(n3884), .A2(n1171), .ZN(n3886) );
  NAND3_X2 U4621 ( .A1(a[26]), .A2(net294426), .A3(net297260), .ZN(n3946) );
  INV_X4 U4622 ( .A(n3946), .ZN(n4013) );
  INV_X4 U4623 ( .A(a[26]), .ZN(net293991) );
  INV_X4 U4624 ( .A(net294426), .ZN(net294425) );
  NOR2_X4 U4625 ( .A1(n4013), .A2(net294285), .ZN(n3891) );
  INV_X4 U4626 ( .A(n3887), .ZN(n3889) );
  INV_X4 U4627 ( .A(n4014), .ZN(n3890) );
  NAND2_X2 U4628 ( .A1(n3892), .A2(n1579), .ZN(n3944) );
  INV_X4 U4629 ( .A(n1579), .ZN(n3894) );
  NAND2_X2 U4630 ( .A1(n3894), .A2(n3893), .ZN(n3942) );
  NAND2_X2 U4631 ( .A1(n3944), .A2(n3942), .ZN(n3895) );
  XNOR2_X2 U4632 ( .A(n3896), .B(n3895), .ZN(n3899) );
  INV_X4 U4633 ( .A(n1610), .ZN(n3897) );
  NAND2_X2 U4634 ( .A1(a[24]), .A2(net297244), .ZN(n3898) );
  NAND2_X2 U4635 ( .A1(n3897), .A2(n3898), .ZN(n3901) );
  INV_X4 U4636 ( .A(n3898), .ZN(n3900) );
  NAND2_X2 U4637 ( .A1(net294393), .A2(net294394), .ZN(n3903) );
  NOR2_X4 U4638 ( .A1(n3913), .A2(net294379), .ZN(n3914) );
  INV_X4 U4639 ( .A(net294366), .ZN(net294358) );
  AOI21_X4 U4640 ( .B1(n1400), .B2(net294322), .A(net294362), .ZN(net294360)
         );
  INV_X4 U4641 ( .A(net294356), .ZN(net294088) );
  XNOR2_X2 U4644 ( .A(n3921), .B(n3920), .ZN(n3926) );
  NAND2_X2 U4645 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  NAND3_X2 U4646 ( .A1(n3933), .A2(net298969), .A3(net294040), .ZN(n3988) );
  NAND2_X2 U4647 ( .A1(a[24]), .A2(net297216), .ZN(n3975) );
  INV_X4 U4648 ( .A(n3975), .ZN(n3974) );
  NAND3_X2 U4649 ( .A1(n3943), .A2(n3942), .A3(n3941), .ZN(n3945) );
  NAND2_X2 U4650 ( .A1(a[26]), .A2(net297226), .ZN(n3965) );
  NAND2_X2 U4651 ( .A1(a[28]), .A2(net297274), .ZN(n3949) );
  INV_X4 U4652 ( .A(n3949), .ZN(n4007) );
  XNOR2_X2 U4653 ( .A(n4007), .B(n1172), .ZN(n3956) );
  INV_X4 U4654 ( .A(n3956), .ZN(n3954) );
  OAI21_X4 U4655 ( .B1(n3953), .B2(n3952), .A(n3951), .ZN(n3955) );
  NAND2_X2 U4656 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  NAND2_X2 U4657 ( .A1(n4008), .A2(n3958), .ZN(n3961) );
  INV_X4 U4658 ( .A(n3961), .ZN(n3960) );
  NAND2_X2 U4659 ( .A1(a[27]), .A2(net297260), .ZN(n3962) );
  INV_X4 U4660 ( .A(n3962), .ZN(n3959) );
  NAND2_X2 U4661 ( .A1(n3960), .A2(n3959), .ZN(n4015) );
  NAND2_X2 U4662 ( .A1(n3962), .A2(n3961), .ZN(n4012) );
  NAND2_X2 U4663 ( .A1(n4015), .A2(n4012), .ZN(n3963) );
  XNOR2_X2 U4664 ( .A(n3964), .B(n3963), .ZN(n3966) );
  NAND2_X2 U4665 ( .A1(n3965), .A2(n1580), .ZN(n3967) );
  NAND3_X2 U4666 ( .A1(n3966), .A2(a[26]), .A3(net297226), .ZN(n3999) );
  XNOR2_X2 U4667 ( .A(n3998), .B(n4000), .ZN(n3968) );
  NAND3_X2 U4668 ( .A1(a[25]), .A2(n3968), .A3(net297244), .ZN(n4027) );
  NAND2_X2 U4669 ( .A1(a[25]), .A2(net297244), .ZN(n3970) );
  INV_X4 U4670 ( .A(n3968), .ZN(n3969) );
  XNOR2_X2 U4671 ( .A(n3972), .B(n3971), .ZN(n3976) );
  INV_X4 U4672 ( .A(n3976), .ZN(n3973) );
  NAND2_X2 U4674 ( .A1(n1114), .A2(n3975), .ZN(n3980) );
  INV_X4 U4675 ( .A(n3980), .ZN(n3977) );
  INV_X4 U4676 ( .A(net294250), .ZN(net294194) );
  OAI21_X4 U4677 ( .B1(n4038), .B2(n3977), .A(net294194), .ZN(n3979) );
  NAND2_X2 U4678 ( .A1(net294251), .A2(net294252), .ZN(n3981) );
  XNOR2_X2 U4679 ( .A(n3978), .B(n3979), .ZN(n3985) );
  XNOR2_X2 U4680 ( .A(n3983), .B(n3982), .ZN(n3984) );
  XNOR2_X2 U4681 ( .A(n3986), .B(n4098), .ZN(net294234) );
  INV_X4 U4682 ( .A(n4098), .ZN(n3990) );
  XNOR2_X2 U4683 ( .A(n3989), .B(n3990), .ZN(n3991) );
  NAND2_X2 U4684 ( .A1(n1285), .A2(n3995), .ZN(net294101) );
  NAND2_X2 U4685 ( .A1(n1501), .A2(net294101), .ZN(net294117) );
  OAI21_X4 U4686 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4041) );
  NAND2_X2 U4687 ( .A1(a[23]), .A2(net297254), .ZN(n4091) );
  INV_X4 U4688 ( .A(n4091), .ZN(n4079) );
  XNOR2_X2 U4689 ( .A(n1261), .B(n4079), .ZN(n4039) );
  NAND2_X2 U4690 ( .A1(a[25]), .A2(net297216), .ZN(n4101) );
  INV_X4 U4691 ( .A(n3998), .ZN(n4001) );
  INV_X4 U4693 ( .A(n4022), .ZN(n4020) );
  INV_X4 U4694 ( .A(n4004), .ZN(n4003) );
  NAND2_X2 U4695 ( .A1(n4003), .A2(n4002), .ZN(n4121) );
  NAND2_X2 U4696 ( .A1(n4007), .A2(n1172), .ZN(n4009) );
  NAND2_X2 U4697 ( .A1(a[28]), .A2(net297260), .ZN(n4116) );
  XNOR2_X2 U4698 ( .A(n4115), .B(n4116), .ZN(n4011) );
  NAND2_X2 U4699 ( .A1(a[27]), .A2(net297228), .ZN(n4111) );
  XNOR2_X2 U4700 ( .A(n4141), .B(n4111), .ZN(n4019) );
  INV_X4 U4701 ( .A(n4012), .ZN(n4017) );
  INV_X4 U4702 ( .A(n4018), .ZN(n4140) );
  XNOR2_X2 U4703 ( .A(n4019), .B(n4140), .ZN(n4021) );
  INV_X4 U4704 ( .A(n4021), .ZN(n4023) );
  NAND2_X2 U4705 ( .A1(n4023), .A2(n4022), .ZN(n4110) );
  NAND2_X2 U4706 ( .A1(n4024), .A2(n4110), .ZN(n4108) );
  NAND2_X2 U4707 ( .A1(a[26]), .A2(net297244), .ZN(n4109) );
  INV_X4 U4708 ( .A(n4109), .ZN(n4025) );
  XNOR2_X2 U4711 ( .A(n4030), .B(n4107), .ZN(n4036) );
  XNOR2_X2 U4712 ( .A(n4039), .B(n4076), .ZN(n4040) );
  INV_X4 U4713 ( .A(n4043), .ZN(n4047) );
  XNOR2_X2 U4714 ( .A(n4047), .B(n4046), .ZN(n4053) );
  OAI21_X4 U4715 ( .B1(n4053), .B2(net297279), .A(n4052), .ZN(n4173) );
  INV_X4 U4716 ( .A(net293935), .ZN(net294092) );
  AOI21_X4 U4717 ( .B1(n4065), .B2(n4066), .A(n4064), .ZN(n4177) );
  NAND2_X2 U4718 ( .A1(n1548), .A2(net294101), .ZN(n4068) );
  INV_X4 U4719 ( .A(n4068), .ZN(n4175) );
  NAND2_X2 U4720 ( .A1(n4073), .A2(n4074), .ZN(product_out[30]) );
  NOR2_X4 U4721 ( .A1(n1613), .A2(n4091), .ZN(n4083) );
  OAI21_X4 U4724 ( .B1(n1369), .B2(n4094), .A(n4093), .ZN(n4170) );
  NAND2_X2 U4725 ( .A1(net294051), .A2(net294052), .ZN(n4095) );
  INV_X4 U4726 ( .A(n4165), .ZN(n4163) );
  NAND2_X2 U4727 ( .A1(\set_product_in_sig/z1 [31]), .A2(net297190), .ZN(n4164) );
  NAND2_X2 U4728 ( .A1(n4163), .A2(n4164), .ZN(n4097) );
  INV_X4 U4729 ( .A(n4097), .ZN(n4161) );
  OAI21_X4 U4730 ( .B1(n4099), .B2(n4100), .A(n4281), .ZN(n4156) );
  INV_X4 U4731 ( .A(n4101), .ZN(n4103) );
  NAND2_X2 U4732 ( .A1(n4103), .A2(n4102), .ZN(n4105) );
  NAND2_X2 U4733 ( .A1(n4104), .A2(n4105), .ZN(n4151) );
  XNOR2_X2 U4735 ( .A(n4141), .B(n4140), .ZN(n4112) );
  NOR2_X2 U4736 ( .A1(n4112), .A2(n4111), .ZN(n4113) );
  NOR2_X4 U4737 ( .A1(n4114), .A2(n4113), .ZN(n4145) );
  NOR2_X4 U4738 ( .A1(n1541), .A2(n4116), .ZN(n4139) );
  INV_X4 U4739 ( .A(a[31]), .ZN(n4117) );
  NOR2_X4 U4740 ( .A1(net294016), .A2(n4117), .ZN(n4120) );
  INV_X4 U4741 ( .A(a[30]), .ZN(n4118) );
  INV_X4 U4742 ( .A(a[24]), .ZN(net294012) );
  FA_X1 U4743 ( .A(n4120), .B(n4119), .CI(net294010), .S(n4124) );
  INV_X4 U4744 ( .A(n4121), .ZN(n4122) );
  INV_X4 U4745 ( .A(a[29]), .ZN(net294006) );
  XNOR2_X2 U4746 ( .A(n4122), .B(net294004), .ZN(n4123) );
  XNOR2_X2 U4747 ( .A(n4124), .B(n4123), .ZN(n4133) );
  INV_X4 U4748 ( .A(a[27]), .ZN(n4125) );
  NOR2_X4 U4749 ( .A1(net297250), .A2(n4125), .ZN(n4128) );
  INV_X4 U4750 ( .A(a[28]), .ZN(n4126) );
  NOR2_X4 U4751 ( .A1(net297234), .A2(n4126), .ZN(n4127) );
  XNOR2_X2 U4752 ( .A(n4128), .B(n4127), .ZN(n4131) );
  NOR2_X4 U4753 ( .A1(net297222), .A2(net293991), .ZN(n4129) );
  INV_X4 U4754 ( .A(a[25]), .ZN(net293988) );
  XNOR2_X2 U4755 ( .A(n4129), .B(net293986), .ZN(n4130) );
  XNOR2_X2 U4756 ( .A(n4131), .B(n4130), .ZN(n4132) );
  XNOR2_X2 U4757 ( .A(n4133), .B(n4132), .ZN(n4137) );
  NOR2_X4 U4758 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  XNOR2_X2 U4759 ( .A(n4137), .B(n4136), .ZN(n4138) );
  XNOR2_X2 U4760 ( .A(n4139), .B(n4138), .ZN(n4143) );
  XNOR2_X2 U4761 ( .A(n4143), .B(n4142), .ZN(n4144) );
  XNOR2_X2 U4762 ( .A(n4145), .B(n4144), .ZN(n4146) );
  XNOR2_X2 U4763 ( .A(n4147), .B(n4146), .ZN(n4148) );
  XNOR2_X2 U4764 ( .A(n4149), .B(n4148), .ZN(n4150) );
  XNOR2_X2 U4765 ( .A(n4151), .B(n4150), .ZN(n4154) );
  INV_X4 U4766 ( .A(n4076), .ZN(n4152) );
  NAND2_X2 U4767 ( .A1(n4152), .A2(n1261), .ZN(n4153) );
  XNOR2_X2 U4768 ( .A(n4154), .B(n4153), .ZN(n4155) );
  XNOR2_X2 U4769 ( .A(n4156), .B(n4155), .ZN(n4159) );
  NOR2_X4 U4770 ( .A1(n4158), .A2(n4157), .ZN(n4172) );
  INV_X4 U4771 ( .A(n4159), .ZN(n4160) );
  NAND2_X2 U4772 ( .A1(n4164), .A2(net297190), .ZN(n4162) );
  NAND2_X2 U4773 ( .A1(n4163), .A2(n4162), .ZN(n4167) );
  NAND2_X2 U4774 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  NAND2_X2 U4775 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  OAI21_X4 U4776 ( .B1(n4170), .B2(n4169), .A(n4168), .ZN(n4171) );
  NOR2_X4 U4777 ( .A1(n4172), .A2(n4171), .ZN(n4185) );
  NAND2_X2 U4778 ( .A1(n1288), .A2(n4173), .ZN(n4174) );
  NAND3_X2 U4779 ( .A1(net293933), .A2(n4175), .A3(n4179), .ZN(n4183) );
  OAI211_X2 U4780 ( .C1(n4177), .C2(n4176), .A(net293927), .B(n1548), .ZN(
        n4182) );
  NAND2_X2 U4781 ( .A1(net294093), .A2(n4178), .ZN(n4180) );
  NAND2_X2 U4782 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  NAND2_X2 U1133 ( .A1(n2776), .A2(net295756), .ZN(n2782) );
  INV_X2 U1140 ( .A(n2782), .ZN(n2779) );
  NAND2_X2 U1142 ( .A1(n1392), .A2(net294330), .ZN(n1391) );
  BUF_X32 U1143 ( .A(n1852), .Z(n4196) );
  INV_X2 U1154 ( .A(n4026), .ZN(n4029) );
  XNOR2_X2 U1155 ( .A(n3339), .B(n3340), .ZN(n4197) );
  OAI21_X4 U1156 ( .B1(n3337), .B2(n3338), .A(n1119), .ZN(n3339) );
  CLKBUF_X3 U1159 ( .A(net294842), .Z(net297593) );
  XNOR2_X2 U1162 ( .A(n2602), .B(n2764), .ZN(n1528) );
  INV_X1 U1166 ( .A(net294793), .ZN(net298389) );
  INV_X8 U1170 ( .A(n2225), .ZN(n2199) );
  OAI21_X2 U1175 ( .B1(n2848), .B2(n2676), .A(n2675), .ZN(n4198) );
  NOR2_X4 U1176 ( .A1(n2674), .A2(n2673), .ZN(n2675) );
  NAND2_X2 U1183 ( .A1(n2011), .A2(n2010), .ZN(n2054) );
  NAND2_X2 U1190 ( .A1(n3301), .A2(n3302), .ZN(n4199) );
  CLKBUF_X3 U1219 ( .A(n3135), .Z(n4200) );
  XNOR2_X2 U1220 ( .A(net296530), .B(n4282), .ZN(n4201) );
  INV_X4 U1226 ( .A(net296425), .ZN(n4282) );
  INV_X8 U1228 ( .A(n2935), .ZN(n3045) );
  XNOR2_X2 U1232 ( .A(n2682), .B(n2773), .ZN(n4202) );
  INV_X2 U1235 ( .A(n1144), .ZN(n4203) );
  INV_X2 U1239 ( .A(n1976), .ZN(n1144) );
  NAND2_X2 U1240 ( .A1(n2028), .A2(n2027), .ZN(n2048) );
  AOI21_X2 U1241 ( .B1(n1127), .B2(n3382), .A(n1115), .ZN(n3234) );
  INV_X4 U1248 ( .A(net294645), .ZN(n1462) );
  INV_X2 U1255 ( .A(n3280), .ZN(n3095) );
  OAI211_X2 U1256 ( .C1(n3096), .C2(n3095), .A(n3278), .B(n3094), .ZN(n3097)
         );
  OAI21_X4 U1258 ( .B1(n3575), .B2(n3576), .A(n4261), .ZN(n4290) );
  CLKBUF_X2 U1259 ( .A(n2295), .Z(n4204) );
  NAND2_X2 U1267 ( .A1(n3301), .A2(n3302), .ZN(n3570) );
  INV_X4 U1270 ( .A(n4199), .ZN(n3303) );
  INV_X16 U1272 ( .A(net296416), .ZN(net298909) );
  OAI21_X2 U1278 ( .B1(n2696), .B2(n2695), .A(n2694), .ZN(n2867) );
  NAND3_X1 U1287 ( .A1(n3938), .A2(n3939), .A3(n3937), .ZN(n3943) );
  NAND2_X2 U1288 ( .A1(n3905), .A2(n3835), .ZN(n3779) );
  XNOR2_X2 U1290 ( .A(n3339), .B(n3340), .ZN(n4205) );
  INV_X4 U1292 ( .A(n3606), .ZN(n3609) );
  NAND2_X2 U1295 ( .A1(n1528), .A2(n2603), .ZN(n2611) );
  OAI21_X1 U1297 ( .B1(n2203), .B2(n2586), .A(net296430), .ZN(n2589) );
  NAND2_X2 U1310 ( .A1(n1802), .A2(n2500), .ZN(n2501) );
  INV_X4 U1324 ( .A(net294658), .ZN(net294652) );
  XOR2_X2 U1325 ( .A(net294806), .B(net294655), .Z(n4206) );
  NAND2_X4 U1326 ( .A1(net294837), .A2(net294658), .ZN(net294806) );
  NAND2_X2 U1333 ( .A1(n1488), .A2(net294651), .ZN(net294655) );
  INV_X1 U1363 ( .A(n4106), .ZN(n4207) );
  AOI21_X4 U1364 ( .B1(n3705), .B2(n3704), .A(n3625), .ZN(n1363) );
  NAND2_X4 U1368 ( .A1(n3705), .A2(n3704), .ZN(n3706) );
  OAI211_X4 U1376 ( .C1(n3738), .C2(n1197), .A(n3737), .B(n3736), .ZN(n3739)
         );
  NAND4_X2 U1378 ( .A1(n2478), .A2(n2103), .A3(n2105), .A4(n1109), .ZN(n4208)
         );
  NAND2_X2 U1382 ( .A1(n2249), .A2(n2312), .ZN(n4211) );
  NAND2_X4 U1383 ( .A1(n4209), .A2(n4210), .ZN(n4212) );
  NAND2_X4 U1393 ( .A1(n4211), .A2(n4212), .ZN(n2251) );
  INV_X4 U1395 ( .A(n2249), .ZN(n4209) );
  INV_X2 U1396 ( .A(n2312), .ZN(n4210) );
  CLKBUF_X3 U1397 ( .A(n1928), .Z(n4213) );
  NAND4_X2 U1418 ( .A1(n2478), .A2(n2103), .A3(n2105), .A4(n1109), .ZN(n2246)
         );
  INV_X8 U1420 ( .A(n3909), .ZN(n4214) );
  INV_X16 U1426 ( .A(n4214), .ZN(n4215) );
  NAND2_X2 U1491 ( .A1(n3687), .A2(net294696), .ZN(n3909) );
  INV_X1 U1494 ( .A(n2571), .ZN(n1577) );
  NAND2_X1 U1501 ( .A1(n1385), .A2(net294228), .ZN(n4218) );
  NAND2_X2 U1504 ( .A1(n4216), .A2(n4217), .ZN(n4219) );
  NAND2_X2 U1527 ( .A1(n4218), .A2(n4219), .ZN(net294218) );
  INV_X4 U1534 ( .A(n1385), .ZN(n4216) );
  INV_X4 U1535 ( .A(net294228), .ZN(n4217) );
  OAI21_X4 U1548 ( .B1(net294218), .B2(net297188), .A(net294219), .ZN(
        net294200) );
  NAND2_X2 U1551 ( .A1(a[14]), .A2(net297485), .ZN(net296099) );
  NAND2_X1 U1561 ( .A1(n2082), .A2(n2149), .ZN(n4222) );
  NAND2_X4 U1573 ( .A1(n4220), .A2(n4221), .ZN(n4223) );
  NAND2_X2 U1581 ( .A1(n4222), .A2(n4223), .ZN(n2083) );
  INV_X4 U1610 ( .A(n2082), .ZN(n4220) );
  INV_X1 U1615 ( .A(n2149), .ZN(n4221) );
  BUF_X4 U1626 ( .A(net294300), .Z(net299137) );
  NAND2_X1 U1631 ( .A1(n1391), .A2(net294366), .ZN(n4226) );
  NAND2_X2 U1651 ( .A1(n4224), .A2(n4225), .ZN(n4227) );
  NAND2_X2 U1660 ( .A1(n4226), .A2(n4227), .ZN(n1390) );
  INV_X4 U1661 ( .A(n1391), .ZN(n4224) );
  INV_X4 U1667 ( .A(net294366), .ZN(n4225) );
  NAND2_X2 U1680 ( .A1(n1390), .A2(net294520), .ZN(n4230) );
  NAND2_X4 U1693 ( .A1(n4228), .A2(n4229), .ZN(n4231) );
  NAND2_X4 U1707 ( .A1(n4230), .A2(n4231), .ZN(n1389) );
  INV_X4 U1711 ( .A(n1390), .ZN(n4228) );
  INV_X4 U1752 ( .A(net294520), .ZN(n4229) );
  INV_X8 U1754 ( .A(n1389), .ZN(n1387) );
  AOI21_X2 U1804 ( .B1(n3396), .B2(n3514), .A(n4277), .ZN(n3397) );
  INV_X4 U1816 ( .A(n3799), .ZN(n3829) );
  INV_X4 U1819 ( .A(net294696), .ZN(net294883) );
  INV_X4 U1836 ( .A(n2472), .ZN(n2475) );
  NAND2_X2 U1840 ( .A1(n3780), .A2(n1571), .ZN(n4234) );
  NAND2_X4 U1850 ( .A1(n4232), .A2(n4233), .ZN(n4235) );
  NAND2_X4 U1879 ( .A1(n4234), .A2(n4235), .ZN(n1570) );
  INV_X4 U1900 ( .A(n3780), .ZN(n4232) );
  INV_X4 U1907 ( .A(n1571), .ZN(n4233) );
  CLKBUF_X2 U1913 ( .A(n1570), .Z(n1656) );
  INV_X4 U1914 ( .A(n3517), .ZN(n3402) );
  NAND2_X2 U1924 ( .A1(n1338), .A2(n4237), .ZN(n4236) );
  INV_X4 U1948 ( .A(n4236), .ZN(n2708) );
  INV_X32 U1949 ( .A(n2707), .ZN(n4237) );
  INV_X2 U1977 ( .A(n1338), .ZN(n2833) );
  INV_X1 U1981 ( .A(n1192), .ZN(n1150) );
  INV_X8 U1983 ( .A(n3102), .ZN(n3371) );
  NAND2_X4 U1988 ( .A1(n2521), .A2(n2555), .ZN(n2522) );
  INV_X2 U1990 ( .A(net294636), .ZN(net298392) );
  CLKBUF_X3 U1991 ( .A(n3099), .Z(n1111) );
  NAND2_X1 U2020 ( .A1(n3418), .A2(n3419), .ZN(n3681) );
  NAND2_X4 U2036 ( .A1(n1137), .A2(n1138), .ZN(n1633) );
  NAND2_X4 U2055 ( .A1(n1135), .A2(n1136), .ZN(n1138) );
  NAND2_X4 U2064 ( .A1(n4268), .A2(n1593), .ZN(n3499) );
  INV_X2 U2072 ( .A(n3263), .ZN(n1135) );
  INV_X2 U2075 ( .A(n3032), .ZN(n1175) );
  INV_X4 U2078 ( .A(n3874), .ZN(n3875) );
  INV_X4 U2089 ( .A(n3597), .ZN(n3599) );
  NAND2_X4 U2094 ( .A1(n2012), .A2(n1954), .ZN(n1182) );
  CLKBUF_X3 U2095 ( .A(net294198), .Z(n4238) );
  INV_X8 U2100 ( .A(net297615), .ZN(net297616) );
  INV_X4 U2123 ( .A(n3507), .ZN(n4287) );
  INV_X8 U2140 ( .A(n3776), .ZN(n3777) );
  CLKBUF_X3 U2151 ( .A(net294086), .Z(n4239) );
  XNOR2_X2 U2152 ( .A(net294354), .B(net299300), .ZN(n3917) );
  INV_X2 U2153 ( .A(net294639), .ZN(n1396) );
  NAND2_X1 U2170 ( .A1(n3831), .A2(n4215), .ZN(net294507) );
  INV_X2 U2178 ( .A(n3039), .ZN(n3040) );
  XNOR2_X1 U2191 ( .A(net294044), .B(net294334), .ZN(net294354) );
  INV_X2 U2193 ( .A(n4037), .ZN(n4032) );
  INV_X4 U2240 ( .A(n3513), .ZN(n3584) );
  INV_X4 U2303 ( .A(n3411), .ZN(n3409) );
  NAND2_X1 U2344 ( .A1(n4041), .A2(n1349), .ZN(n4242) );
  NAND2_X4 U2359 ( .A1(n4240), .A2(n4241), .ZN(n4243) );
  NAND2_X4 U2379 ( .A1(n4242), .A2(n4243), .ZN(n4092) );
  INV_X2 U2382 ( .A(n4089), .ZN(n4240) );
  INV_X2 U2387 ( .A(n1349), .ZN(n4241) );
  OAI21_X4 U2388 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4093) );
  OAI21_X4 U2433 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4089) );
  NAND3_X2 U2468 ( .A1(net294320), .A2(net294322), .A3(n4266), .ZN(n3931) );
  NAND2_X4 U2478 ( .A1(n1362), .A2(n3239), .ZN(n3240) );
  NAND2_X4 U2479 ( .A1(net295618), .A2(n3061), .ZN(n4272) );
  NAND2_X4 U2491 ( .A1(n1932), .A2(n1982), .ZN(n4244) );
  NAND2_X2 U2493 ( .A1(n4245), .A2(n1984), .ZN(n1937) );
  INV_X4 U2494 ( .A(n4244), .ZN(n4245) );
  NAND2_X4 U2495 ( .A1(n1917), .A2(n1916), .ZN(n1982) );
  INV_X4 U2506 ( .A(n1937), .ZN(n1938) );
  INV_X2 U2508 ( .A(n2643), .ZN(n4246) );
  INV_X2 U2513 ( .A(n4246), .ZN(n4247) );
  INV_X8 U2519 ( .A(n3003), .ZN(n3006) );
  NOR2_X2 U2537 ( .A1(n3200), .A2(n3199), .ZN(n3211) );
  BUF_X32 U2635 ( .A(n3221), .Z(n4248) );
  INV_X1 U2636 ( .A(n2819), .ZN(n1147) );
  NAND2_X4 U2649 ( .A1(n2150), .A2(n2151), .ZN(n4249) );
  BUF_X32 U2670 ( .A(n2644), .Z(n4250) );
  NAND2_X1 U2673 ( .A1(n2264), .A2(n2367), .ZN(n2169) );
  NAND2_X4 U2682 ( .A1(n3097), .A2(n3098), .ZN(n3177) );
  BUF_X16 U2690 ( .A(n2646), .Z(n1539) );
  INV_X2 U2708 ( .A(n1618), .ZN(n3297) );
  NAND2_X2 U2727 ( .A1(n2167), .A2(n2166), .ZN(n2367) );
  INV_X8 U2728 ( .A(n2630), .ZN(n1758) );
  NAND2_X4 U2734 ( .A1(n2536), .A2(n2535), .ZN(n2538) );
  INV_X8 U2739 ( .A(n3558), .ZN(n3717) );
  NOR2_X4 U2751 ( .A1(n3115), .A2(n3313), .ZN(n3131) );
  INV_X4 U2755 ( .A(n1499), .ZN(n3079) );
  NAND2_X2 U2762 ( .A1(n3469), .A2(n3470), .ZN(n4044) );
  INV_X8 U2763 ( .A(n3347), .ZN(n3469) );
  NAND2_X4 U2771 ( .A1(n3614), .A2(n3613), .ZN(n3692) );
  INV_X4 U2779 ( .A(n3685), .ZN(n3572) );
  INV_X4 U2805 ( .A(n3902), .ZN(n1533) );
  NAND4_X4 U2813 ( .A1(a[15]), .A2(n4276), .A3(net295732), .A4(net297260), 
        .ZN(n3144) );
  INV_X1 U2814 ( .A(n1657), .ZN(n4106) );
  NAND2_X2 U2819 ( .A1(n3908), .A2(n3907), .ZN(n4251) );
  NAND2_X4 U2847 ( .A1(n2302), .A2(n1632), .ZN(n2479) );
  INV_X4 U2857 ( .A(n2729), .ZN(n4252) );
  INV_X4 U2894 ( .A(n4252), .ZN(n4253) );
  NAND2_X2 U2909 ( .A1(n2095), .A2(n2094), .ZN(n2477) );
  NAND2_X4 U2915 ( .A1(n1280), .A2(n3083), .ZN(n1117) );
  NOR2_X4 U2917 ( .A1(n3083), .A2(n1280), .ZN(n1504) );
  NAND2_X1 U2929 ( .A1(n1690), .A2(n2908), .ZN(n2740) );
  INV_X8 U2934 ( .A(n2908), .ZN(n2624) );
  INV_X2 U2952 ( .A(n3091), .ZN(n4254) );
  NAND2_X2 U2954 ( .A1(n2620), .A2(n2621), .ZN(n2665) );
  INV_X2 U2975 ( .A(n4249), .ZN(n4255) );
  INV_X4 U2981 ( .A(n4255), .ZN(n4256) );
  NAND2_X4 U2985 ( .A1(n2276), .A2(n2173), .ZN(n2163) );
  NAND2_X2 U2987 ( .A1(n1353), .A2(n3552), .ZN(n3443) );
  INV_X8 U2993 ( .A(n2395), .ZN(n2255) );
  OAI21_X2 U3001 ( .B1(n1689), .B2(n3557), .A(n3789), .ZN(n4286) );
  NAND2_X1 U3068 ( .A1(n1280), .A2(n3083), .ZN(n1616) );
  NAND2_X4 U3075 ( .A1(n2526), .A2(n2654), .ZN(n2738) );
  NAND2_X4 U3120 ( .A1(n1305), .A2(n2655), .ZN(n2627) );
  NAND2_X2 U3172 ( .A1(n2256), .A2(n1309), .ZN(n2353) );
  INV_X2 U3184 ( .A(n2472), .ZN(n1778) );
  INV_X8 U3223 ( .A(n3554), .ZN(n1689) );
  OAI211_X2 U3228 ( .C1(n1803), .C2(n2319), .A(n2318), .B(n1625), .ZN(n2333)
         );
  NAND2_X2 U3236 ( .A1(n3223), .A2(n3224), .ZN(n3306) );
  NAND2_X4 U3248 ( .A1(n1943), .A2(n1942), .ZN(n1944) );
  INV_X8 U3250 ( .A(n2560), .ZN(n2653) );
  AND2_X2 U3256 ( .A1(n2255), .A2(n2398), .ZN(n4257) );
  NAND2_X4 U3270 ( .A1(a[4]), .A2(net297216), .ZN(n2398) );
  INV_X2 U3271 ( .A(n3283), .ZN(n3089) );
  BUF_X4 U3282 ( .A(n1590), .Z(n1314) );
  NAND2_X4 U3334 ( .A1(n1190), .A2(n2245), .ZN(n1590) );
  NAND2_X2 U3347 ( .A1(n2045), .A2(n2044), .ZN(n4258) );
  NAND2_X2 U3352 ( .A1(n2045), .A2(n2044), .ZN(n2176) );
  NAND2_X2 U3371 ( .A1(n3453), .A2(n3856), .ZN(n3454) );
  XOR2_X2 U3397 ( .A(n2078), .B(n2077), .Z(n1626) );
  NOR2_X4 U3400 ( .A1(n2094), .A2(n2076), .ZN(n2077) );
  INV_X2 U3436 ( .A(n2520), .ZN(n4259) );
  INV_X4 U3445 ( .A(n2520), .ZN(n1651) );
  NOR2_X4 U3446 ( .A1(n3083), .A2(n1280), .ZN(n4260) );
  BUF_X4 U3463 ( .A(n2234), .Z(n1505) );
  CLKBUF_X3 U3483 ( .A(n3574), .Z(n4261) );
  NAND3_X2 U3499 ( .A1(n2286), .A2(n1493), .A3(n2284), .ZN(n4262) );
  OAI21_X4 U3520 ( .B1(n3260), .B2(n3164), .A(n1198), .ZN(n1242) );
  CLKBUF_X3 U3525 ( .A(net294088), .Z(net298149) );
  INV_X2 U3571 ( .A(n3728), .ZN(n3731) );
  CLKBUF_X2 U3586 ( .A(n2412), .Z(n4263) );
  OAI21_X1 U3587 ( .B1(net295018), .B2(net295019), .A(net295020), .ZN(n4264)
         );
  INV_X4 U3589 ( .A(n3225), .ZN(n3226) );
  INV_X2 U3604 ( .A(n3225), .ZN(n1324) );
  NAND2_X4 U3657 ( .A1(n4084), .A2(net294068), .ZN(n4094) );
  INV_X16 U3668 ( .A(n3082), .ZN(n3083) );
  INV_X4 U3670 ( .A(net294611), .ZN(net295585) );
  INV_X4 U3679 ( .A(n4270), .ZN(n4265) );
  INV_X4 U3706 ( .A(n1597), .ZN(n4270) );
  INV_X8 U3718 ( .A(n3124), .ZN(n3072) );
  NAND2_X2 U3753 ( .A1(n2884), .A2(n2917), .ZN(n2744) );
  INV_X2 U3783 ( .A(net294510), .ZN(n4266) );
  INV_X1 U3807 ( .A(n1226), .ZN(n1151) );
  INV_X1 U3808 ( .A(n3906), .ZN(n4267) );
  INV_X4 U3858 ( .A(n3607), .ZN(n3673) );
  NAND2_X4 U3927 ( .A1(n3565), .A2(n1276), .ZN(n4268) );
  AND2_X4 U3930 ( .A1(n3487), .A2(n3486), .ZN(n1276) );
  INV_X8 U3964 ( .A(n3036), .ZN(n4269) );
  INV_X8 U3974 ( .A(n3161), .ZN(n3036) );
  INV_X1 U4002 ( .A(net294285), .ZN(n4271) );
  AOI21_X4 U4046 ( .B1(n3089), .B2(n3278), .A(n3088), .ZN(n3098) );
  NAND2_X4 U4052 ( .A1(n2661), .A2(n2625), .ZN(n2362) );
  INV_X1 U4120 ( .A(n3625), .ZN(n3701) );
  NAND2_X2 U4147 ( .A1(n3168), .A2(n3169), .ZN(n1559) );
  NAND2_X4 U4232 ( .A1(n4178), .A2(net293931), .ZN(n4179) );
  NAND2_X4 U4240 ( .A1(n4174), .A2(net293935), .ZN(net293931) );
  NAND3_X1 U4278 ( .A1(n4057), .A2(n4059), .A3(n4058), .ZN(n3551) );
  INV_X8 U4296 ( .A(n4260), .ZN(n3278) );
  AND2_X4 U4299 ( .A1(n1353), .A2(n3553), .ZN(n1306) );
  INV_X4 U4315 ( .A(net294447), .ZN(n1256) );
  NAND2_X2 U4343 ( .A1(net294447), .A2(net294448), .ZN(net294442) );
  XNOR2_X1 U4358 ( .A(net294447), .B(net294394), .ZN(net294628) );
  INV_X2 U4365 ( .A(net295995), .ZN(net296417) );
  NAND2_X2 U4366 ( .A1(n2317), .A2(n2316), .ZN(n4273) );
  NAND2_X4 U4367 ( .A1(n3301), .A2(n3302), .ZN(n1361) );
  INV_X4 U4368 ( .A(n3878), .ZN(n3879) );
  NAND2_X4 U4376 ( .A1(n3329), .A2(n3330), .ZN(n3392) );
  NAND2_X2 U4390 ( .A1(net294083), .A2(net294068), .ZN(net294228) );
  NAND2_X4 U4399 ( .A1(n3973), .A2(n3974), .ZN(n4274) );
  NAND2_X4 U4400 ( .A1(n2204), .A2(n1930), .ZN(n2323) );
  AOI21_X2 U4439 ( .B1(n3627), .B2(n3626), .A(n3701), .ZN(n3636) );
  INV_X2 U4456 ( .A(n4110), .ZN(n4114) );
  INV_X2 U4457 ( .A(net299240), .ZN(net295934) );
  NAND2_X2 U4469 ( .A1(n3664), .A2(n3665), .ZN(n4275) );
  XNOR2_X1 U4482 ( .A(n4076), .B(n1261), .ZN(n4281) );
  INV_X8 U4486 ( .A(net294790), .ZN(net294787) );
  INV_X4 U4495 ( .A(net295733), .ZN(n4276) );
  INV_X4 U4509 ( .A(net295626), .ZN(net295733) );
  OAI21_X1 U4510 ( .B1(net298860), .B2(net294048), .A(net295587), .ZN(n3186)
         );
  INV_X8 U4528 ( .A(net294995), .ZN(net294940) );
  BUF_X4 U4534 ( .A(n4284), .Z(n1240) );
  INV_X1 U4551 ( .A(n3764), .ZN(n3762) );
  NOR2_X4 U4559 ( .A1(n3324), .A2(n3323), .ZN(n4277) );
  INV_X4 U4566 ( .A(n4277), .ZN(n3511) );
  INV_X2 U4597 ( .A(net294535), .ZN(n4278) );
  INV_X4 U4609 ( .A(n4278), .ZN(n4279) );
  NAND2_X4 U4611 ( .A1(n3363), .A2(n3362), .ZN(n3571) );
  BUF_X8 U4642 ( .A(n4108), .Z(n4280) );
  NAND2_X4 U4643 ( .A1(n2288), .A2(n2400), .ZN(n2289) );
  AND2_X2 U4673 ( .A1(n3633), .A2(n3625), .ZN(n1563) );
  NAND2_X1 U4692 ( .A1(net297196), .A2(n3625), .ZN(n3567) );
  INV_X8 U4709 ( .A(n3028), .ZN(n3029) );
  NAND2_X2 U4710 ( .A1(n2745), .A2(n2619), .ZN(n1329) );
  INV_X4 U4722 ( .A(n3106), .ZN(n3108) );
  NAND2_X2 U4723 ( .A1(n2397), .A2(n1503), .ZN(n2355) );
  INV_X8 U4734 ( .A(n3503), .ZN(n3577) );
  INV_X2 U4783 ( .A(n3481), .ZN(n3480) );
  NAND3_X1 U4784 ( .A1(n2188), .A2(n2187), .A3(n2186), .ZN(n1503) );
  INV_X1 U4785 ( .A(net296771), .ZN(net298605) );
  INV_X2 U4786 ( .A(net296329), .ZN(net296425) );
  INV_X4 U4787 ( .A(net296329), .ZN(n1346) );
  INV_X4 U4788 ( .A(net297484), .ZN(net298051) );
  NAND2_X4 U4789 ( .A1(n2556), .A2(n2557), .ZN(n2558) );
  INV_X4 U4790 ( .A(n1914), .ZN(n1739) );
  INV_X1 U4791 ( .A(n1510), .ZN(n1511) );
  OAI211_X2 U4792 ( .C1(n1381), .C2(n3599), .A(n3598), .B(net294913), .ZN(
        n4283) );
  NAND3_X4 U4793 ( .A1(a[20]), .A2(net295008), .A3(net297226), .ZN(net294913)
         );
  NAND2_X2 U4794 ( .A1(n3265), .A2(n3266), .ZN(n4284) );
  INV_X8 U4795 ( .A(n3267), .ZN(n3265) );
  NOR2_X4 U4796 ( .A1(n1788), .A2(n1690), .ZN(n2905) );
  INV_X8 U4797 ( .A(net294044), .ZN(n4285) );
  INV_X8 U4798 ( .A(net294329), .ZN(net294044) );
  NAND2_X4 U4799 ( .A1(net294438), .A2(net294406), .ZN(net294532) );
  INV_X4 U4800 ( .A(n3579), .ZN(n1513) );
  NOR2_X2 U4801 ( .A1(n3107), .A2(n3106), .ZN(n3112) );
  NAND2_X1 U4802 ( .A1(n1521), .A2(n3490), .ZN(n3372) );
  NAND2_X4 U4803 ( .A1(n1149), .A2(n1222), .ZN(n3626) );
  INV_X4 U4804 ( .A(n4287), .ZN(n4288) );
  NAND2_X1 U4805 ( .A1(n3244), .A2(net298655), .ZN(n3245) );
  INV_X8 U4806 ( .A(n3710), .ZN(n3785) );
  OAI21_X4 U4807 ( .B1(n2185), .B2(n2152), .A(n4256), .ZN(n2153) );
  NAND2_X4 U4808 ( .A1(n3686), .A2(n3685), .ZN(n3728) );
  INV_X2 U4809 ( .A(n3732), .ZN(n3733) );
  INV_X8 U4810 ( .A(n2312), .ZN(n2313) );
  INV_X2 U4811 ( .A(n3333), .ZN(n3391) );
  XNOR2_X1 U4812 ( .A(net294401), .B(net294402), .ZN(net299052) );
  INV_X2 U4813 ( .A(n4274), .ZN(n4038) );
  NAND2_X4 U4814 ( .A1(n3416), .A2(n3415), .ZN(n4289) );
  INV_X8 U4815 ( .A(n1588), .ZN(n3416) );
  INV_X8 U4816 ( .A(n3559), .ZN(n3627) );
  NAND2_X4 U4817 ( .A1(n3631), .A2(n3471), .ZN(n3559) );
  INV_X4 U4818 ( .A(n3272), .ZN(n3301) );
  NAND2_X4 U4819 ( .A1(n1609), .A2(n1163), .ZN(n2315) );
  CLKBUF_X3 U4820 ( .A(n3518), .Z(n4291) );
  NAND3_X2 U4821 ( .A1(n2687), .A2(n1629), .A3(n2686), .ZN(n2691) );
  INV_X2 U4822 ( .A(n1128), .ZN(n1422) );
  AOI22_X1 U4823 ( .A1(n3297), .A2(n2648), .B1(n2648), .B2(net297188), .ZN(
        n4292) );
  NAND2_X2 U4824 ( .A1(n3564), .A2(n3424), .ZN(n4293) );
  INV_X32 U4825 ( .A(control[1]), .ZN(net297170) );
  INV_X4 U4826 ( .A(n1393), .ZN(n1388) );
  NAND2_X4 U4827 ( .A1(n3727), .A2(n3800), .ZN(net294790) );
  XNOR2_X2 U4828 ( .A(n4294), .B(n1657), .ZN(n4030) );
  INV_X32 U4829 ( .A(n4101), .ZN(n4294) );
  NAND3_X2 U4830 ( .A1(n2133), .A2(n2135), .A3(n2134), .ZN(n2237) );
  OAI21_X4 U4831 ( .B1(n3648), .B2(n4295), .A(n3646), .ZN(n3653) );
  INV_X1 U4832 ( .A(n3588), .ZN(n4295) );
  INV_X8 U4833 ( .A(n3645), .ZN(n3648) );
  AOI22_X2 U4834 ( .A1(n4296), .A2(n1984), .B1(n4297), .B2(n1982), .ZN(n1991)
         );
  INV_X1 U4835 ( .A(n1879), .ZN(n4296) );
  INV_X2 U4836 ( .A(n2115), .ZN(n4297) );
  NAND3_X4 U4837 ( .A1(n3286), .A2(n3285), .A3(n3284), .ZN(n1244) );
  NAND2_X4 U4838 ( .A1(n1522), .A2(n3166), .ZN(n3382) );
  NOR2_X4 U4839 ( .A1(net294779), .A2(n4298), .ZN(n4299) );
  INV_X4 U4840 ( .A(n3536), .ZN(n4298) );
  INV_X4 U4841 ( .A(n4299), .ZN(n3537) );
  AOI21_X4 U4842 ( .B1(n1210), .B2(n1211), .A(n3151), .ZN(n4300) );
  INV_X8 U4843 ( .A(n4300), .ZN(n3400) );
  INV_X2 U4844 ( .A(n3157), .ZN(n3330) );
  NOR2_X4 U4845 ( .A1(net294580), .A2(n4301), .ZN(n4302) );
  INV_X2 U4846 ( .A(net294640), .ZN(n4301) );
  INV_X4 U4847 ( .A(n4302), .ZN(net294577) );
  OAI21_X4 U4848 ( .B1(n4001), .B2(n4303), .A(n3999), .ZN(n4022) );
  INV_X2 U4849 ( .A(n3967), .ZN(n4303) );
  NAND2_X4 U4850 ( .A1(n2738), .A2(n2627), .ZN(n2537) );
  NAND3_X2 U4851 ( .A1(n1685), .A2(n1686), .A3(n2784), .ZN(n2852) );
  OAI21_X2 U4852 ( .B1(n1520), .B2(net294048), .A(n3360), .ZN(n3361) );
  NAND2_X4 U4853 ( .A1(n3404), .A2(n1645), .ZN(n1254) );
  INV_X4 U4854 ( .A(n3403), .ZN(n3404) );
  NOR3_X4 U4855 ( .A1(net297170), .A2(n1786), .A3(control[0]), .ZN(n1785) );
  XNOR2_X2 U4856 ( .A(n4082), .B(n4083), .ZN(n4084) );
  OAI21_X4 U4857 ( .B1(n2741), .B2(n2742), .A(n2917), .ZN(n2668) );
  XNOR2_X2 U4858 ( .A(n1811), .B(n1812), .ZN(n1818) );
  OAI221_X4 U4859 ( .B1(n3076), .B2(n3116), .C1(n3075), .C2(n3074), .A(n3073), 
        .ZN(n3077) );
  INV_X4 U4860 ( .A(n3312), .ZN(n3076) );
  OAI21_X4 U4861 ( .B1(n3463), .B2(n4304), .A(n3570), .ZN(n3310) );
  INV_X1 U4862 ( .A(n3374), .ZN(n4304) );
endmodule

