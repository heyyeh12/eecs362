
module and_32 ( a, b, z );
  input [31:0] a;
  input [31:0] b;
  output [31:0] z;


  AND2_X2 U1 ( .A1(b[9]), .A2(a[9]), .ZN(z[9]) );
  AND2_X2 U2 ( .A1(b[8]), .A2(a[8]), .ZN(z[8]) );
  AND2_X2 U3 ( .A1(b[7]), .A2(a[7]), .ZN(z[7]) );
  AND2_X2 U4 ( .A1(b[6]), .A2(a[6]), .ZN(z[6]) );
  AND2_X2 U5 ( .A1(b[5]), .A2(a[5]), .ZN(z[5]) );
  AND2_X2 U6 ( .A1(b[4]), .A2(a[4]), .ZN(z[4]) );
  AND2_X2 U7 ( .A1(b[3]), .A2(a[3]), .ZN(z[3]) );
  AND2_X2 U8 ( .A1(b[31]), .A2(a[31]), .ZN(z[31]) );
  AND2_X2 U9 ( .A1(b[30]), .A2(a[30]), .ZN(z[30]) );
  AND2_X2 U10 ( .A1(b[2]), .A2(a[2]), .ZN(z[2]) );
  AND2_X2 U11 ( .A1(b[29]), .A2(a[29]), .ZN(z[29]) );
  AND2_X2 U12 ( .A1(b[28]), .A2(a[28]), .ZN(z[28]) );
  AND2_X2 U13 ( .A1(b[27]), .A2(a[27]), .ZN(z[27]) );
  AND2_X2 U14 ( .A1(b[26]), .A2(a[26]), .ZN(z[26]) );
  AND2_X2 U15 ( .A1(b[25]), .A2(a[25]), .ZN(z[25]) );
  AND2_X2 U16 ( .A1(b[24]), .A2(a[24]), .ZN(z[24]) );
  AND2_X2 U17 ( .A1(b[23]), .A2(a[23]), .ZN(z[23]) );
  AND2_X2 U18 ( .A1(b[22]), .A2(a[22]), .ZN(z[22]) );
  AND2_X2 U19 ( .A1(b[21]), .A2(a[21]), .ZN(z[21]) );
  AND2_X2 U20 ( .A1(b[20]), .A2(a[20]), .ZN(z[20]) );
  AND2_X2 U21 ( .A1(b[1]), .A2(a[1]), .ZN(z[1]) );
  AND2_X2 U22 ( .A1(b[19]), .A2(a[19]), .ZN(z[19]) );
  AND2_X2 U23 ( .A1(b[18]), .A2(a[18]), .ZN(z[18]) );
  AND2_X2 U24 ( .A1(b[17]), .A2(a[17]), .ZN(z[17]) );
  AND2_X2 U25 ( .A1(b[16]), .A2(a[16]), .ZN(z[16]) );
  AND2_X2 U26 ( .A1(b[15]), .A2(a[15]), .ZN(z[15]) );
  AND2_X2 U27 ( .A1(b[14]), .A2(a[14]), .ZN(z[14]) );
  AND2_X2 U28 ( .A1(b[13]), .A2(a[13]), .ZN(z[13]) );
  AND2_X2 U29 ( .A1(b[12]), .A2(a[12]), .ZN(z[12]) );
  AND2_X2 U30 ( .A1(b[11]), .A2(a[11]), .ZN(z[11]) );
  AND2_X2 U31 ( .A1(b[10]), .A2(a[10]), .ZN(z[10]) );
  AND2_X2 U32 ( .A1(b[0]), .A2(a[0]), .ZN(z[0]) );
endmodule

