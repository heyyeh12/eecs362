
module mem_wb ( clk, rst, ctrl, valid_d, instr_d, regDst_d, memRd_d, regWr_d, 
        link_d, fp_d, dSize_d, rd_d, aluRes_d, memRdData_d, reg31Val_d, 
        busFP_d, busA_d, instr_q, regDst_q, memRd_q, regWr_q, link_q, fp_q, 
        dSize_q, rd_q, aluRes_q, memRdData_q, reg31Val_q, busFP_q, busA_q, 
        valid_q );
  input [1:0] ctrl;
  input [31:0] instr_d;
  input [1:0] dSize_d;
  input [4:0] rd_d;
  input [31:0] aluRes_d;
  input [31:0] memRdData_d;
  input [31:0] reg31Val_d;
  input [31:0] busFP_d;
  input [31:0] busA_d;
  output [31:0] instr_q;
  output [1:0] dSize_q;
  output [4:0] rd_q;
  output [31:0] aluRes_q;
  output [31:0] memRdData_q;
  output [31:0] reg31Val_q;
  output [31:0] busFP_q;
  output [31:0] busA_q;
  input clk, rst, valid_d, regDst_d, memRd_d, regWr_d, link_d, fp_d;
  output regDst_q, memRd_q, regWr_q, link_q, fp_q, valid_q;
  wire   n1, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309;

  DFF_X1 memRdData_q_reg_31_ ( .D(n289), .CK(clk), .Q(memRdData_q[31]) );
  DFF_X1 memRdData_q_reg_30_ ( .D(n288), .CK(clk), .Q(memRdData_q[30]) );
  DFF_X1 memRdData_q_reg_29_ ( .D(n287), .CK(clk), .Q(memRdData_q[29]) );
  DFF_X1 memRdData_q_reg_28_ ( .D(n286), .CK(clk), .Q(memRdData_q[28]) );
  DFF_X1 memRdData_q_reg_27_ ( .D(n285), .CK(clk), .Q(memRdData_q[27]) );
  DFF_X1 memRdData_q_reg_26_ ( .D(n284), .CK(clk), .Q(memRdData_q[26]) );
  DFF_X1 memRdData_q_reg_25_ ( .D(n283), .CK(clk), .Q(memRdData_q[25]) );
  DFF_X1 memRdData_q_reg_24_ ( .D(n282), .CK(clk), .Q(memRdData_q[24]) );
  DFF_X1 memRdData_q_reg_23_ ( .D(n281), .CK(clk), .Q(memRdData_q[23]) );
  DFF_X1 memRdData_q_reg_22_ ( .D(n280), .CK(clk), .Q(memRdData_q[22]) );
  DFF_X1 memRdData_q_reg_21_ ( .D(n279), .CK(clk), .Q(memRdData_q[21]) );
  DFF_X1 memRdData_q_reg_20_ ( .D(n278), .CK(clk), .Q(memRdData_q[20]) );
  DFF_X1 memRdData_q_reg_19_ ( .D(n277), .CK(clk), .Q(memRdData_q[19]) );
  DFF_X1 memRdData_q_reg_18_ ( .D(n276), .CK(clk), .Q(memRdData_q[18]) );
  DFF_X1 memRdData_q_reg_17_ ( .D(n275), .CK(clk), .Q(memRdData_q[17]) );
  DFF_X1 memRdData_q_reg_16_ ( .D(n274), .CK(clk), .Q(memRdData_q[16]) );
  DFF_X1 memRdData_q_reg_15_ ( .D(n273), .CK(clk), .Q(memRdData_q[15]) );
  DFF_X1 memRdData_q_reg_14_ ( .D(n272), .CK(clk), .Q(memRdData_q[14]) );
  DFF_X1 memRdData_q_reg_13_ ( .D(n271), .CK(clk), .Q(memRdData_q[13]) );
  DFF_X1 memRdData_q_reg_12_ ( .D(n270), .CK(clk), .Q(memRdData_q[12]) );
  DFF_X1 memRdData_q_reg_11_ ( .D(n269), .CK(clk), .Q(memRdData_q[11]) );
  DFF_X1 memRdData_q_reg_10_ ( .D(n268), .CK(clk), .Q(memRdData_q[10]) );
  DFF_X1 memRdData_q_reg_9_ ( .D(n267), .CK(clk), .Q(memRdData_q[9]) );
  DFF_X1 memRdData_q_reg_8_ ( .D(n266), .CK(clk), .Q(memRdData_q[8]) );
  DFF_X1 memRdData_q_reg_7_ ( .D(n265), .CK(clk), .Q(memRdData_q[7]) );
  DFF_X1 memRdData_q_reg_6_ ( .D(n264), .CK(clk), .Q(memRdData_q[6]) );
  DFF_X1 memRdData_q_reg_5_ ( .D(n263), .CK(clk), .Q(memRdData_q[5]) );
  DFF_X1 memRdData_q_reg_4_ ( .D(n262), .CK(clk), .Q(memRdData_q[4]) );
  DFF_X1 memRdData_q_reg_3_ ( .D(n261), .CK(clk), .Q(memRdData_q[3]) );
  DFF_X1 memRdData_q_reg_2_ ( .D(n260), .CK(clk), .Q(memRdData_q[2]) );
  DFF_X1 memRdData_q_reg_1_ ( .D(n259), .CK(clk), .Q(memRdData_q[1]) );
  DFF_X1 memRdData_q_reg_0_ ( .D(n258), .CK(clk), .Q(memRdData_q[0]) );
  DFF_X1 reg31Val_q_reg_31_ ( .D(n257), .CK(clk), .Q(reg31Val_q[31]) );
  DFF_X1 reg31Val_q_reg_30_ ( .D(n256), .CK(clk), .Q(reg31Val_q[30]) );
  DFF_X1 reg31Val_q_reg_29_ ( .D(n255), .CK(clk), .Q(reg31Val_q[29]) );
  DFF_X1 reg31Val_q_reg_28_ ( .D(n254), .CK(clk), .Q(reg31Val_q[28]) );
  DFF_X1 reg31Val_q_reg_27_ ( .D(n253), .CK(clk), .Q(reg31Val_q[27]) );
  DFF_X1 reg31Val_q_reg_26_ ( .D(n252), .CK(clk), .Q(reg31Val_q[26]) );
  DFF_X1 reg31Val_q_reg_25_ ( .D(n251), .CK(clk), .Q(reg31Val_q[25]) );
  DFF_X1 reg31Val_q_reg_24_ ( .D(n250), .CK(clk), .Q(reg31Val_q[24]) );
  DFF_X1 reg31Val_q_reg_23_ ( .D(n249), .CK(clk), .Q(reg31Val_q[23]) );
  DFF_X1 reg31Val_q_reg_22_ ( .D(n248), .CK(clk), .Q(reg31Val_q[22]) );
  DFF_X1 reg31Val_q_reg_21_ ( .D(n247), .CK(clk), .Q(reg31Val_q[21]) );
  DFF_X1 reg31Val_q_reg_20_ ( .D(n246), .CK(clk), .Q(reg31Val_q[20]) );
  DFF_X1 reg31Val_q_reg_19_ ( .D(n245), .CK(clk), .Q(reg31Val_q[19]) );
  DFF_X1 reg31Val_q_reg_18_ ( .D(n244), .CK(clk), .Q(reg31Val_q[18]) );
  DFF_X1 reg31Val_q_reg_17_ ( .D(n243), .CK(clk), .Q(reg31Val_q[17]) );
  DFF_X1 reg31Val_q_reg_16_ ( .D(n242), .CK(clk), .Q(reg31Val_q[16]) );
  DFF_X1 reg31Val_q_reg_15_ ( .D(n241), .CK(clk), .Q(reg31Val_q[15]) );
  DFF_X1 reg31Val_q_reg_14_ ( .D(n240), .CK(clk), .Q(reg31Val_q[14]) );
  DFF_X1 reg31Val_q_reg_13_ ( .D(n239), .CK(clk), .Q(reg31Val_q[13]) );
  DFF_X1 reg31Val_q_reg_12_ ( .D(n238), .CK(clk), .Q(reg31Val_q[12]) );
  DFF_X1 reg31Val_q_reg_11_ ( .D(n237), .CK(clk), .Q(reg31Val_q[11]) );
  DFF_X1 reg31Val_q_reg_10_ ( .D(n236), .CK(clk), .Q(reg31Val_q[10]) );
  DFF_X1 reg31Val_q_reg_9_ ( .D(n235), .CK(clk), .Q(reg31Val_q[9]) );
  DFF_X1 reg31Val_q_reg_8_ ( .D(n234), .CK(clk), .Q(reg31Val_q[8]) );
  DFF_X1 reg31Val_q_reg_7_ ( .D(n233), .CK(clk), .Q(reg31Val_q[7]) );
  DFF_X1 reg31Val_q_reg_6_ ( .D(n232), .CK(clk), .Q(reg31Val_q[6]) );
  DFF_X1 reg31Val_q_reg_5_ ( .D(n231), .CK(clk), .Q(reg31Val_q[5]) );
  DFF_X1 reg31Val_q_reg_4_ ( .D(n230), .CK(clk), .Q(reg31Val_q[4]) );
  DFF_X1 reg31Val_q_reg_3_ ( .D(n229), .CK(clk), .Q(reg31Val_q[3]) );
  DFF_X1 reg31Val_q_reg_2_ ( .D(n228), .CK(clk), .Q(reg31Val_q[2]) );
  DFF_X1 reg31Val_q_reg_1_ ( .D(n227), .CK(clk), .Q(reg31Val_q[1]) );
  DFF_X1 reg31Val_q_reg_0_ ( .D(n226), .CK(clk), .Q(reg31Val_q[0]) );
  DFF_X1 link_q_reg ( .D(n225), .CK(clk), .Q(link_q) );
  DFFR_X1 instr_q_reg_31_ ( .D(n224), .CK(clk), .RN(rst), .Q(instr_q[31]) );
  DFFR_X1 instr_q_reg_30_ ( .D(n223), .CK(clk), .RN(rst), .Q(instr_q[30]) );
  DFFR_X1 instr_q_reg_29_ ( .D(n222), .CK(clk), .RN(rst), .Q(instr_q[29]) );
  DFFR_X1 instr_q_reg_28_ ( .D(n221), .CK(clk), .RN(rst), .Q(instr_q[28]) );
  DFFR_X1 instr_q_reg_27_ ( .D(n220), .CK(clk), .RN(rst), .Q(instr_q[27]) );
  DFFR_X1 instr_q_reg_26_ ( .D(n219), .CK(clk), .RN(rst), .Q(instr_q[26]) );
  DFFR_X1 instr_q_reg_25_ ( .D(n218), .CK(clk), .RN(rst), .Q(instr_q[25]) );
  DFFR_X1 instr_q_reg_24_ ( .D(n217), .CK(clk), .RN(rst), .Q(instr_q[24]) );
  DFFR_X1 instr_q_reg_23_ ( .D(n216), .CK(clk), .RN(rst), .Q(instr_q[23]) );
  DFFR_X1 instr_q_reg_22_ ( .D(n215), .CK(clk), .RN(rst), .Q(instr_q[22]) );
  DFFR_X1 instr_q_reg_21_ ( .D(n214), .CK(clk), .RN(rst), .Q(instr_q[21]) );
  DFFR_X1 instr_q_reg_20_ ( .D(n213), .CK(clk), .RN(rst), .Q(instr_q[20]) );
  DFFR_X1 instr_q_reg_19_ ( .D(n212), .CK(clk), .RN(rst), .Q(instr_q[19]) );
  DFFR_X1 instr_q_reg_18_ ( .D(n211), .CK(clk), .RN(rst), .Q(instr_q[18]) );
  DFFR_X1 instr_q_reg_17_ ( .D(n210), .CK(clk), .RN(rst), .Q(instr_q[17]) );
  DFFR_X1 instr_q_reg_16_ ( .D(n209), .CK(clk), .RN(rst), .Q(instr_q[16]) );
  DFFR_X1 instr_q_reg_15_ ( .D(n208), .CK(clk), .RN(rst), .Q(instr_q[15]) );
  DFFR_X1 instr_q_reg_14_ ( .D(n207), .CK(clk), .RN(rst), .Q(instr_q[14]) );
  DFFR_X1 instr_q_reg_13_ ( .D(n206), .CK(clk), .RN(rst), .Q(instr_q[13]) );
  DFFR_X1 instr_q_reg_12_ ( .D(n205), .CK(clk), .RN(rst), .Q(instr_q[12]) );
  DFFR_X1 instr_q_reg_11_ ( .D(n204), .CK(clk), .RN(rst), .Q(instr_q[11]) );
  DFFR_X1 instr_q_reg_10_ ( .D(n203), .CK(clk), .RN(rst), .Q(instr_q[10]) );
  DFFR_X1 instr_q_reg_9_ ( .D(n202), .CK(clk), .RN(rst), .Q(instr_q[9]) );
  DFFR_X1 instr_q_reg_8_ ( .D(n201), .CK(clk), .RN(rst), .Q(instr_q[8]) );
  DFFR_X1 instr_q_reg_7_ ( .D(n200), .CK(clk), .RN(rst), .Q(instr_q[7]) );
  DFFR_X1 instr_q_reg_6_ ( .D(n199), .CK(clk), .RN(rst), .Q(instr_q[6]) );
  DFFR_X1 instr_q_reg_5_ ( .D(n198), .CK(clk), .RN(rst), .Q(instr_q[5]) );
  DFFS_X1 instr_q_reg_4_ ( .D(n197), .CK(clk), .SN(rst), .Q(instr_q[4]) );
  DFFR_X1 instr_q_reg_3_ ( .D(n196), .CK(clk), .RN(rst), .Q(instr_q[3]) );
  DFFS_X1 instr_q_reg_2_ ( .D(n195), .CK(clk), .SN(rst), .Q(instr_q[2]) );
  DFFR_X1 instr_q_reg_1_ ( .D(n194), .CK(clk), .RN(rst), .Q(instr_q[1]) );
  DFFS_X1 instr_q_reg_0_ ( .D(n193), .CK(clk), .SN(rst), .Q(instr_q[0]) );
  DFFR_X1 regWr_q_reg ( .D(n192), .CK(clk), .RN(rst), .Q(regWr_q) );
  DFFR_X1 valid_q_reg ( .D(n191), .CK(clk), .RN(rst), .Q(valid_q) );
  DFF_X1 fp_q_reg ( .D(n190), .CK(clk), .Q(fp_q) );
  DFF_X1 regDst_q_reg ( .D(n189), .CK(clk), .Q(regDst_q) );
  DFF_X1 memRd_q_reg ( .D(n188), .CK(clk), .Q(memRd_q) );
  DFF_X1 dSize_q_reg_1_ ( .D(n187), .CK(clk), .Q(dSize_q[1]) );
  DFF_X1 dSize_q_reg_0_ ( .D(n186), .CK(clk), .Q(dSize_q[0]) );
  DFF_X1 rd_q_reg_4_ ( .D(n185), .CK(clk), .Q(rd_q[4]) );
  DFF_X1 rd_q_reg_3_ ( .D(n184), .CK(clk), .Q(rd_q[3]) );
  DFF_X1 rd_q_reg_2_ ( .D(n183), .CK(clk), .Q(rd_q[2]) );
  DFF_X1 rd_q_reg_1_ ( .D(n182), .CK(clk), .Q(rd_q[1]) );
  DFF_X1 rd_q_reg_0_ ( .D(n181), .CK(clk), .Q(rd_q[0]) );
  DFF_X1 aluRes_q_reg_31_ ( .D(n180), .CK(clk), .Q(aluRes_q[31]) );
  DFF_X1 aluRes_q_reg_30_ ( .D(n179), .CK(clk), .Q(aluRes_q[30]) );
  DFF_X1 aluRes_q_reg_29_ ( .D(n178), .CK(clk), .Q(aluRes_q[29]) );
  DFF_X1 aluRes_q_reg_28_ ( .D(n177), .CK(clk), .Q(aluRes_q[28]) );
  DFF_X1 aluRes_q_reg_27_ ( .D(n176), .CK(clk), .Q(aluRes_q[27]) );
  DFF_X1 aluRes_q_reg_26_ ( .D(n175), .CK(clk), .Q(aluRes_q[26]) );
  DFF_X1 aluRes_q_reg_25_ ( .D(n174), .CK(clk), .Q(aluRes_q[25]) );
  DFF_X1 aluRes_q_reg_24_ ( .D(n173), .CK(clk), .Q(aluRes_q[24]) );
  DFF_X1 aluRes_q_reg_23_ ( .D(n172), .CK(clk), .Q(aluRes_q[23]) );
  DFF_X1 aluRes_q_reg_22_ ( .D(n171), .CK(clk), .Q(aluRes_q[22]) );
  DFF_X1 aluRes_q_reg_21_ ( .D(n170), .CK(clk), .Q(aluRes_q[21]) );
  DFF_X1 aluRes_q_reg_20_ ( .D(n169), .CK(clk), .Q(aluRes_q[20]) );
  DFF_X1 aluRes_q_reg_19_ ( .D(n168), .CK(clk), .Q(aluRes_q[19]) );
  DFF_X1 aluRes_q_reg_18_ ( .D(n167), .CK(clk), .Q(aluRes_q[18]) );
  DFF_X1 aluRes_q_reg_17_ ( .D(n166), .CK(clk), .Q(aluRes_q[17]) );
  DFF_X1 aluRes_q_reg_16_ ( .D(n165), .CK(clk), .Q(aluRes_q[16]) );
  DFF_X1 aluRes_q_reg_15_ ( .D(n164), .CK(clk), .Q(aluRes_q[15]) );
  DFF_X1 aluRes_q_reg_14_ ( .D(n163), .CK(clk), .Q(aluRes_q[14]) );
  DFF_X1 aluRes_q_reg_13_ ( .D(n162), .CK(clk), .Q(aluRes_q[13]) );
  DFF_X1 aluRes_q_reg_12_ ( .D(n161), .CK(clk), .Q(aluRes_q[12]) );
  DFF_X1 aluRes_q_reg_11_ ( .D(n160), .CK(clk), .Q(aluRes_q[11]) );
  DFF_X1 aluRes_q_reg_10_ ( .D(n159), .CK(clk), .Q(aluRes_q[10]) );
  DFF_X1 aluRes_q_reg_9_ ( .D(n158), .CK(clk), .Q(aluRes_q[9]) );
  DFF_X1 aluRes_q_reg_8_ ( .D(n157), .CK(clk), .Q(aluRes_q[8]) );
  DFF_X1 aluRes_q_reg_7_ ( .D(n156), .CK(clk), .Q(aluRes_q[7]) );
  DFF_X1 aluRes_q_reg_6_ ( .D(n155), .CK(clk), .Q(aluRes_q[6]) );
  DFF_X1 aluRes_q_reg_5_ ( .D(n154), .CK(clk), .Q(aluRes_q[5]) );
  DFF_X1 aluRes_q_reg_4_ ( .D(n153), .CK(clk), .Q(aluRes_q[4]) );
  DFF_X1 aluRes_q_reg_3_ ( .D(n152), .CK(clk), .Q(aluRes_q[3]) );
  DFF_X1 aluRes_q_reg_2_ ( .D(n151), .CK(clk), .Q(aluRes_q[2]) );
  DFF_X1 aluRes_q_reg_1_ ( .D(n150), .CK(clk), .Q(aluRes_q[1]) );
  DFF_X1 aluRes_q_reg_0_ ( .D(n149), .CK(clk), .Q(aluRes_q[0]) );
  INV_X1 U3 ( .A(n1), .ZN(n191) );
  AOI22_X1 U4 ( .A1(valid_d), .A2(n309), .B1(valid_q), .B2(n308), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n192) );
  AOI22_X1 U6 ( .A1(regWr_d), .A2(n309), .B1(regWr_q), .B2(n3), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n189) );
  AOI22_X1 U8 ( .A1(regDst_q), .A2(n302), .B1(regDst_d), .B2(n295), .ZN(n5) );
  INV_X1 U9 ( .A(n8), .ZN(n235) );
  AOI22_X1 U10 ( .A1(reg31Val_q[9]), .A2(n303), .B1(reg31Val_d[9]), .B2(n295), 
        .ZN(n8) );
  INV_X1 U11 ( .A(n9), .ZN(n234) );
  AOI22_X1 U12 ( .A1(reg31Val_q[8]), .A2(n302), .B1(reg31Val_d[8]), .B2(n296), 
        .ZN(n9) );
  INV_X1 U13 ( .A(n10), .ZN(n233) );
  AOI22_X1 U14 ( .A1(reg31Val_q[7]), .A2(n303), .B1(reg31Val_d[7]), .B2(n296), 
        .ZN(n10) );
  INV_X1 U15 ( .A(n11), .ZN(n232) );
  AOI22_X1 U16 ( .A1(reg31Val_q[6]), .A2(n302), .B1(reg31Val_d[6]), .B2(n295), 
        .ZN(n11) );
  INV_X1 U17 ( .A(n12), .ZN(n231) );
  AOI22_X1 U18 ( .A1(reg31Val_q[5]), .A2(n303), .B1(reg31Val_d[5]), .B2(n295), 
        .ZN(n12) );
  INV_X1 U19 ( .A(n13), .ZN(n230) );
  AOI22_X1 U20 ( .A1(reg31Val_q[4]), .A2(n302), .B1(reg31Val_d[4]), .B2(n296), 
        .ZN(n13) );
  INV_X1 U21 ( .A(n14), .ZN(n229) );
  AOI22_X1 U22 ( .A1(reg31Val_q[3]), .A2(n303), .B1(reg31Val_d[3]), .B2(n296), 
        .ZN(n14) );
  INV_X1 U23 ( .A(n15), .ZN(n257) );
  AOI22_X1 U24 ( .A1(reg31Val_q[31]), .A2(n303), .B1(reg31Val_d[31]), .B2(n296), .ZN(n15) );
  INV_X1 U25 ( .A(n16), .ZN(n256) );
  AOI22_X1 U26 ( .A1(reg31Val_q[30]), .A2(n303), .B1(reg31Val_d[30]), .B2(n296), .ZN(n16) );
  INV_X1 U27 ( .A(n17), .ZN(n228) );
  AOI22_X1 U28 ( .A1(reg31Val_q[2]), .A2(n303), .B1(reg31Val_d[2]), .B2(n296), 
        .ZN(n17) );
  INV_X1 U29 ( .A(n18), .ZN(n255) );
  AOI22_X1 U30 ( .A1(reg31Val_q[29]), .A2(n303), .B1(reg31Val_d[29]), .B2(n296), .ZN(n18) );
  INV_X1 U31 ( .A(n19), .ZN(n254) );
  AOI22_X1 U32 ( .A1(reg31Val_q[28]), .A2(n303), .B1(reg31Val_d[28]), .B2(n296), .ZN(n19) );
  INV_X1 U33 ( .A(n20), .ZN(n253) );
  AOI22_X1 U34 ( .A1(reg31Val_q[27]), .A2(n303), .B1(reg31Val_d[27]), .B2(n296), .ZN(n20) );
  INV_X1 U35 ( .A(n21), .ZN(n252) );
  AOI22_X1 U36 ( .A1(reg31Val_q[26]), .A2(n303), .B1(reg31Val_d[26]), .B2(n296), .ZN(n21) );
  INV_X1 U37 ( .A(n22), .ZN(n251) );
  AOI22_X1 U38 ( .A1(reg31Val_q[25]), .A2(n303), .B1(reg31Val_d[25]), .B2(n296), .ZN(n22) );
  INV_X1 U39 ( .A(n23), .ZN(n250) );
  AOI22_X1 U40 ( .A1(reg31Val_q[24]), .A2(n303), .B1(reg31Val_d[24]), .B2(n296), .ZN(n23) );
  INV_X1 U41 ( .A(n24), .ZN(n249) );
  AOI22_X1 U42 ( .A1(reg31Val_q[23]), .A2(n303), .B1(reg31Val_d[23]), .B2(n296), .ZN(n24) );
  INV_X1 U43 ( .A(n25), .ZN(n248) );
  AOI22_X1 U44 ( .A1(reg31Val_q[22]), .A2(n303), .B1(reg31Val_d[22]), .B2(n296), .ZN(n25) );
  INV_X1 U45 ( .A(n26), .ZN(n247) );
  AOI22_X1 U46 ( .A1(reg31Val_q[21]), .A2(n303), .B1(reg31Val_d[21]), .B2(n295), .ZN(n26) );
  INV_X1 U47 ( .A(n27), .ZN(n246) );
  AOI22_X1 U48 ( .A1(reg31Val_q[20]), .A2(n303), .B1(reg31Val_d[20]), .B2(n295), .ZN(n27) );
  INV_X1 U49 ( .A(n28), .ZN(n227) );
  AOI22_X1 U50 ( .A1(reg31Val_q[1]), .A2(n303), .B1(reg31Val_d[1]), .B2(n295), 
        .ZN(n28) );
  INV_X1 U51 ( .A(n29), .ZN(n245) );
  AOI22_X1 U52 ( .A1(reg31Val_q[19]), .A2(n303), .B1(reg31Val_d[19]), .B2(n295), .ZN(n29) );
  INV_X1 U53 ( .A(n30), .ZN(n244) );
  AOI22_X1 U54 ( .A1(reg31Val_q[18]), .A2(n303), .B1(reg31Val_d[18]), .B2(n295), .ZN(n30) );
  INV_X1 U55 ( .A(n31), .ZN(n243) );
  AOI22_X1 U56 ( .A1(reg31Val_q[17]), .A2(n303), .B1(reg31Val_d[17]), .B2(n295), .ZN(n31) );
  INV_X1 U57 ( .A(n32), .ZN(n242) );
  AOI22_X1 U58 ( .A1(reg31Val_q[16]), .A2(n303), .B1(reg31Val_d[16]), .B2(n295), .ZN(n32) );
  INV_X1 U59 ( .A(n33), .ZN(n241) );
  AOI22_X1 U60 ( .A1(reg31Val_q[15]), .A2(n303), .B1(reg31Val_d[15]), .B2(n295), .ZN(n33) );
  INV_X1 U61 ( .A(n34), .ZN(n240) );
  AOI22_X1 U62 ( .A1(reg31Val_q[14]), .A2(n303), .B1(reg31Val_d[14]), .B2(n295), .ZN(n34) );
  INV_X1 U63 ( .A(n35), .ZN(n239) );
  AOI22_X1 U64 ( .A1(reg31Val_q[13]), .A2(n303), .B1(reg31Val_d[13]), .B2(n295), .ZN(n35) );
  INV_X1 U65 ( .A(n36), .ZN(n238) );
  AOI22_X1 U66 ( .A1(reg31Val_q[12]), .A2(n303), .B1(reg31Val_d[12]), .B2(n295), .ZN(n36) );
  INV_X1 U67 ( .A(n37), .ZN(n237) );
  AOI22_X1 U68 ( .A1(reg31Val_q[11]), .A2(n303), .B1(reg31Val_d[11]), .B2(n294), .ZN(n37) );
  INV_X1 U69 ( .A(n38), .ZN(n236) );
  AOI22_X1 U70 ( .A1(reg31Val_q[10]), .A2(n303), .B1(reg31Val_d[10]), .B2(n293), .ZN(n38) );
  INV_X1 U71 ( .A(n39), .ZN(n226) );
  AOI22_X1 U72 ( .A1(reg31Val_q[0]), .A2(n303), .B1(reg31Val_d[0]), .B2(n294), 
        .ZN(n39) );
  INV_X1 U73 ( .A(n40), .ZN(n185) );
  AOI22_X1 U74 ( .A1(rd_q[4]), .A2(n303), .B1(rd_d[4]), .B2(n293), .ZN(n40) );
  INV_X1 U75 ( .A(n41), .ZN(n184) );
  AOI22_X1 U76 ( .A1(rd_q[3]), .A2(n302), .B1(rd_d[3]), .B2(n293), .ZN(n41) );
  INV_X1 U77 ( .A(n42), .ZN(n183) );
  AOI22_X1 U78 ( .A1(rd_q[2]), .A2(n302), .B1(rd_d[2]), .B2(n294), .ZN(n42) );
  INV_X1 U79 ( .A(n43), .ZN(n182) );
  AOI22_X1 U80 ( .A1(rd_q[1]), .A2(n302), .B1(rd_d[1]), .B2(n293), .ZN(n43) );
  INV_X1 U81 ( .A(n44), .ZN(n181) );
  AOI22_X1 U82 ( .A1(rd_q[0]), .A2(n302), .B1(rd_d[0]), .B2(n294), .ZN(n44) );
  INV_X1 U83 ( .A(n45), .ZN(n188) );
  AOI22_X1 U84 ( .A1(memRd_q), .A2(n302), .B1(memRd_d), .B2(n293), .ZN(n45) );
  INV_X1 U85 ( .A(n46), .ZN(n267) );
  AOI22_X1 U86 ( .A1(memRdData_q[9]), .A2(n302), .B1(memRdData_d[9]), .B2(n294), .ZN(n46) );
  INV_X1 U87 ( .A(n47), .ZN(n266) );
  AOI22_X1 U88 ( .A1(memRdData_q[8]), .A2(n302), .B1(memRdData_d[8]), .B2(n293), .ZN(n47) );
  INV_X1 U89 ( .A(n48), .ZN(n265) );
  AOI22_X1 U90 ( .A1(memRdData_q[7]), .A2(n302), .B1(memRdData_d[7]), .B2(n294), .ZN(n48) );
  INV_X1 U91 ( .A(n49), .ZN(n264) );
  AOI22_X1 U92 ( .A1(memRdData_q[6]), .A2(n302), .B1(memRdData_d[6]), .B2(n294), .ZN(n49) );
  INV_X1 U93 ( .A(n50), .ZN(n263) );
  AOI22_X1 U94 ( .A1(memRdData_q[5]), .A2(n302), .B1(memRdData_d[5]), .B2(n294), .ZN(n50) );
  INV_X1 U95 ( .A(n51), .ZN(n262) );
  AOI22_X1 U96 ( .A1(memRdData_q[4]), .A2(n302), .B1(memRdData_d[4]), .B2(n294), .ZN(n51) );
  INV_X1 U97 ( .A(n52), .ZN(n261) );
  AOI22_X1 U98 ( .A1(memRdData_q[3]), .A2(n302), .B1(memRdData_d[3]), .B2(n294), .ZN(n52) );
  INV_X1 U99 ( .A(n53), .ZN(n289) );
  AOI22_X1 U100 ( .A1(memRdData_q[31]), .A2(n302), .B1(memRdData_d[31]), .B2(
        n294), .ZN(n53) );
  INV_X1 U101 ( .A(n54), .ZN(n288) );
  AOI22_X1 U102 ( .A1(memRdData_q[30]), .A2(n302), .B1(memRdData_d[30]), .B2(
        n294), .ZN(n54) );
  INV_X1 U103 ( .A(n55), .ZN(n260) );
  AOI22_X1 U104 ( .A1(memRdData_q[2]), .A2(n302), .B1(memRdData_d[2]), .B2(
        n294), .ZN(n55) );
  INV_X1 U105 ( .A(n56), .ZN(n287) );
  AOI22_X1 U106 ( .A1(memRdData_q[29]), .A2(n302), .B1(memRdData_d[29]), .B2(
        n294), .ZN(n56) );
  INV_X1 U107 ( .A(n57), .ZN(n286) );
  AOI22_X1 U108 ( .A1(memRdData_q[28]), .A2(n302), .B1(memRdData_d[28]), .B2(
        n294), .ZN(n57) );
  INV_X1 U109 ( .A(n58), .ZN(n285) );
  AOI22_X1 U110 ( .A1(memRdData_q[27]), .A2(n302), .B1(memRdData_d[27]), .B2(
        n294), .ZN(n58) );
  INV_X1 U111 ( .A(n59), .ZN(n284) );
  AOI22_X1 U112 ( .A1(memRdData_q[26]), .A2(n302), .B1(memRdData_d[26]), .B2(
        n293), .ZN(n59) );
  INV_X1 U113 ( .A(n60), .ZN(n283) );
  AOI22_X1 U114 ( .A1(memRdData_q[25]), .A2(n302), .B1(memRdData_d[25]), .B2(
        n293), .ZN(n60) );
  INV_X1 U115 ( .A(n61), .ZN(n282) );
  AOI22_X1 U116 ( .A1(memRdData_q[24]), .A2(n302), .B1(memRdData_d[24]), .B2(
        n293), .ZN(n61) );
  INV_X1 U117 ( .A(n62), .ZN(n281) );
  AOI22_X1 U118 ( .A1(memRdData_q[23]), .A2(n302), .B1(memRdData_d[23]), .B2(
        n293), .ZN(n62) );
  INV_X1 U119 ( .A(n63), .ZN(n280) );
  AOI22_X1 U120 ( .A1(memRdData_q[22]), .A2(n302), .B1(memRdData_d[22]), .B2(
        n293), .ZN(n63) );
  INV_X1 U121 ( .A(n64), .ZN(n279) );
  AOI22_X1 U122 ( .A1(memRdData_q[21]), .A2(n302), .B1(memRdData_d[21]), .B2(
        n293), .ZN(n64) );
  INV_X1 U123 ( .A(n65), .ZN(n278) );
  AOI22_X1 U124 ( .A1(memRdData_q[20]), .A2(n302), .B1(memRdData_d[20]), .B2(
        n293), .ZN(n65) );
  INV_X1 U125 ( .A(n66), .ZN(n259) );
  AOI22_X1 U126 ( .A1(memRdData_q[1]), .A2(n302), .B1(memRdData_d[1]), .B2(
        n293), .ZN(n66) );
  INV_X1 U127 ( .A(n67), .ZN(n277) );
  AOI22_X1 U128 ( .A1(memRdData_q[19]), .A2(n302), .B1(memRdData_d[19]), .B2(
        n293), .ZN(n67) );
  INV_X1 U129 ( .A(n68), .ZN(n276) );
  AOI22_X1 U130 ( .A1(memRdData_q[18]), .A2(n301), .B1(memRdData_d[18]), .B2(
        n293), .ZN(n68) );
  INV_X1 U131 ( .A(n69), .ZN(n275) );
  AOI22_X1 U132 ( .A1(memRdData_q[17]), .A2(n301), .B1(memRdData_d[17]), .B2(
        n293), .ZN(n69) );
  INV_X1 U133 ( .A(n70), .ZN(n274) );
  AOI22_X1 U134 ( .A1(memRdData_q[16]), .A2(n301), .B1(memRdData_d[16]), .B2(
        n291), .ZN(n70) );
  INV_X1 U135 ( .A(n71), .ZN(n273) );
  AOI22_X1 U136 ( .A1(memRdData_q[15]), .A2(n301), .B1(memRdData_d[15]), .B2(
        n292), .ZN(n71) );
  INV_X1 U137 ( .A(n72), .ZN(n272) );
  AOI22_X1 U138 ( .A1(memRdData_q[14]), .A2(n301), .B1(memRdData_d[14]), .B2(
        n291), .ZN(n72) );
  INV_X1 U139 ( .A(n73), .ZN(n271) );
  AOI22_X1 U140 ( .A1(memRdData_q[13]), .A2(n301), .B1(memRdData_d[13]), .B2(
        n292), .ZN(n73) );
  INV_X1 U141 ( .A(n74), .ZN(n270) );
  AOI22_X1 U142 ( .A1(memRdData_q[12]), .A2(n301), .B1(memRdData_d[12]), .B2(
        n291), .ZN(n74) );
  INV_X1 U143 ( .A(n75), .ZN(n269) );
  AOI22_X1 U144 ( .A1(memRdData_q[11]), .A2(n301), .B1(memRdData_d[11]), .B2(
        n292), .ZN(n75) );
  INV_X1 U145 ( .A(n76), .ZN(n268) );
  AOI22_X1 U146 ( .A1(memRdData_q[10]), .A2(n301), .B1(memRdData_d[10]), .B2(
        n291), .ZN(n76) );
  INV_X1 U147 ( .A(n77), .ZN(n258) );
  AOI22_X1 U148 ( .A1(memRdData_q[0]), .A2(n301), .B1(memRdData_d[0]), .B2(
        n292), .ZN(n77) );
  INV_X1 U149 ( .A(n78), .ZN(n225) );
  AOI22_X1 U150 ( .A1(link_q), .A2(n301), .B1(link_d), .B2(n304), .ZN(n78) );
  INV_X1 U151 ( .A(n79), .ZN(n202) );
  AOI22_X1 U152 ( .A1(instr_d[9]), .A2(n309), .B1(instr_q[9]), .B2(n3), .ZN(
        n79) );
  INV_X1 U153 ( .A(n80), .ZN(n201) );
  AOI22_X1 U154 ( .A1(instr_d[8]), .A2(n309), .B1(instr_q[8]), .B2(n3), .ZN(
        n80) );
  INV_X1 U155 ( .A(n81), .ZN(n200) );
  AOI22_X1 U156 ( .A1(instr_d[7]), .A2(n309), .B1(instr_q[7]), .B2(n3), .ZN(
        n81) );
  INV_X1 U157 ( .A(n82), .ZN(n199) );
  AOI22_X1 U158 ( .A1(instr_d[6]), .A2(n309), .B1(instr_q[6]), .B2(n3), .ZN(
        n82) );
  INV_X1 U159 ( .A(n83), .ZN(n198) );
  AOI22_X1 U160 ( .A1(instr_d[5]), .A2(n309), .B1(instr_q[5]), .B2(n3), .ZN(
        n83) );
  INV_X1 U161 ( .A(n84), .ZN(n197) );
  AOI221_X1 U162 ( .B1(instr_q[4]), .B2(n308), .C1(instr_d[4]), .C2(n309), .A(
        n85), .ZN(n84) );
  INV_X1 U163 ( .A(n86), .ZN(n196) );
  AOI22_X1 U164 ( .A1(instr_d[3]), .A2(n309), .B1(instr_q[3]), .B2(n3), .ZN(
        n86) );
  INV_X1 U165 ( .A(n87), .ZN(n224) );
  AOI22_X1 U166 ( .A1(instr_d[31]), .A2(n309), .B1(instr_q[31]), .B2(n308), 
        .ZN(n87) );
  INV_X1 U167 ( .A(n88), .ZN(n223) );
  AOI22_X1 U168 ( .A1(instr_d[30]), .A2(n309), .B1(instr_q[30]), .B2(n3), .ZN(
        n88) );
  INV_X1 U169 ( .A(n89), .ZN(n195) );
  AOI221_X1 U170 ( .B1(instr_q[2]), .B2(n3), .C1(instr_d[2]), .C2(n309), .A(
        n85), .ZN(n89) );
  INV_X1 U171 ( .A(n90), .ZN(n222) );
  AOI22_X1 U172 ( .A1(instr_d[29]), .A2(n309), .B1(instr_q[29]), .B2(n308), 
        .ZN(n90) );
  INV_X1 U173 ( .A(n91), .ZN(n221) );
  AOI22_X1 U174 ( .A1(instr_d[28]), .A2(n309), .B1(instr_q[28]), .B2(n308), 
        .ZN(n91) );
  INV_X1 U175 ( .A(n92), .ZN(n220) );
  AOI22_X1 U176 ( .A1(instr_d[27]), .A2(n309), .B1(instr_q[27]), .B2(n308), 
        .ZN(n92) );
  INV_X1 U177 ( .A(n93), .ZN(n219) );
  AOI22_X1 U178 ( .A1(instr_d[26]), .A2(n309), .B1(instr_q[26]), .B2(n308), 
        .ZN(n93) );
  INV_X1 U179 ( .A(n94), .ZN(n218) );
  AOI22_X1 U180 ( .A1(instr_d[25]), .A2(n309), .B1(instr_q[25]), .B2(n308), 
        .ZN(n94) );
  INV_X1 U181 ( .A(n95), .ZN(n217) );
  AOI22_X1 U182 ( .A1(instr_d[24]), .A2(n309), .B1(instr_q[24]), .B2(n308), 
        .ZN(n95) );
  INV_X1 U183 ( .A(n96), .ZN(n216) );
  AOI22_X1 U184 ( .A1(instr_d[23]), .A2(n309), .B1(instr_q[23]), .B2(n308), 
        .ZN(n96) );
  INV_X1 U185 ( .A(n97), .ZN(n215) );
  AOI22_X1 U186 ( .A1(instr_d[22]), .A2(n309), .B1(instr_q[22]), .B2(n308), 
        .ZN(n97) );
  INV_X1 U187 ( .A(n98), .ZN(n214) );
  AOI22_X1 U188 ( .A1(instr_d[21]), .A2(n309), .B1(instr_q[21]), .B2(n308), 
        .ZN(n98) );
  INV_X1 U189 ( .A(n99), .ZN(n213) );
  AOI22_X1 U190 ( .A1(instr_d[20]), .A2(n309), .B1(instr_q[20]), .B2(n308), 
        .ZN(n99) );
  INV_X1 U191 ( .A(n100), .ZN(n194) );
  AOI22_X1 U192 ( .A1(instr_d[1]), .A2(n309), .B1(instr_q[1]), .B2(n308), .ZN(
        n100) );
  INV_X1 U193 ( .A(n101), .ZN(n212) );
  AOI22_X1 U194 ( .A1(instr_d[19]), .A2(n309), .B1(instr_q[19]), .B2(n308), 
        .ZN(n101) );
  INV_X1 U195 ( .A(n102), .ZN(n211) );
  AOI22_X1 U196 ( .A1(instr_d[18]), .A2(n309), .B1(instr_q[18]), .B2(n308), 
        .ZN(n102) );
  INV_X1 U197 ( .A(n103), .ZN(n210) );
  AOI22_X1 U198 ( .A1(instr_d[17]), .A2(n309), .B1(instr_q[17]), .B2(n308), 
        .ZN(n103) );
  INV_X1 U199 ( .A(n104), .ZN(n209) );
  AOI22_X1 U200 ( .A1(instr_d[16]), .A2(n309), .B1(instr_q[16]), .B2(n308), 
        .ZN(n104) );
  INV_X1 U201 ( .A(n105), .ZN(n208) );
  AOI22_X1 U202 ( .A1(instr_d[15]), .A2(n309), .B1(instr_q[15]), .B2(n308), 
        .ZN(n105) );
  INV_X1 U203 ( .A(n106), .ZN(n207) );
  AOI22_X1 U204 ( .A1(instr_d[14]), .A2(n309), .B1(instr_q[14]), .B2(n308), 
        .ZN(n106) );
  INV_X1 U205 ( .A(n107), .ZN(n206) );
  AOI22_X1 U206 ( .A1(instr_d[13]), .A2(n309), .B1(instr_q[13]), .B2(n308), 
        .ZN(n107) );
  INV_X1 U207 ( .A(n108), .ZN(n205) );
  AOI22_X1 U208 ( .A1(instr_d[12]), .A2(n309), .B1(instr_q[12]), .B2(n308), 
        .ZN(n108) );
  INV_X1 U209 ( .A(n109), .ZN(n204) );
  AOI22_X1 U210 ( .A1(instr_d[11]), .A2(n309), .B1(instr_q[11]), .B2(n308), 
        .ZN(n109) );
  INV_X1 U211 ( .A(n110), .ZN(n203) );
  AOI22_X1 U212 ( .A1(instr_d[10]), .A2(n309), .B1(instr_q[10]), .B2(n308), 
        .ZN(n110) );
  INV_X1 U213 ( .A(n111), .ZN(n193) );
  AOI221_X1 U214 ( .B1(instr_q[0]), .B2(n308), .C1(instr_d[0]), .C2(n309), .A(
        n85), .ZN(n111) );
  NOR2_X1 U215 ( .A1(n3), .A2(ctrl[0]), .ZN(n85) );
  INV_X1 U216 ( .A(n112), .ZN(n3) );
  OAI21_X1 U217 ( .B1(ctrl[1]), .B2(ctrl[0]), .A(n113), .ZN(n112) );
  INV_X1 U218 ( .A(n114), .ZN(n190) );
  AOI22_X1 U219 ( .A1(fp_q), .A2(n301), .B1(fp_d), .B2(n291), .ZN(n114) );
  INV_X1 U220 ( .A(n115), .ZN(n187) );
  AOI22_X1 U221 ( .A1(dSize_q[1]), .A2(n301), .B1(dSize_d[1]), .B2(n292), .ZN(
        n115) );
  INV_X1 U222 ( .A(n116), .ZN(n186) );
  AOI22_X1 U223 ( .A1(dSize_q[0]), .A2(n301), .B1(dSize_d[0]), .B2(n292), .ZN(
        n116) );
  INV_X1 U224 ( .A(n117), .ZN(n158) );
  AOI22_X1 U225 ( .A1(aluRes_q[9]), .A2(n301), .B1(aluRes_d[9]), .B2(n292), 
        .ZN(n117) );
  INV_X1 U226 ( .A(n118), .ZN(n157) );
  AOI22_X1 U227 ( .A1(aluRes_q[8]), .A2(n301), .B1(aluRes_d[8]), .B2(n292), 
        .ZN(n118) );
  INV_X1 U228 ( .A(n119), .ZN(n156) );
  AOI22_X1 U229 ( .A1(aluRes_q[7]), .A2(n301), .B1(aluRes_d[7]), .B2(n292), 
        .ZN(n119) );
  INV_X1 U230 ( .A(n120), .ZN(n155) );
  AOI22_X1 U231 ( .A1(aluRes_q[6]), .A2(n301), .B1(aluRes_d[6]), .B2(n292), 
        .ZN(n120) );
  INV_X1 U232 ( .A(n121), .ZN(n154) );
  AOI22_X1 U233 ( .A1(aluRes_q[5]), .A2(n301), .B1(aluRes_d[5]), .B2(n292), 
        .ZN(n121) );
  INV_X1 U234 ( .A(n122), .ZN(n153) );
  AOI22_X1 U235 ( .A1(aluRes_q[4]), .A2(n301), .B1(aluRes_d[4]), .B2(n292), 
        .ZN(n122) );
  INV_X1 U236 ( .A(n123), .ZN(n152) );
  AOI22_X1 U237 ( .A1(aluRes_q[3]), .A2(n301), .B1(aluRes_d[3]), .B2(n292), 
        .ZN(n123) );
  INV_X1 U238 ( .A(n124), .ZN(n180) );
  AOI22_X1 U239 ( .A1(aluRes_q[31]), .A2(n301), .B1(aluRes_d[31]), .B2(n292), 
        .ZN(n124) );
  INV_X1 U240 ( .A(n125), .ZN(n179) );
  AOI22_X1 U241 ( .A1(aluRes_q[30]), .A2(n301), .B1(aluRes_d[30]), .B2(n292), 
        .ZN(n125) );
  INV_X1 U242 ( .A(n126), .ZN(n151) );
  AOI22_X1 U243 ( .A1(aluRes_q[2]), .A2(n301), .B1(aluRes_d[2]), .B2(n292), 
        .ZN(n126) );
  INV_X1 U244 ( .A(n127), .ZN(n178) );
  AOI22_X1 U245 ( .A1(aluRes_q[29]), .A2(n301), .B1(aluRes_d[29]), .B2(n291), 
        .ZN(n127) );
  INV_X1 U246 ( .A(n128), .ZN(n177) );
  AOI22_X1 U247 ( .A1(aluRes_q[28]), .A2(n301), .B1(aluRes_d[28]), .B2(n291), 
        .ZN(n128) );
  INV_X1 U248 ( .A(n129), .ZN(n176) );
  AOI22_X1 U249 ( .A1(aluRes_q[27]), .A2(n301), .B1(aluRes_d[27]), .B2(n291), 
        .ZN(n129) );
  INV_X1 U250 ( .A(n130), .ZN(n175) );
  AOI22_X1 U251 ( .A1(aluRes_q[26]), .A2(n300), .B1(aluRes_d[26]), .B2(n291), 
        .ZN(n130) );
  INV_X1 U252 ( .A(n131), .ZN(n174) );
  AOI22_X1 U253 ( .A1(aluRes_q[25]), .A2(n300), .B1(aluRes_d[25]), .B2(n291), 
        .ZN(n131) );
  INV_X1 U254 ( .A(n132), .ZN(n173) );
  AOI22_X1 U255 ( .A1(aluRes_q[24]), .A2(n300), .B1(aluRes_d[24]), .B2(n291), 
        .ZN(n132) );
  INV_X1 U256 ( .A(n133), .ZN(n172) );
  AOI22_X1 U257 ( .A1(aluRes_q[23]), .A2(n300), .B1(aluRes_d[23]), .B2(n291), 
        .ZN(n133) );
  INV_X1 U258 ( .A(n134), .ZN(n171) );
  AOI22_X1 U259 ( .A1(aluRes_q[22]), .A2(n300), .B1(aluRes_d[22]), .B2(n291), 
        .ZN(n134) );
  INV_X1 U260 ( .A(n135), .ZN(n170) );
  AOI22_X1 U261 ( .A1(aluRes_q[21]), .A2(n300), .B1(aluRes_d[21]), .B2(n291), 
        .ZN(n135) );
  INV_X1 U262 ( .A(n136), .ZN(n169) );
  AOI22_X1 U263 ( .A1(aluRes_q[20]), .A2(n300), .B1(aluRes_d[20]), .B2(n291), 
        .ZN(n136) );
  INV_X1 U264 ( .A(n137), .ZN(n150) );
  AOI22_X1 U265 ( .A1(aluRes_q[1]), .A2(n300), .B1(aluRes_d[1]), .B2(n291), 
        .ZN(n137) );
  INV_X1 U266 ( .A(n138), .ZN(n168) );
  AOI22_X1 U267 ( .A1(aluRes_q[19]), .A2(n300), .B1(aluRes_d[19]), .B2(n290), 
        .ZN(n138) );
  INV_X1 U268 ( .A(n139), .ZN(n167) );
  AOI22_X1 U269 ( .A1(aluRes_q[18]), .A2(n300), .B1(aluRes_d[18]), .B2(n290), 
        .ZN(n139) );
  INV_X1 U270 ( .A(n140), .ZN(n166) );
  AOI22_X1 U271 ( .A1(aluRes_q[17]), .A2(n300), .B1(aluRes_d[17]), .B2(n290), 
        .ZN(n140) );
  INV_X1 U272 ( .A(n141), .ZN(n165) );
  AOI22_X1 U273 ( .A1(aluRes_q[16]), .A2(n300), .B1(aluRes_d[16]), .B2(n290), 
        .ZN(n141) );
  INV_X1 U274 ( .A(n142), .ZN(n164) );
  AOI22_X1 U275 ( .A1(aluRes_q[15]), .A2(n300), .B1(aluRes_d[15]), .B2(n290), 
        .ZN(n142) );
  INV_X1 U276 ( .A(n143), .ZN(n163) );
  AOI22_X1 U277 ( .A1(aluRes_q[14]), .A2(n300), .B1(aluRes_d[14]), .B2(n290), 
        .ZN(n143) );
  INV_X1 U278 ( .A(n144), .ZN(n162) );
  AOI22_X1 U279 ( .A1(aluRes_q[13]), .A2(n300), .B1(aluRes_d[13]), .B2(n290), 
        .ZN(n144) );
  INV_X1 U280 ( .A(n145), .ZN(n161) );
  AOI22_X1 U281 ( .A1(aluRes_q[12]), .A2(n300), .B1(aluRes_d[12]), .B2(n290), 
        .ZN(n145) );
  INV_X1 U282 ( .A(n146), .ZN(n160) );
  AOI22_X1 U283 ( .A1(aluRes_q[11]), .A2(n300), .B1(aluRes_d[11]), .B2(n290), 
        .ZN(n146) );
  INV_X1 U284 ( .A(n147), .ZN(n159) );
  AOI22_X1 U285 ( .A1(aluRes_q[10]), .A2(n300), .B1(aluRes_d[10]), .B2(n290), 
        .ZN(n147) );
  INV_X1 U286 ( .A(n148), .ZN(n149) );
  AOI22_X1 U287 ( .A1(aluRes_q[0]), .A2(n300), .B1(aluRes_d[0]), .B2(n290), 
        .ZN(n148) );
  NAND2_X1 U289 ( .A1(rst), .A2(n309), .ZN(n6) );
  NAND2_X1 U291 ( .A1(ctrl[1]), .A2(ctrl[0]), .ZN(n113) );
  INV_X4 U292 ( .A(n6), .ZN(n307) );
  INV_X4 U293 ( .A(n300), .ZN(n290) );
  INV_X4 U294 ( .A(n305), .ZN(n300) );
  INV_X4 U295 ( .A(n305), .ZN(n301) );
  INV_X4 U296 ( .A(n305), .ZN(n299) );
  INV_X4 U297 ( .A(n299), .ZN(n291) );
  INV_X4 U298 ( .A(n299), .ZN(n292) );
  INV_X4 U299 ( .A(n307), .ZN(n306) );
  INV_X4 U300 ( .A(n306), .ZN(n305) );
  INV_X4 U301 ( .A(n113), .ZN(n309) );
  INV_X4 U302 ( .A(n305), .ZN(n298) );
  INV_X4 U303 ( .A(n298), .ZN(n293) );
  INV_X4 U304 ( .A(n298), .ZN(n294) );
  INV_X4 U305 ( .A(n305), .ZN(n297) );
  INV_X4 U306 ( .A(n297), .ZN(n295) );
  INV_X4 U307 ( .A(n297), .ZN(n296) );
  INV_X4 U308 ( .A(n112), .ZN(n308) );
  INV_X4 U309 ( .A(n306), .ZN(n304) );
  INV_X4 U310 ( .A(n304), .ZN(n302) );
  INV_X4 U311 ( .A(n304), .ZN(n303) );
endmodule

