
module multiplier ( a, b, control, product_in, product_out );
  input [31:0] a;
  input [31:0] b;
  input [1:0] control;
  input [31:0] product_in;
  output [31:0] product_out;
  wire   net327996, net327997, net327998, net327999, net328000, net328003,
         net328013, net328016, net328019, net328020, net328021, net328023,
         net328024, net328025, net328026, net328028, net328029, net328030,
         net328031, net328035, net328039, net328046, net328051, net328068,
         net328083, net328105, net328110, net328113, net328117, net328118,
         net328120, net328122, net328123, net328125, net328128, net328142,
         net328147, net328158, net328160, net328162, net328168, net328172,
         net328177, net328179, net328180, net328183, net328192, net328222,
         net328229, net328231, net328232, net328233, net328234, net328235,
         net328244, net328245, net328247, net328250, net328253, net328254,
         net328259, net328260, net328264, net328268, net328272, net328274,
         net328309, net328331, net328338, net328385, net328388, net328389,
         net328392, net328393, net328403, net328404, net328406, net328408,
         net328409, net328414, net328415, net328450, net328470, net328483,
         net328484, net328485, net328491, net328527, net328528, net328533,
         net328555, net328562, net328563, net328564, net328568, net328573,
         net328574, net328575, net328582, net328585, net328588, net328595,
         net328596, net328597, net328599, net328601, net328602, net328603,
         net328604, net328605, net328606, net328607, net328615, net328616,
         net328712, net328734, net328736, net328737, net328738, net328741,
         net328748, net328750, net328751, net328752, net328790, net328791,
         net328851, net328853, net328855, net328856, net328860, net328861,
         net328864, net328865, net328866, net328869, net328871, net328872,
         net328911, net328912, net328916, net328936, net328937, net328980,
         net328981, net328982, net328983, net328984, net329000, net329006,
         net329014, net329015, net329017, net329018, net329019, net329033,
         net329043, net329052, net329055, net329112, net329193, net329194,
         net329225, net329230, net329289, net329295, net329297, net329340,
         net329343, net329344, net329345, net329352, net329395, net329397,
         net329398, net329399, net329404, net329407, net329410, net329441,
         net329445, net329451, net329453, net329454, net329456, net329457,
         net329459, net329464, net329465, net329467, net329472, net329545,
         net329547, net329549, net329552, net329556, net329559, net329560,
         net329592, net329593, net329598, net329690, net329737, net329743,
         net329750, net329751, net329753, net329754, net329755, net329802,
         net329803, net329808, net329810, net329812, net329813, net329824,
         net329857, net329858, net329859, net329860, net329866, net329868,
         net329873, net329876, net329918, net329965, net329970, net329972,
         net329973, net329974, net329986, net329988, net329990, net329992,
         net329994, net330021, net330024, net330025, net330028, net330029,
         net330033, net330037, net330038, net330039, net330040, net330042,
         net330043, net330044, net330067, net330088, net330089, net330098,
         net330110, net330126, net330127, net330130, net330131, net330134,
         net330142, net330173, net330197, net330204, net330213, net330234,
         net330238, net330239, net330327, net330330, net330331, net330334,
         net330336, net330337, net330338, net330377, net330379, net330382,
         net330383, net330384, net330406, net330456, net330457, net330458,
         net330459, net330509, net330510, net330512, net330513, net330595,
         net330596, net330598, net330600, net330601, net330612, net330649,
         net330650, net330651, net330652, net330653, net330654, net330705,
         net330730, net330737, net330738, net330741, net330742, net330751,
         net330752, net330786, net330808, net330819, net330822, net330834,
         net330839, net330843, net330850, net330853, net330854, net330855,
         net330858, net330860, net330861, net330862, net330863, net330876,
         net330910, net330911, net330912, net330913, net330915, net330916,
         net330917, net330918, net330942, net330965, net330983, net330986,
         net330987, net330990, net330991, net330998, net330999, net331000,
         net331025, net331028, net331029, net331032, net331037, net331055,
         net331069, net331070, net331073, net331083, net331084, net331086,
         net331090, net331091, net331092, net331096, net331097, net331098,
         net331113, net331115, net331119, net331123, net331124, net331125,
         net331126, net331129, net331130, net331131, net331132, net331137,
         net331138, net331143, net331144, net331145, net331154, net331169,
         net331176, net331177, net331178, net331180, net331181, net331182,
         net331189, net331192, net331193, net331194, net331195, net331196,
         net331198, net331199, net331200, net331201, net331202, net331204,
         net331211, net331213, net331221, net331226, net331227, net331228,
         net331234, net331235, net331237, net331238, net331243, net331244,
         net331245, net331247, net331251, net331261, net331262, net331271,
         net331277, net331287, net331299, net331295, net331293, net331311,
         net331307, net331305, net331323, net331329, net331343, net331341,
         net331353, net331351, net331349, net331359, net331357, net331363,
         net331362, net331480, net331479, net331478, net331477, net331476,
         net331506, net331520, net331583, net331614, net331799, net331798,
         net331896, net331895, net331939, net331938, net332007, net332006,
         net332018, net332050, net332088, net332214, net332292, net332287,
         net332364, net332463, net332462, net332586, net332585, net332584,
         net332690, net332747, net332761, net332836, net332856, net332855,
         net332891, net332947, net332946, net332977, net332988, net332987,
         net333045, net333044, net333079, net333078, net333222, net333237,
         net333280, net333277, net333276, net333275, net333311, net333315,
         net333336, net333424, net333501, net333500, net333532, net333531,
         net333530, net333569, net333577, net333615, net333614, net333621,
         net333659, net333678, net333677, net333770, net333795, net333802,
         net333816, net333862, net333869, net333879, net333915, net333918,
         net333944, net333991, net334005, net334039, net334044, net334167,
         net334211, net334240, net334239, net334298, net334308, net334385,
         net334433, net334437, net334464, net328137, net328922, net328873,
         net331072, net328919, net334227, net332666, net330128, net329471,
         net332895, net332894, net328921, net328918, net328584, net328567,
         net328475, net330335, net330332, net330237, net330026, net333874,
         net333853, net331127, net331066, net331064, net331063, net331061,
         net331264, net328472, net332558, net328617, net328614, net328612,
         net328487, net328236, net329821, net329818, net329466, net333618,
         net331058, net330955, net330954, net330746, net332668, net328111,
         net328109, net327991, net332028, net328525, net328167, net328149,
         net328027, net329985, net329815, net329811, net329452, net334334,
         net330925, net330856, net330748, net330614, net331170, net329409,
         net329334, net332583, net332378, net328182, net328181, net328151,
         net328148, net328134, net328132, net328131, net328130, net328129,
         net328127, net328126, net328047, net331272, net331212, net329339,
         net329073, net329020, net331273, net331254, net331017, net334415,
         net330859, net330745, net333894, net332821, net332819, net332231,
         net332230, net329978, net329971, net329968, net329967, net329966,
         net329819, net329817, net329816, net329470, net333890, net333519,
         net331034, net331033, net331030, net330599, net330247, net330246,
         net330245, net330244, net328854, net328583, net328579, net328578,
         net328576, net328524, net328230, net330386, net330385, net329989,
         net329980, net329872, net329455, net331263, net327992, net331283,
         net331282, net329919, net329558, net329557, net329469, net329463,
         net329462, net329461, net329338, net329337, net329336, net331499,
         net331128, net331068, net331062, net330994, net328917, net328794,
         net328593, net329069, net329068, net328920, net331613, net331253,
         net331059, net331031, net328249, net328006, net334441, net332820,
         net329981, net332266, net332265, net332264, net331863, net331862,
         net331861, net331860, net331270, net331269, net328608, net328570,
         net328569, net328474, net328473, net328405, net328176, net328174,
         net328173, net328171, net328170, net328169, net331284, net329291,
         net329072, net329071, net329070, net329021, net328742, net328740,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1153, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493;

  NAND2_X2 U1133 ( .A1(net329812), .A2(net329811), .ZN(net329808) );
  NAND2_X4 U1134 ( .A1(n4396), .A2(n1291), .ZN(n3348) );
  OAI21_X2 U1135 ( .B1(n3922), .B2(net331295), .A(n3496), .ZN(n3191) );
  NAND2_X2 U1137 ( .A1(net329470), .A2(net329465), .ZN(net329802) );
  NAND2_X4 U1138 ( .A1(n3099), .A2(n3100), .ZN(n3333) );
  INV_X4 U1139 ( .A(net330509), .ZN(n1104) );
  INV_X4 U1140 ( .A(net330509), .ZN(net330384) );
  INV_X4 U1142 ( .A(n4099), .ZN(n4101) );
  INV_X4 U1143 ( .A(net330204), .ZN(net333500) );
  INV_X4 U1144 ( .A(n4297), .ZN(n4096) );
  INV_X8 U1145 ( .A(n4298), .ZN(n1795) );
  INV_X8 U1146 ( .A(n3410), .ZN(n2024) );
  OAI21_X1 U1147 ( .B1(n3923), .B2(net331295), .A(n2409), .ZN(n1417) );
  XNOR2_X1 U1148 ( .A(n3189), .B(n3188), .ZN(n3174) );
  INV_X1 U1149 ( .A(n2842), .ZN(n1105) );
  NAND2_X4 U1150 ( .A1(n2924), .A2(n1146), .ZN(n2841) );
  AND2_X2 U1151 ( .A1(n1622), .A2(n1115), .ZN(n1106) );
  NAND2_X4 U1152 ( .A1(n1299), .A2(n2956), .ZN(n1622) );
  INV_X8 U1154 ( .A(n3587), .ZN(n3411) );
  AND2_X2 U1155 ( .A1(n2736), .A2(n2739), .ZN(n1107) );
  INV_X4 U1156 ( .A(n1107), .ZN(n3484) );
  NAND2_X4 U1157 ( .A1(n1234), .A2(n1235), .ZN(n1108) );
  NAND2_X4 U1159 ( .A1(n3347), .A2(n3110), .ZN(n1291) );
  NAND3_X1 U1160 ( .A1(net333853), .A2(net330652), .A3(net330654), .ZN(
        net330819) );
  NAND2_X2 U1161 ( .A1(n2874), .A2(n2924), .ZN(n2875) );
  INV_X4 U1162 ( .A(n2679), .ZN(n1109) );
  INV_X8 U1163 ( .A(n1109), .ZN(n1110) );
  OAI211_X2 U1166 ( .C1(n3204), .C2(n1659), .A(n3203), .B(n1191), .ZN(n1167)
         );
  NAND2_X4 U1167 ( .A1(net330752), .A2(n1631), .ZN(n2183) );
  INV_X2 U1168 ( .A(n1359), .ZN(n2904) );
  AOI21_X2 U1169 ( .B1(n4125), .B2(n4124), .A(n3936), .ZN(n3926) );
  INV_X2 U1170 ( .A(n3618), .ZN(n3621) );
  NAND2_X2 U1171 ( .A1(n1369), .A2(n4286), .ZN(n4331) );
  INV_X2 U1172 ( .A(n4286), .ZN(n4287) );
  NAND2_X1 U1173 ( .A1(n4028), .A2(n4027), .ZN(n1111) );
  BUF_X8 U1174 ( .A(net329018), .Z(n1433) );
  NOR2_X4 U1175 ( .A1(n2770), .A2(n2771), .ZN(n2772) );
  NAND2_X2 U1176 ( .A1(net331357), .A2(a[10]), .ZN(n2562) );
  INV_X8 U1178 ( .A(n1801), .ZN(n3415) );
  XNOR2_X2 U1179 ( .A(n4444), .B(n1287), .ZN(n1738) );
  INV_X8 U1180 ( .A(n3567), .ZN(n1287) );
  OAI21_X2 U1183 ( .B1(n3213), .B2(n1636), .A(n1115), .ZN(n3214) );
  NAND2_X1 U1184 ( .A1(n3287), .A2(n3286), .ZN(n1113) );
  NAND2_X1 U1185 ( .A1(n3747), .A2(n1404), .ZN(n3750) );
  INV_X8 U1186 ( .A(n3164), .ZN(n1114) );
  INV_X8 U1187 ( .A(n3409), .ZN(n3164) );
  NAND2_X2 U1188 ( .A1(n1602), .A2(net330089), .ZN(net329471) );
  INV_X1 U1189 ( .A(n3488), .ZN(n3312) );
  NAND3_X2 U1191 ( .A1(n1646), .A2(a[10]), .A3(n2037), .ZN(n1115) );
  INV_X4 U1192 ( .A(n3827), .ZN(n1139) );
  NOR2_X2 U1194 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  INV_X1 U1195 ( .A(net328236), .ZN(net328233) );
  NAND3_X4 U1197 ( .A1(n1399), .A2(net330088), .A3(n2914), .ZN(n2917) );
  NAND2_X2 U1198 ( .A1(net330044), .A2(n1601), .ZN(net330088) );
  INV_X4 U1199 ( .A(n4004), .ZN(n4005) );
  INV_X8 U1200 ( .A(n2664), .ZN(n2578) );
  NOR2_X4 U1201 ( .A1(n4254), .A2(n4253), .ZN(n1412) );
  CLKBUF_X2 U1202 ( .A(n2918), .Z(n1116) );
  INV_X2 U1203 ( .A(n3555), .ZN(n3559) );
  CLKBUF_X2 U1204 ( .A(net329073), .Z(n1117) );
  INV_X4 U1205 ( .A(n4284), .ZN(n4181) );
  AND2_X4 U1206 ( .A1(n3742), .A2(n3741), .ZN(n1644) );
  INV_X4 U1207 ( .A(n3932), .ZN(n2017) );
  INV_X2 U1208 ( .A(n4024), .ZN(n1118) );
  OAI21_X2 U1209 ( .B1(net328233), .B2(net328234), .A(net328235), .ZN(
        net328232) );
  INV_X4 U1210 ( .A(n2240), .ZN(n2264) );
  INV_X2 U1211 ( .A(n2910), .ZN(n2882) );
  NAND2_X1 U1212 ( .A1(n3102), .A2(n2910), .ZN(n3000) );
  NAND2_X2 U1213 ( .A1(n3270), .A2(n3269), .ZN(n3435) );
  INV_X4 U1214 ( .A(n4146), .ZN(n4150) );
  INV_X8 U1215 ( .A(n2892), .ZN(n2893) );
  NAND2_X2 U1216 ( .A1(n2892), .A2(n2983), .ZN(n2987) );
  INV_X4 U1217 ( .A(net328122), .ZN(net328180) );
  XNOR2_X2 U1219 ( .A(net329291), .B(n1433), .ZN(n1119) );
  INV_X4 U1220 ( .A(n2787), .ZN(n1667) );
  NAND2_X2 U1222 ( .A1(n3165), .A2(n3407), .ZN(n3167) );
  NAND3_X1 U1223 ( .A1(n3095), .A2(n3407), .A3(n3408), .ZN(n3096) );
  NAND3_X2 U1224 ( .A1(n3617), .A2(n3616), .A3(n3615), .ZN(n1120) );
  NAND2_X2 U1225 ( .A1(net329070), .A2(net328873), .ZN(n1500) );
  INV_X8 U1227 ( .A(net329345), .ZN(net329459) );
  NAND3_X2 U1228 ( .A1(n3671), .A2(n3670), .A3(n3669), .ZN(n3673) );
  INV_X4 U1229 ( .A(n3794), .ZN(n3792) );
  INV_X4 U1230 ( .A(n2938), .ZN(n3046) );
  XNOR2_X2 U1231 ( .A(n1139), .B(n3663), .ZN(n1121) );
  XNOR2_X1 U1232 ( .A(n1139), .B(n3663), .ZN(net328029) );
  NAND2_X2 U1233 ( .A1(net331226), .A2(net330991), .ZN(n2063) );
  NAND3_X1 U1234 ( .A1(n3211), .A2(n3092), .A3(n3007), .ZN(n1122) );
  NAND4_X4 U1235 ( .A1(n2077), .A2(n2076), .A3(net331253), .A4(a[3]), .ZN(
        n2078) );
  XNOR2_X2 U1237 ( .A(net328597), .B(n3907), .ZN(n1711) );
  XNOR2_X2 U1238 ( .A(n3907), .B(net328614), .ZN(n1123) );
  INV_X8 U1239 ( .A(net328597), .ZN(net328614) );
  OAI21_X4 U1240 ( .B1(net331311), .B2(net330173), .A(n2813), .ZN(n1124) );
  INV_X4 U1241 ( .A(n2814), .ZN(n2813) );
  NAND2_X4 U1243 ( .A1(n1900), .A2(n1901), .ZN(n2434) );
  NAND2_X2 U1244 ( .A1(n4447), .A2(n1900), .ZN(n1163) );
  INV_X2 U1246 ( .A(net334441), .ZN(n1126) );
  NAND2_X2 U1247 ( .A1(n1962), .A2(n1961), .ZN(n3811) );
  INV_X4 U1248 ( .A(n2786), .ZN(n2787) );
  NAND2_X1 U1249 ( .A1(n4429), .A2(n2110), .ZN(n2113) );
  NAND2_X2 U1250 ( .A1(n2084), .A2(n2083), .ZN(n2110) );
  XNOR2_X2 U1251 ( .A(net330954), .B(net331058), .ZN(n1127) );
  INV_X4 U1252 ( .A(n1127), .ZN(net331055) );
  NAND2_X4 U1254 ( .A1(n2791), .A2(n2848), .ZN(n2792) );
  OAI21_X4 U1255 ( .B1(n2577), .B2(n2576), .A(n2575), .ZN(n1625) );
  INV_X4 U1256 ( .A(n1407), .ZN(n1252) );
  NAND2_X4 U1257 ( .A1(n3030), .A2(n2848), .ZN(n1129) );
  NAND2_X2 U1258 ( .A1(n4066), .A2(n4065), .ZN(n1974) );
  NAND2_X2 U1259 ( .A1(n1414), .A2(n3712), .ZN(n3804) );
  INV_X2 U1260 ( .A(net333044), .ZN(net333045) );
  INV_X4 U1261 ( .A(n3011), .ZN(n2754) );
  NAND2_X4 U1262 ( .A1(n2590), .A2(n1153), .ZN(n1156) );
  INV_X2 U1263 ( .A(net328872), .ZN(n1130) );
  INV_X8 U1264 ( .A(n1130), .ZN(n1131) );
  NAND2_X2 U1265 ( .A1(net329454), .A2(net329593), .ZN(net329970) );
  INV_X4 U1266 ( .A(net329970), .ZN(n1556) );
  INV_X4 U1267 ( .A(net329021), .ZN(net333991) );
  NAND2_X4 U1268 ( .A1(n2484), .A2(n2485), .ZN(n1132) );
  NOR2_X2 U1269 ( .A1(n1403), .A2(n3554), .ZN(net334433) );
  INV_X4 U1270 ( .A(net334433), .ZN(net328856) );
  NAND2_X2 U1272 ( .A1(net328737), .A2(net328738), .ZN(net328736) );
  NAND2_X4 U1273 ( .A1(n4305), .A2(n4304), .ZN(n1134) );
  NAND2_X4 U1274 ( .A1(n4305), .A2(n4304), .ZN(n1135) );
  INV_X2 U1275 ( .A(n1427), .ZN(n1190) );
  OAI21_X2 U1276 ( .B1(n4423), .B2(n3318), .A(n3194), .ZN(n2999) );
  INV_X4 U1277 ( .A(n2999), .ZN(n3088) );
  INV_X8 U1278 ( .A(n3653), .ZN(n1267) );
  NOR2_X1 U1279 ( .A1(n3662), .A2(n3661), .ZN(n1155) );
  NOR2_X2 U1280 ( .A1(n1155), .A2(n3963), .ZN(n3964) );
  NAND2_X4 U1281 ( .A1(n3971), .A2(n3970), .ZN(n4017) );
  NOR4_X4 U1283 ( .A1(n4198), .A2(n1580), .A3(n1137), .A4(n4197), .ZN(n1136)
         );
  INV_X32 U1284 ( .A(n4206), .ZN(n1137) );
  INV_X8 U1285 ( .A(n4207), .ZN(n4198) );
  NAND2_X1 U1286 ( .A1(net328035), .A2(n4194), .ZN(n4208) );
  INV_X2 U1287 ( .A(n4208), .ZN(n4197) );
  AOI21_X2 U1288 ( .B1(n2978), .B2(n3093), .A(n3091), .ZN(n1698) );
  INV_X4 U1289 ( .A(n1698), .ZN(n2995) );
  NAND2_X4 U1290 ( .A1(n3378), .A2(net329397), .ZN(n1138) );
  INV_X8 U1291 ( .A(n3752), .ZN(n3827) );
  INV_X4 U1293 ( .A(n3071), .ZN(n1662) );
  OAI221_X2 U1294 ( .B1(n4430), .B2(net328712), .C1(n3922), .C2(net331363), 
        .A(n3921), .ZN(n1140) );
  INV_X8 U1295 ( .A(n2024), .ZN(n2025) );
  NAND2_X2 U1297 ( .A1(n3225), .A2(n3226), .ZN(n1141) );
  INV_X4 U1298 ( .A(n3411), .ZN(n1142) );
  NOR2_X1 U1299 ( .A1(n1125), .A2(n3841), .ZN(n3569) );
  NAND3_X2 U1300 ( .A1(net330654), .A2(net330652), .A3(net333853), .ZN(n1143)
         );
  INV_X4 U1301 ( .A(n1314), .ZN(n2559) );
  NAND2_X2 U1302 ( .A1(n2574), .A2(n2573), .ZN(n2163) );
  NAND4_X2 U1304 ( .A1(control[1]), .A2(b[1]), .A3(control[0]), .A4(a[2]), 
        .ZN(n1202) );
  INV_X4 U1305 ( .A(n3158), .ZN(n1894) );
  NAND3_X2 U1306 ( .A1(n4106), .A2(n4135), .A3(net331299), .ZN(n4114) );
  NAND2_X4 U1307 ( .A1(n4135), .A2(net332584), .ZN(n4193) );
  OAI211_X4 U1308 ( .C1(n4105), .C2(n1173), .A(n4104), .B(n4103), .ZN(n4135)
         );
  CLKBUF_X3 U1310 ( .A(n3627), .Z(n1144) );
  XNOR2_X2 U1311 ( .A(n2994), .B(n2997), .ZN(n2968) );
  NAND2_X2 U1312 ( .A1(n2778), .A2(n2779), .ZN(n1146) );
  NOR2_X4 U1313 ( .A1(n2108), .A2(n2109), .ZN(n1145) );
  NAND2_X4 U1314 ( .A1(n1847), .A2(n1848), .ZN(n2108) );
  INV_X1 U1315 ( .A(net330650), .ZN(net331000) );
  INV_X32 U1316 ( .A(control[0]), .ZN(n1326) );
  INV_X1 U1317 ( .A(n1128), .ZN(n1637) );
  INV_X2 U1318 ( .A(n2776), .ZN(n2779) );
  NAND2_X1 U1320 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  INV_X4 U1321 ( .A(n1739), .ZN(n3155) );
  NAND2_X2 U1322 ( .A1(n3226), .A2(n1739), .ZN(n3157) );
  INV_X8 U1323 ( .A(n1230), .ZN(n1939) );
  INV_X1 U1324 ( .A(net328385), .ZN(n1148) );
  INV_X2 U1325 ( .A(n1148), .ZN(n1149) );
  INV_X2 U1326 ( .A(n2449), .ZN(n2447) );
  INV_X4 U1327 ( .A(n4130), .ZN(n3934) );
  NOR3_X2 U1328 ( .A1(n4130), .A2(net328254), .A3(n4131), .ZN(n4133) );
  NAND2_X4 U1329 ( .A1(n3231), .A2(n1850), .ZN(n1150) );
  NAND2_X2 U1330 ( .A1(n3231), .A2(n1850), .ZN(n3420) );
  NAND2_X4 U1331 ( .A1(n1365), .A2(n3170), .ZN(n3320) );
  NAND2_X2 U1332 ( .A1(n2103), .A2(n2102), .ZN(n1151) );
  NAND2_X4 U1333 ( .A1(n2101), .A2(n2100), .ZN(n2102) );
  NAND2_X4 U1336 ( .A1(n2588), .A2(n2589), .ZN(n1153) );
  INV_X8 U1337 ( .A(n2587), .ZN(n2588) );
  INV_X2 U1338 ( .A(n3253), .ZN(n1160) );
  INV_X2 U1339 ( .A(n3103), .ZN(n3027) );
  INV_X8 U1340 ( .A(net331069), .ZN(n1521) );
  INV_X4 U1341 ( .A(n4093), .ZN(n3956) );
  NAND2_X4 U1345 ( .A1(n2889), .A2(n3023), .ZN(n2909) );
  INV_X4 U1346 ( .A(n3662), .ZN(n3720) );
  INV_X2 U1347 ( .A(n4225), .ZN(n3837) );
  INV_X4 U1348 ( .A(n3837), .ZN(n1404) );
  NAND2_X2 U1349 ( .A1(n2590), .A2(net330028), .ZN(net330033) );
  NAND2_X2 U1350 ( .A1(n2587), .A2(n2586), .ZN(n2590) );
  INV_X1 U1351 ( .A(net329441), .ZN(n1157) );
  OAI211_X4 U1352 ( .C1(n1160), .C2(n3141), .A(n3249), .B(n3248), .ZN(n3144)
         );
  NAND2_X1 U1353 ( .A1(n1281), .A2(n3765), .ZN(n1961) );
  AND2_X2 U1354 ( .A1(n3150), .A2(n1655), .ZN(n1158) );
  XNOR2_X2 U1355 ( .A(net328864), .B(net328865), .ZN(n1159) );
  INV_X4 U1356 ( .A(n4213), .ZN(n3187) );
  NAND2_X2 U1357 ( .A1(n4145), .A2(net328231), .ZN(n4189) );
  NAND4_X4 U1359 ( .A1(n2131), .A2(n2130), .A3(n1207), .A4(n2026), .ZN(n2133)
         );
  INV_X4 U1361 ( .A(n2290), .ZN(n2675) );
  INV_X4 U1363 ( .A(n1313), .ZN(n1161) );
  NAND2_X4 U1364 ( .A1(net331068), .A2(net330650), .ZN(net331062) );
  INV_X2 U1365 ( .A(net334005), .ZN(n1162) );
  INV_X8 U1366 ( .A(net330247), .ZN(net334005) );
  INV_X1 U1367 ( .A(net331090), .ZN(n1164) );
  NAND2_X2 U1368 ( .A1(n1588), .A2(n1587), .ZN(net331058) );
  XOR2_X2 U1369 ( .A(n4274), .B(n4276), .Z(n1165) );
  XNOR2_X2 U1372 ( .A(n4467), .B(n3288), .ZN(n1166) );
  OAI21_X2 U1374 ( .B1(n4297), .B2(n4298), .A(n4296), .ZN(n4299) );
  INV_X2 U1375 ( .A(n3317), .ZN(n1659) );
  NAND2_X2 U1376 ( .A1(n4119), .A2(n4118), .ZN(net328260) );
  INV_X2 U1377 ( .A(n4127), .ZN(n4128) );
  AOI21_X4 U1378 ( .B1(net329754), .B2(net329345), .A(net329755), .ZN(n3109)
         );
  OAI21_X1 U1379 ( .B1(n1364), .B2(net331363), .A(n4111), .ZN(n1168) );
  NAND2_X4 U1380 ( .A1(net331066), .A2(n1597), .ZN(net331064) );
  NAND2_X4 U1381 ( .A1(n2073), .A2(n2072), .ZN(n1169) );
  NAND4_X4 U1382 ( .A1(n1310), .A2(b[8]), .A3(control[1]), .A4(a[3]), .ZN(
        n1170) );
  NAND2_X1 U1383 ( .A1(net328574), .A2(net328575), .ZN(n3908) );
  INV_X2 U1384 ( .A(n3121), .ZN(n2929) );
  OAI21_X2 U1386 ( .B1(n3273), .B2(n3277), .A(net333678), .ZN(n3424) );
  NAND2_X2 U1388 ( .A1(net330911), .A2(net330614), .ZN(net330910) );
  NOR2_X2 U1389 ( .A1(net330384), .A2(net334415), .ZN(net330601) );
  NAND2_X2 U1390 ( .A1(n1322), .A2(n1323), .ZN(net329818) );
  NAND2_X2 U1391 ( .A1(n3130), .A2(n3129), .ZN(n3250) );
  INV_X1 U1392 ( .A(n2035), .ZN(n1172) );
  INV_X32 U1393 ( .A(n2036), .ZN(n2034) );
  NAND2_X2 U1394 ( .A1(n4219), .A2(n4220), .ZN(n4224) );
  NAND2_X4 U1395 ( .A1(n2592), .A2(n2655), .ZN(n1817) );
  NAND2_X4 U1396 ( .A1(n3028), .A2(net329876), .ZN(n3029) );
  INV_X2 U1398 ( .A(net333045), .ZN(n1173) );
  NAND3_X4 U1399 ( .A1(n4428), .A2(control[0]), .A3(b[16]), .ZN(n1174) );
  NAND2_X1 U1400 ( .A1(a[8]), .A2(n2206), .ZN(n2209) );
  INV_X4 U1401 ( .A(n2096), .ZN(n2026) );
  INV_X2 U1402 ( .A(net329974), .ZN(net329978) );
  INV_X4 U1403 ( .A(n2279), .ZN(n2161) );
  INV_X8 U1404 ( .A(n2278), .ZN(n2162) );
  NOR2_X4 U1405 ( .A1(n3964), .A2(n3965), .ZN(n3966) );
  INV_X2 U1406 ( .A(n3961), .ZN(n3965) );
  OAI21_X4 U1407 ( .B1(n4388), .B2(n2758), .A(n2545), .ZN(n2463) );
  CLKBUF_X3 U1408 ( .A(net332977), .Z(net334437) );
  NAND2_X4 U1409 ( .A1(n4416), .A2(n2599), .ZN(n3019) );
  INV_X8 U1411 ( .A(net328405), .ZN(net328474) );
  OAI21_X4 U1412 ( .B1(net329821), .B2(net333532), .A(net329592), .ZN(
        net329743) );
  INV_X4 U1413 ( .A(net329456), .ZN(net329821) );
  NAND2_X4 U1414 ( .A1(n2598), .A2(n2597), .ZN(n1933) );
  INV_X4 U1417 ( .A(net328524), .ZN(net328234) );
  NAND2_X1 U1418 ( .A1(net329824), .A2(net329990), .ZN(net329974) );
  NOR2_X2 U1419 ( .A1(n2677), .A2(n1721), .ZN(n2678) );
  INV_X8 U1422 ( .A(n2435), .ZN(n2362) );
  INV_X4 U1424 ( .A(n3067), .ZN(n1276) );
  NAND2_X4 U1425 ( .A1(n1367), .A2(n1271), .ZN(net328570) );
  BUF_X4 U1426 ( .A(n3680), .Z(n1759) );
  NAND2_X4 U1427 ( .A1(n1864), .A2(n1863), .ZN(n2553) );
  NAND2_X2 U1428 ( .A1(net327991), .A2(net327992), .ZN(n1479) );
  NAND2_X2 U1429 ( .A1(net328491), .A2(n4072), .ZN(n1231) );
  OAI21_X4 U1430 ( .B1(n3878), .B2(n3877), .A(n3876), .ZN(n1175) );
  NAND4_X4 U1431 ( .A1(net331193), .A2(b[9]), .A3(control[1]), .A4(a[2]), .ZN(
        n1176) );
  NAND2_X2 U1432 ( .A1(n4060), .A2(n4059), .ZN(n1179) );
  NAND2_X4 U1433 ( .A1(n1177), .A2(n1178), .ZN(n1180) );
  NAND2_X4 U1434 ( .A1(n1179), .A2(n1180), .ZN(n4062) );
  INV_X4 U1435 ( .A(n4060), .ZN(n1177) );
  INV_X4 U1436 ( .A(n4059), .ZN(n1178) );
  NAND2_X2 U1437 ( .A1(n1758), .A2(n1757), .ZN(n1183) );
  NAND2_X4 U1438 ( .A1(n1181), .A2(n1182), .ZN(n1184) );
  NAND2_X4 U1439 ( .A1(n1183), .A2(n1184), .ZN(net327997) );
  INV_X4 U1440 ( .A(n1757), .ZN(n1181) );
  INV_X4 U1441 ( .A(n1758), .ZN(n1182) );
  INV_X8 U1443 ( .A(n4062), .ZN(n4063) );
  NAND2_X4 U1444 ( .A1(n4061), .A2(n4062), .ZN(n4180) );
  NAND2_X2 U1445 ( .A1(net330839), .A2(a[5]), .ZN(n2279) );
  NAND2_X4 U1446 ( .A1(n2740), .A2(n2739), .ZN(n2979) );
  CLKBUF_X3 U1447 ( .A(n2399), .Z(n1676) );
  INV_X4 U1448 ( .A(n3387), .ZN(n1908) );
  INV_X4 U1450 ( .A(n3574), .ZN(n1725) );
  OAI21_X2 U1451 ( .B1(n3105), .B2(n3104), .A(n3333), .ZN(n3106) );
  NAND2_X2 U1452 ( .A1(n4093), .A2(n4090), .ZN(n4100) );
  INV_X4 U1453 ( .A(n3967), .ZN(n1665) );
  INV_X4 U1454 ( .A(n3419), .ZN(n1301) );
  NOR2_X2 U1456 ( .A1(n4014), .A2(n3947), .ZN(n3949) );
  NOR2_X4 U1457 ( .A1(n3947), .A2(n1280), .ZN(n1281) );
  INV_X8 U1458 ( .A(n1730), .ZN(n3480) );
  NAND2_X4 U1459 ( .A1(n1490), .A2(n1491), .ZN(n1730) );
  NAND2_X2 U1460 ( .A1(n4130), .A2(net328260), .ZN(n4033) );
  NOR2_X2 U1461 ( .A1(n3228), .A2(n1940), .ZN(n3232) );
  NAND2_X2 U1462 ( .A1(n3397), .A2(n1246), .ZN(n3399) );
  INV_X2 U1463 ( .A(n3397), .ZN(n3314) );
  BUF_X32 U1464 ( .A(n2521), .Z(n1185) );
  NAND2_X4 U1465 ( .A1(n1708), .A2(n3072), .ZN(n3074) );
  INV_X8 U1466 ( .A(n2901), .ZN(n2903) );
  NAND2_X4 U1467 ( .A1(n2606), .A2(n2605), .ZN(n1186) );
  INV_X8 U1468 ( .A(n2604), .ZN(n2605) );
  NAND2_X4 U1469 ( .A1(n2980), .A2(n2982), .ZN(n2824) );
  NAND2_X2 U1470 ( .A1(n3187), .A2(n4212), .ZN(n3501) );
  OAI21_X2 U1471 ( .B1(n2419), .B2(n2418), .A(n1983), .ZN(n1187) );
  INV_X4 U1472 ( .A(n2336), .ZN(n1188) );
  INV_X4 U1473 ( .A(n1188), .ZN(n1189) );
  XNOR2_X2 U1474 ( .A(n2610), .B(n2630), .ZN(n1706) );
  NAND2_X2 U1475 ( .A1(n2610), .A2(n2630), .ZN(n1241) );
  INV_X4 U1477 ( .A(n1190), .ZN(n1191) );
  NAND2_X4 U1478 ( .A1(n3187), .A2(n4212), .ZN(n1192) );
  NAND2_X2 U1480 ( .A1(n3081), .A2(n3490), .ZN(n3086) );
  NAND2_X2 U1481 ( .A1(n1192), .A2(n1355), .ZN(n3313) );
  XNOR2_X2 U1482 ( .A(n3835), .B(n1672), .ZN(product_out[25]) );
  INV_X2 U1483 ( .A(n2039), .ZN(n1203) );
  INV_X4 U1484 ( .A(n3245), .ZN(n1193) );
  INV_X4 U1486 ( .A(n3431), .ZN(n3245) );
  INV_X8 U1487 ( .A(n1537), .ZN(n1536) );
  NOR2_X4 U1488 ( .A1(n1560), .A2(n1559), .ZN(n1194) );
  NOR2_X2 U1489 ( .A1(n1560), .A2(n1559), .ZN(n1195) );
  INV_X8 U1490 ( .A(n1561), .ZN(n1560) );
  NAND3_X2 U1491 ( .A1(net331251), .A2(n1293), .A3(b[24]), .ZN(n1210) );
  INV_X8 U1492 ( .A(n2375), .ZN(n1702) );
  INV_X8 U1493 ( .A(net328249), .ZN(net331613) );
  AOI22_X4 U1494 ( .A1(b[27]), .A2(net331613), .B1(b[19]), .B2(net328035), 
        .ZN(n1512) );
  AOI22_X4 U1495 ( .A1(b[28]), .A2(net331613), .B1(b[20]), .B2(net328035), 
        .ZN(n1566) );
  CLKBUF_X2 U1496 ( .A(n2247), .Z(n1196) );
  NAND2_X4 U1497 ( .A1(n2631), .A2(n2632), .ZN(n2547) );
  INV_X16 U1498 ( .A(control[1]), .ZN(net332836) );
  INV_X4 U1499 ( .A(net331030), .ZN(net331034) );
  OAI21_X4 U1500 ( .B1(n1203), .B2(n2207), .A(n2105), .ZN(n2167) );
  NAND3_X4 U1501 ( .A1(net331193), .A2(control[1]), .A3(b[8]), .ZN(n1197) );
  NAND4_X4 U1502 ( .A1(net331284), .A2(net331283), .A3(n1204), .A4(n1324), 
        .ZN(net328105) );
  NOR2_X2 U1503 ( .A1(n2677), .A2(n1717), .ZN(n2165) );
  NAND2_X4 U1504 ( .A1(n3875), .A2(n3995), .ZN(n1198) );
  NAND2_X2 U1505 ( .A1(n3875), .A2(n3995), .ZN(n3996) );
  NAND2_X4 U1506 ( .A1(n3871), .A2(n3872), .ZN(n3875) );
  NAND4_X4 U1507 ( .A1(a[3]), .A2(b[16]), .A3(control[0]), .A4(net331200), 
        .ZN(n1199) );
  INV_X8 U1508 ( .A(n2056), .ZN(n2070) );
  NAND3_X4 U1509 ( .A1(net331192), .A2(control[0]), .A3(b[17]), .ZN(n1200) );
  OAI21_X4 U1511 ( .B1(n4029), .B2(net331295), .A(net328415), .ZN(n4036) );
  NAND2_X2 U1512 ( .A1(net331154), .A2(net331084), .ZN(n2061) );
  INV_X4 U1513 ( .A(net331145), .ZN(net331084) );
  NAND3_X4 U1515 ( .A1(n1293), .A2(b[9]), .A3(control[1]), .ZN(n1204) );
  INV_X4 U1516 ( .A(n2096), .ZN(n1205) );
  NAND2_X4 U1517 ( .A1(n2055), .A2(n2054), .ZN(n2056) );
  INV_X8 U1518 ( .A(n2862), .ZN(n2936) );
  INV_X2 U1519 ( .A(n3255), .ZN(n3141) );
  INV_X4 U1521 ( .A(n2226), .ZN(n1898) );
  INV_X2 U1522 ( .A(net329230), .ZN(net329289) );
  INV_X4 U1523 ( .A(n2179), .ZN(n1206) );
  NAND4_X4 U1525 ( .A1(a[2]), .A2(b[17]), .A3(control[0]), .A4(net331253), 
        .ZN(n1208) );
  NAND3_X4 U1526 ( .A1(net329919), .A2(n1311), .A3(b[24]), .ZN(n1209) );
  NAND2_X1 U1527 ( .A1(a[20]), .A2(net331323), .ZN(net328861) );
  INV_X8 U1528 ( .A(net328068), .ZN(net331311) );
  AND2_X4 U1529 ( .A1(a[14]), .A2(net331343), .ZN(n1211) );
  AND2_X2 U1530 ( .A1(a[14]), .A2(n2034), .ZN(n1212) );
  INV_X32 U1531 ( .A(control[0]), .ZN(net331254) );
  AND2_X4 U1532 ( .A1(a[22]), .A2(net331349), .ZN(n1213) );
  AND2_X4 U1533 ( .A1(a[24]), .A2(net331349), .ZN(n1214) );
  AND2_X4 U1534 ( .A1(a[28]), .A2(net331349), .ZN(n1215) );
  INV_X8 U1535 ( .A(n2081), .ZN(n2046) );
  AND2_X2 U1536 ( .A1(a[30]), .A2(n1719), .ZN(n1216) );
  NAND2_X4 U1537 ( .A1(n2568), .A2(n2567), .ZN(n2684) );
  NAND2_X2 U1538 ( .A1(n2441), .A2(n2440), .ZN(n2360) );
  AND2_X2 U1539 ( .A1(n2441), .A2(n2440), .ZN(n1217) );
  AND2_X4 U1540 ( .A1(n3645), .A2(n3696), .ZN(n1218) );
  INV_X4 U1541 ( .A(net330991), .ZN(net333874) );
  INV_X8 U1542 ( .A(net333874), .ZN(net333879) );
  INV_X8 U1543 ( .A(net329445), .ZN(net329441) );
  INV_X1 U1544 ( .A(net331798), .ZN(net331799) );
  INV_X4 U1545 ( .A(n2844), .ZN(n1283) );
  INV_X2 U1546 ( .A(net330327), .ZN(net332018) );
  INV_X8 U1547 ( .A(net329750), .ZN(n1277) );
  INV_X4 U1548 ( .A(n1392), .ZN(net328869) );
  NAND2_X4 U1549 ( .A1(n4393), .A2(n4006), .ZN(n3899) );
  NAND2_X4 U1550 ( .A1(n3804), .A2(n3803), .ZN(net328737) );
  INV_X8 U1551 ( .A(n2693), .ZN(n2003) );
  NAND2_X4 U1552 ( .A1(n1998), .A2(n1997), .ZN(n3016) );
  NAND2_X4 U1553 ( .A1(net328389), .A2(n1700), .ZN(n4076) );
  NAND2_X4 U1554 ( .A1(n3103), .A2(n3102), .ZN(n1940) );
  NAND2_X4 U1555 ( .A1(n3230), .A2(n3229), .ZN(n3332) );
  NAND2_X4 U1556 ( .A1(n2429), .A2(n2428), .ZN(n2430) );
  NAND2_X4 U1557 ( .A1(n3091), .A2(n3211), .ZN(n3409) );
  NAND2_X4 U1558 ( .A1(n4361), .A2(n4363), .ZN(n4303) );
  INV_X8 U1559 ( .A(net328854), .ZN(net328576) );
  NAND2_X4 U1560 ( .A1(n3201), .A2(n3200), .ZN(n1427) );
  OAI21_X4 U1561 ( .B1(n3206), .B2(n2976), .A(n2835), .ZN(n2891) );
  INV_X4 U1562 ( .A(n3726), .ZN(n3581) );
  XNOR2_X1 U1563 ( .A(n3395), .B(n1337), .ZN(n1219) );
  OAI221_X4 U1564 ( .B1(n4430), .B2(net328712), .C1(n3922), .C2(net331363), 
        .A(n3921), .ZN(n1647) );
  AND2_X2 U1565 ( .A1(n3310), .A2(n1246), .ZN(n1220) );
  INV_X2 U1566 ( .A(n3570), .ZN(n1360) );
  INV_X4 U1567 ( .A(n2192), .ZN(n2146) );
  NAND2_X2 U1568 ( .A1(n2926), .A2(n2925), .ZN(n2942) );
  INV_X2 U1569 ( .A(n2374), .ZN(n2292) );
  INV_X2 U1570 ( .A(n2445), .ZN(n2286) );
  CLKBUF_X2 U1572 ( .A(n2112), .Z(n1221) );
  NAND2_X2 U1573 ( .A1(n2219), .A2(n2573), .ZN(n2220) );
  NAND2_X1 U1575 ( .A1(n1222), .A2(n2390), .ZN(n1225) );
  NAND2_X2 U1576 ( .A1(n1224), .A2(n1225), .ZN(n1691) );
  INV_X2 U1577 ( .A(n2389), .ZN(n1222) );
  INV_X2 U1578 ( .A(n2390), .ZN(n1223) );
  NAND2_X2 U1579 ( .A1(n2388), .A2(n2019), .ZN(n1228) );
  NAND2_X4 U1580 ( .A1(n1226), .A2(n1227), .ZN(n1229) );
  NAND2_X4 U1581 ( .A1(n1228), .A2(n1229), .ZN(n2529) );
  INV_X4 U1582 ( .A(n2388), .ZN(n1226) );
  INV_X4 U1583 ( .A(n2019), .ZN(n1227) );
  NAND2_X4 U1584 ( .A1(n3044), .A2(n1661), .ZN(n1230) );
  NAND2_X2 U1585 ( .A1(n3552), .A2(n3551), .ZN(n1234) );
  NAND2_X4 U1586 ( .A1(n1232), .A2(n1233), .ZN(n1235) );
  NAND2_X4 U1587 ( .A1(n1234), .A2(n1235), .ZN(net329193) );
  INV_X4 U1588 ( .A(n3552), .ZN(n1232) );
  INV_X4 U1589 ( .A(n3551), .ZN(n1233) );
  INV_X4 U1590 ( .A(n3708), .ZN(n1236) );
  INV_X8 U1591 ( .A(n1236), .ZN(n1237) );
  NAND3_X1 U1592 ( .A1(a[19]), .A2(n3550), .A3(net331341), .ZN(n3708) );
  NAND2_X4 U1594 ( .A1(net330860), .A2(net330859), .ZN(net334044) );
  NAND2_X4 U1595 ( .A1(n1851), .A2(n1852), .ZN(net328406) );
  NOR2_X4 U1596 ( .A1(net334308), .A2(net331295), .ZN(n4295) );
  NAND2_X4 U1597 ( .A1(n3415), .A2(n3416), .ZN(n1329) );
  NAND4_X2 U1598 ( .A1(n1850), .A2(n3334), .A3(n1673), .A4(n3102), .ZN(n3219)
         );
  OAI21_X4 U1599 ( .B1(n1927), .B2(n1418), .A(n3583), .ZN(n3584) );
  XNOR2_X1 U1600 ( .A(n3472), .B(n1959), .ZN(n1692) );
  INV_X1 U1601 ( .A(n2738), .ZN(n1238) );
  NAND2_X4 U1602 ( .A1(n1239), .A2(n1240), .ZN(n1242) );
  NAND2_X4 U1603 ( .A1(n1242), .A2(n1241), .ZN(n2612) );
  INV_X4 U1604 ( .A(n2610), .ZN(n1239) );
  INV_X4 U1605 ( .A(n2630), .ZN(n1240) );
  INV_X2 U1606 ( .A(net328247), .ZN(n1243) );
  INV_X2 U1608 ( .A(net331263), .ZN(net331181) );
  OAI221_X4 U1609 ( .B1(n1925), .B2(n3589), .C1(n3588), .C2(n1142), .A(n3586), 
        .ZN(n3597) );
  NAND2_X4 U1610 ( .A1(n4058), .A2(n4156), .ZN(n4157) );
  INV_X4 U1611 ( .A(n4157), .ZN(n4059) );
  NOR2_X4 U1612 ( .A1(net328120), .A2(n1581), .ZN(net331938) );
  INV_X4 U1613 ( .A(n1400), .ZN(n4196) );
  NAND2_X2 U1614 ( .A1(net331154), .A2(n2129), .ZN(n2098) );
  INV_X4 U1615 ( .A(n3334), .ZN(n3228) );
  INV_X2 U1617 ( .A(n2770), .ZN(n1394) );
  INV_X4 U1618 ( .A(n4493), .ZN(n1244) );
  INV_X2 U1619 ( .A(n3293), .ZN(n1245) );
  INV_X4 U1620 ( .A(n3312), .ZN(n1246) );
  OAI21_X2 U1621 ( .B1(n2896), .B2(net331293), .A(net330067), .ZN(n1247) );
  NAND2_X2 U1622 ( .A1(n2811), .A2(n2812), .ZN(n1250) );
  NAND2_X4 U1623 ( .A1(n1248), .A2(n1249), .ZN(n1251) );
  NAND2_X4 U1624 ( .A1(n1250), .A2(n1251), .ZN(n2814) );
  INV_X4 U1625 ( .A(n2811), .ZN(n1248) );
  INV_X4 U1626 ( .A(n2812), .ZN(n1249) );
  INV_X4 U1627 ( .A(net329466), .ZN(net333677) );
  XNOR2_X2 U1628 ( .A(n2801), .B(n2802), .ZN(n1407) );
  INV_X4 U1629 ( .A(n2804), .ZN(n3013) );
  INV_X2 U1630 ( .A(n3881), .ZN(n3879) );
  AND2_X2 U1631 ( .A1(net329981), .A2(n1253), .ZN(n1254) );
  INV_X4 U1632 ( .A(net329815), .ZN(n1253) );
  NAND4_X2 U1633 ( .A1(n2867), .A2(n2868), .A3(a[13]), .A4(n2034), .ZN(n3038)
         );
  NAND2_X1 U1634 ( .A1(net330337), .A2(net330338), .ZN(n1598) );
  INV_X4 U1635 ( .A(n1538), .ZN(n1309) );
  NAND2_X4 U1636 ( .A1(n3993), .A2(n4152), .ZN(n4151) );
  NAND4_X4 U1637 ( .A1(a[25]), .A2(n3992), .A3(n4047), .A4(n2034), .ZN(n4152)
         );
  NAND2_X4 U1638 ( .A1(n3988), .A2(n3987), .ZN(n3992) );
  NAND2_X4 U1639 ( .A1(net328244), .A2(net331295), .ZN(net328122) );
  INV_X4 U1640 ( .A(n3770), .ZN(n3776) );
  NAND2_X2 U1641 ( .A1(n2642), .A2(n2641), .ZN(n1257) );
  NAND2_X2 U1642 ( .A1(n1255), .A2(n1256), .ZN(n1258) );
  NAND2_X2 U1643 ( .A1(n1257), .A2(n1258), .ZN(n2699) );
  INV_X4 U1644 ( .A(n2642), .ZN(n1255) );
  INV_X4 U1645 ( .A(n2641), .ZN(n1256) );
  INV_X4 U1646 ( .A(n2636), .ZN(n2701) );
  NAND2_X4 U1647 ( .A1(n2861), .A2(n1487), .ZN(n1784) );
  NAND2_X2 U1648 ( .A1(n1329), .A2(n3586), .ZN(n3419) );
  INV_X8 U1649 ( .A(n3402), .ZN(n1879) );
  NAND2_X2 U1650 ( .A1(n1113), .A2(n4455), .ZN(n3288) );
  NAND2_X2 U1651 ( .A1(n2353), .A2(n2354), .ZN(n2268) );
  INV_X1 U1652 ( .A(n2896), .ZN(n1716) );
  INV_X8 U1653 ( .A(n1909), .ZN(n1259) );
  NAND2_X2 U1654 ( .A1(n2060), .A2(n2059), .ZN(n1262) );
  NAND2_X4 U1655 ( .A1(n1260), .A2(n1261), .ZN(n1263) );
  NAND2_X4 U1656 ( .A1(n1263), .A2(n1262), .ZN(n2106) );
  INV_X8 U1657 ( .A(n2060), .ZN(n1260) );
  INV_X8 U1658 ( .A(n1169), .ZN(n1261) );
  NAND3_X4 U1659 ( .A1(net328918), .A2(net328584), .A3(net328920), .ZN(
        net328794) );
  INV_X4 U1660 ( .A(n1926), .ZN(net330038) );
  NAND2_X4 U1661 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
  INV_X2 U1662 ( .A(n4387), .ZN(n1683) );
  INV_X4 U1663 ( .A(net331273), .ZN(net331861) );
  NAND2_X1 U1664 ( .A1(n3151), .A2(n1264), .ZN(n1265) );
  NAND2_X2 U1665 ( .A1(n1158), .A2(n1447), .ZN(n1266) );
  NAND2_X2 U1666 ( .A1(n1265), .A2(n1266), .ZN(n1728) );
  INV_X1 U1667 ( .A(n1447), .ZN(n1264) );
  NAND2_X2 U1668 ( .A1(n3653), .A2(n1268), .ZN(n1269) );
  NAND2_X2 U1669 ( .A1(n1267), .A2(n3705), .ZN(n1270) );
  NAND2_X2 U1670 ( .A1(n1269), .A2(n1270), .ZN(n3654) );
  INV_X2 U1671 ( .A(n3705), .ZN(n1268) );
  BUF_X4 U1672 ( .A(n3355), .Z(n1447) );
  NOR2_X1 U1673 ( .A1(n1628), .A2(n3954), .ZN(n3957) );
  NOR2_X2 U1674 ( .A1(n3805), .A2(n3855), .ZN(n3806) );
  INV_X4 U1675 ( .A(n3808), .ZN(n3805) );
  NAND2_X4 U1676 ( .A1(net330839), .A2(a[0]), .ZN(net331143) );
  INV_X8 U1677 ( .A(n3506), .ZN(n1906) );
  NAND2_X4 U1678 ( .A1(n1199), .A2(net331244), .ZN(n2053) );
  NAND2_X4 U1679 ( .A1(n1430), .A2(n1431), .ZN(n3469) );
  INV_X4 U1680 ( .A(net328234), .ZN(n1271) );
  NAND2_X2 U1681 ( .A1(n3897), .A2(n3898), .ZN(n1274) );
  NAND2_X4 U1682 ( .A1(n1272), .A2(n1273), .ZN(n1275) );
  NAND2_X4 U1683 ( .A1(n1274), .A2(n1275), .ZN(net328574) );
  INV_X4 U1684 ( .A(n3897), .ZN(n1272) );
  INV_X4 U1685 ( .A(n3898), .ZN(n1273) );
  INV_X4 U1686 ( .A(n2627), .ZN(n2830) );
  NAND2_X2 U1687 ( .A1(n4466), .A2(n3067), .ZN(n1278) );
  NAND2_X4 U1688 ( .A1(n1276), .A2(n1277), .ZN(n1279) );
  NAND2_X4 U1689 ( .A1(n1278), .A2(n1279), .ZN(n3098) );
  INV_X4 U1691 ( .A(n4020), .ZN(n3293) );
  INV_X4 U1692 ( .A(n3948), .ZN(n1280) );
  INV_X4 U1693 ( .A(net329455), .ZN(net332050) );
  NAND2_X4 U1695 ( .A1(n2196), .A2(n2197), .ZN(n2255) );
  NAND2_X4 U1696 ( .A1(n2256), .A2(n2255), .ZN(n2321) );
  NAND2_X4 U1699 ( .A1(n1438), .A2(n1439), .ZN(n1441) );
  INV_X8 U1700 ( .A(n2053), .ZN(n2071) );
  NAND2_X4 U1701 ( .A1(n1541), .A2(net330382), .ZN(n1539) );
  INV_X2 U1702 ( .A(net328583), .ZN(n1282) );
  NAND2_X1 U1703 ( .A1(n2844), .A2(n2842), .ZN(n1284) );
  NAND2_X2 U1704 ( .A1(n1283), .A2(n1105), .ZN(n1285) );
  NAND2_X2 U1705 ( .A1(n1285), .A2(n1284), .ZN(n2791) );
  INV_X4 U1707 ( .A(net332231), .ZN(n1315) );
  NAND2_X4 U1708 ( .A1(n1594), .A2(n1330), .ZN(net329466) );
  NAND2_X4 U1709 ( .A1(n2397), .A2(n2398), .ZN(n2509) );
  NAND2_X4 U1710 ( .A1(n2508), .A2(n2509), .ZN(n2406) );
  NAND2_X2 U1711 ( .A1(n3467), .A2(n3527), .ZN(n1430) );
  NAND2_X2 U1712 ( .A1(net329810), .A2(net329471), .ZN(net330040) );
  INV_X4 U1713 ( .A(net329471), .ZN(net329469) );
  INV_X4 U1714 ( .A(n3978), .ZN(n3973) );
  OAI21_X2 U1715 ( .B1(n4285), .B2(n4284), .A(n4283), .ZN(n4286) );
  INV_X4 U1716 ( .A(n3585), .ZN(n3588) );
  INV_X8 U1717 ( .A(n2741), .ZN(n1286) );
  INV_X8 U1718 ( .A(n2962), .ZN(n2741) );
  NAND2_X4 U1719 ( .A1(n3679), .A2(n4421), .ZN(n3682) );
  NOR2_X2 U1720 ( .A1(net328180), .A2(net328181), .ZN(net328127) );
  NAND2_X2 U1721 ( .A1(n1970), .A2(n3567), .ZN(n1289) );
  NAND2_X4 U1722 ( .A1(n1287), .A2(n4444), .ZN(n1290) );
  NAND2_X4 U1723 ( .A1(n1289), .A2(n1290), .ZN(net328245) );
  INV_X2 U1725 ( .A(n1328), .ZN(n3893) );
  OAI21_X4 U1726 ( .B1(n4026), .B2(net331363), .A(n4025), .ZN(n4027) );
  NAND2_X2 U1727 ( .A1(net328260), .A2(n1111), .ZN(net328415) );
  INV_X4 U1729 ( .A(n2519), .ZN(n2520) );
  INV_X4 U1730 ( .A(n4300), .ZN(n4373) );
  NAND2_X2 U1731 ( .A1(n1390), .A2(n3154), .ZN(n1440) );
  NAND2_X4 U1732 ( .A1(n3584), .A2(n3963), .ZN(n3663) );
  OAI21_X4 U1733 ( .B1(n2825), .B2(n2824), .A(n1687), .ZN(n2895) );
  XOR2_X2 U1734 ( .A(n4289), .B(net328192), .Z(n1292) );
  XOR2_X1 U1735 ( .A(n4343), .B(n1292), .Z(n4290) );
  INV_X32 U1736 ( .A(control[0]), .ZN(n1293) );
  INV_X32 U1737 ( .A(control[0]), .ZN(n1294) );
  NAND2_X4 U1738 ( .A1(n3684), .A2(n1688), .ZN(n3428) );
  NOR2_X2 U1739 ( .A1(net328234), .A2(net328404), .ZN(net328568) );
  INV_X2 U1741 ( .A(n3711), .ZN(n1295) );
  INV_X4 U1742 ( .A(n1295), .ZN(n1296) );
  NOR2_X4 U1743 ( .A1(net329743), .A2(n3111), .ZN(n3115) );
  INV_X4 U1745 ( .A(n4255), .ZN(n4081) );
  NAND2_X2 U1749 ( .A1(n1804), .A2(n1805), .ZN(n3955) );
  NAND3_X2 U1750 ( .A1(n4087), .A2(n4086), .A3(n4085), .ZN(n3857) );
  INV_X8 U1751 ( .A(n3469), .ZN(n3522) );
  NAND2_X4 U1752 ( .A1(n3149), .A2(n3236), .ZN(n3153) );
  NAND2_X2 U1753 ( .A1(net328259), .A2(net328268), .ZN(n1945) );
  INV_X2 U1754 ( .A(n2855), .ZN(n2673) );
  INV_X2 U1755 ( .A(n4047), .ZN(n3991) );
  NOR2_X4 U1756 ( .A1(n3974), .A2(n3886), .ZN(n3890) );
  NAND2_X4 U1757 ( .A1(n3892), .A2(n3893), .ZN(n3900) );
  INV_X4 U1758 ( .A(n3154), .ZN(n1438) );
  NAND2_X2 U1759 ( .A1(n3299), .A2(n1167), .ZN(n3304) );
  NAND2_X4 U1760 ( .A1(n1896), .A2(n1897), .ZN(n1297) );
  NAND2_X2 U1761 ( .A1(n1896), .A2(n1897), .ZN(n3216) );
  INV_X1 U1762 ( .A(net328260), .ZN(n1583) );
  INV_X2 U1763 ( .A(n2416), .ZN(n2418) );
  INV_X4 U1764 ( .A(n3534), .ZN(n1298) );
  INV_X2 U1765 ( .A(n3534), .ZN(n3629) );
  NAND2_X2 U1766 ( .A1(n1504), .A2(net328236), .ZN(net328569) );
  OAI21_X4 U1767 ( .B1(n1252), .B2(n3014), .A(n3012), .ZN(n3018) );
  INV_X8 U1768 ( .A(n3212), .ZN(n3091) );
  NAND2_X4 U1769 ( .A1(n1300), .A2(n1301), .ZN(n1302) );
  NAND2_X4 U1770 ( .A1(n3418), .A2(n1302), .ZN(n3477) );
  INV_X2 U1771 ( .A(n3508), .ZN(n1300) );
  INV_X2 U1772 ( .A(n3992), .ZN(n3990) );
  INV_X1 U1773 ( .A(n3863), .ZN(n3788) );
  AOI21_X2 U1774 ( .B1(net328487), .B2(n1507), .A(net328567), .ZN(n1505) );
  INV_X2 U1775 ( .A(net328487), .ZN(net328483) );
  OR2_X4 U1776 ( .A1(n1313), .A2(a[6]), .ZN(n1354) );
  NAND2_X4 U1777 ( .A1(n2318), .A2(n2319), .ZN(n1303) );
  INV_X8 U1778 ( .A(n2317), .ZN(n2318) );
  NAND2_X2 U1780 ( .A1(n4139), .A2(n4082), .ZN(n3914) );
  NAND2_X2 U1781 ( .A1(net331798), .A2(n1456), .ZN(n1458) );
  NAND2_X4 U1782 ( .A1(n2535), .A2(n2534), .ZN(n2602) );
  INV_X1 U1783 ( .A(net334308), .ZN(net328179) );
  INV_X8 U1784 ( .A(n4480), .ZN(n2571) );
  OAI21_X1 U1785 ( .B1(n2701), .B2(n2700), .A(n2837), .ZN(n3009) );
  INV_X8 U1786 ( .A(net329454), .ZN(net329873) );
  NAND2_X4 U1787 ( .A1(n2241), .A2(n2421), .ZN(n2249) );
  NAND2_X4 U1788 ( .A1(net329069), .A2(net329068), .ZN(net328920) );
  XNOR2_X2 U1789 ( .A(net329559), .B(net329560), .ZN(net329339) );
  NAND2_X4 U1790 ( .A1(n4280), .A2(n4279), .ZN(n4316) );
  OAI21_X2 U1791 ( .B1(net329858), .B2(net329859), .A(net329598), .ZN(
        net329857) );
  NAND2_X4 U1792 ( .A1(n2710), .A2(n2711), .ZN(n2712) );
  NAND2_X1 U1793 ( .A1(n2545), .A2(n2544), .ZN(n1428) );
  AND2_X4 U1794 ( .A1(n2441), .A2(n2440), .ZN(n1415) );
  NAND2_X4 U1795 ( .A1(net330839), .A2(a[2]), .ZN(net331145) );
  INV_X1 U1796 ( .A(n4152), .ZN(n4153) );
  INV_X8 U1797 ( .A(n3122), .ZN(n3135) );
  NAND3_X2 U1798 ( .A1(n2755), .A2(net333944), .A3(n4458), .ZN(n2697) );
  INV_X2 U1799 ( .A(n4147), .ZN(n4268) );
  INV_X8 U1800 ( .A(n3509), .ZN(n1909) );
  NAND2_X1 U1801 ( .A1(net329441), .A2(net329690), .ZN(n1305) );
  NAND2_X4 U1802 ( .A1(n1304), .A2(n1157), .ZN(n1306) );
  NAND2_X4 U1803 ( .A1(n1305), .A2(n1306), .ZN(net329556) );
  INV_X4 U1804 ( .A(net329690), .ZN(n1304) );
  NAND2_X4 U1805 ( .A1(n2401), .A2(n2402), .ZN(n2403) );
  INV_X1 U1806 ( .A(n2563), .ZN(n2569) );
  NOR2_X4 U1807 ( .A1(n1159), .A2(net328861), .ZN(n1307) );
  INV_X4 U1808 ( .A(n1307), .ZN(net328588) );
  XNOR2_X2 U1809 ( .A(net330331), .B(n1309), .ZN(n1308) );
  INV_X32 U1810 ( .A(control[0]), .ZN(n1310) );
  INV_X32 U1811 ( .A(control[0]), .ZN(n1311) );
  INV_X32 U1812 ( .A(control[0]), .ZN(n1312) );
  INV_X2 U1813 ( .A(n2574), .ZN(n2576) );
  NAND2_X4 U1814 ( .A1(n2433), .A2(n2531), .ZN(n2496) );
  INV_X4 U1816 ( .A(net330843), .ZN(net332690) );
  NAND2_X4 U1818 ( .A1(n3003), .A2(n3002), .ZN(n3007) );
  INV_X8 U1819 ( .A(n2676), .ZN(n2575) );
  NAND2_X4 U1820 ( .A1(n3274), .A2(n3423), .ZN(n3383) );
  INV_X4 U1821 ( .A(n2878), .ZN(n1996) );
  NOR2_X2 U1822 ( .A1(net330600), .A2(net330599), .ZN(n1551) );
  NAND3_X4 U1823 ( .A1(n2785), .A2(net333501), .A3(net333869), .ZN(n1314) );
  INV_X8 U1824 ( .A(net332230), .ZN(net332231) );
  NAND2_X2 U1826 ( .A1(net332836), .A2(n1325), .ZN(net328249) );
  AND2_X2 U1827 ( .A1(net330043), .A2(net330042), .ZN(n1607) );
  NAND2_X4 U1828 ( .A1(control[0]), .A2(net331195), .ZN(n2077) );
  INV_X2 U1829 ( .A(n4448), .ZN(net329755) );
  INV_X2 U1830 ( .A(n4270), .ZN(n1988) );
  NOR2_X2 U1832 ( .A1(net328389), .A2(n1988), .ZN(n4074) );
  AOI21_X2 U1833 ( .B1(n1822), .B2(n4269), .A(n4268), .ZN(n4272) );
  INV_X8 U1834 ( .A(net330742), .ZN(net330247) );
  NOR2_X4 U1835 ( .A1(n1294), .A2(b[1]), .ZN(net331202) );
  NAND2_X4 U1836 ( .A1(net333659), .A2(net329992), .ZN(net329872) );
  NAND2_X2 U1837 ( .A1(a[8]), .A2(n2207), .ZN(n2208) );
  NAND2_X4 U1838 ( .A1(n3067), .A2(n3100), .ZN(n3066) );
  NAND2_X4 U1839 ( .A1(n2104), .A2(a[1]), .ZN(net331144) );
  INV_X8 U1840 ( .A(net331144), .ZN(net331204) );
  NAND2_X1 U1841 ( .A1(n4316), .A2(n4315), .ZN(n4317) );
  INV_X8 U1842 ( .A(n3363), .ZN(n3455) );
  NAND2_X2 U1843 ( .A1(n3595), .A2(n1329), .ZN(n3596) );
  NAND2_X2 U1844 ( .A1(net328172), .A2(net328171), .ZN(net331480) );
  NOR2_X2 U1845 ( .A1(n1319), .A2(n1568), .ZN(n1318) );
  OAI22_X1 U1846 ( .A1(net328712), .A2(n4108), .B1(n1733), .B2(net331363), 
        .ZN(n3500) );
  OAI22_X1 U1847 ( .A1(net328712), .A2(net328250), .B1(n1243), .B2(net331363), 
        .ZN(n3572) );
  OAI22_X1 U1848 ( .A1(n3816), .A2(net328712), .B1(n1133), .B2(net331363), 
        .ZN(n3182) );
  OAI22_X1 U1849 ( .A1(net328712), .A2(n3173), .B1(n3923), .B2(net331363), 
        .ZN(n3189) );
  NAND2_X2 U1850 ( .A1(n3476), .A2(n3477), .ZN(n1490) );
  NAND2_X2 U1851 ( .A1(n2693), .A2(net330327), .ZN(n2004) );
  INV_X4 U1852 ( .A(net331272), .ZN(net331860) );
  INV_X8 U1853 ( .A(n2057), .ZN(n2073) );
  INV_X8 U1854 ( .A(n4138), .ZN(n4259) );
  INV_X8 U1855 ( .A(n3298), .ZN(n4018) );
  NAND2_X2 U1856 ( .A1(n3622), .A2(n3435), .ZN(n3377) );
  NAND2_X4 U1857 ( .A1(n4291), .A2(n1685), .ZN(n4294) );
  NAND2_X1 U1859 ( .A1(n2693), .A2(net332018), .ZN(n1316) );
  NAND2_X2 U1860 ( .A1(n2003), .A2(net330327), .ZN(n1317) );
  INV_X4 U1862 ( .A(n3598), .ZN(n3764) );
  XNOR2_X2 U1863 ( .A(net328916), .B(net328751), .ZN(n1600) );
  INV_X4 U1864 ( .A(n3392), .ZN(n1443) );
  INV_X4 U1865 ( .A(net328137), .ZN(net328244) );
  NAND3_X1 U1866 ( .A1(n3220), .A2(n3218), .A3(n3219), .ZN(n3221) );
  INV_X8 U1867 ( .A(n2731), .ZN(n2738) );
  NAND2_X2 U1868 ( .A1(n3392), .A2(n3404), .ZN(n1445) );
  XNOR2_X2 U1871 ( .A(n4333), .B(n4332), .ZN(n1368) );
  AOI21_X2 U1872 ( .B1(n1615), .B2(n2855), .A(n2857), .ZN(n2770) );
  OAI211_X4 U1873 ( .C1(net329754), .C2(net333577), .A(net329803), .B(
        net329802), .ZN(n3067) );
  OR2_X2 U1874 ( .A1(n2376), .A2(n2377), .ZN(n1319) );
  NAND2_X2 U1875 ( .A1(net329819), .A2(n1555), .ZN(n1322) );
  NAND2_X4 U1876 ( .A1(n1320), .A2(n1321), .ZN(n1323) );
  INV_X1 U1877 ( .A(net329819), .ZN(n1320) );
  INV_X4 U1878 ( .A(n1555), .ZN(n1321) );
  NAND3_X4 U1879 ( .A1(n2454), .A2(n2456), .A3(n2455), .ZN(n2780) );
  NOR2_X1 U1880 ( .A1(n2105), .A2(n1345), .ZN(n2107) );
  NAND2_X4 U1881 ( .A1(net333615), .A2(net330730), .ZN(n2227) );
  NAND3_X4 U1882 ( .A1(control[0]), .A2(control[1]), .A3(b[1]), .ZN(n1324) );
  NAND2_X4 U1883 ( .A1(net329020), .A2(n1117), .ZN(net329291) );
  XNOR2_X2 U1884 ( .A(n3377), .B(n3430), .ZN(n1373) );
  NAND2_X4 U1885 ( .A1(n1957), .A2(n3766), .ZN(n4084) );
  NAND2_X2 U1886 ( .A1(net328588), .A2(net328582), .ZN(n3808) );
  NAND3_X4 U1887 ( .A1(n2210), .A2(net331357), .A3(a[7]), .ZN(n2280) );
  NAND2_X4 U1888 ( .A1(n2209), .A2(n2208), .ZN(n2210) );
  INV_X4 U1889 ( .A(net330134), .ZN(net330234) );
  NAND2_X4 U1890 ( .A1(n4468), .A2(n1536), .ZN(net330134) );
  INV_X4 U1891 ( .A(net329193), .ZN(n1503) );
  INV_X16 U1892 ( .A(control[0]), .ZN(n1325) );
  NAND3_X4 U1893 ( .A1(control[0]), .A2(control[1]), .A3(b[0]), .ZN(n1327) );
  NAND2_X4 U1894 ( .A1(n1197), .A2(n2045), .ZN(n2081) );
  AND2_X4 U1895 ( .A1(net332558), .A2(net328027), .ZN(net334308) );
  INV_X8 U1896 ( .A(n3379), .ZN(n3378) );
  NAND2_X4 U1897 ( .A1(net329467), .A2(n1399), .ZN(n2878) );
  NAND2_X4 U1898 ( .A1(net328236), .A2(net328524), .ZN(net331476) );
  NOR2_X1 U1899 ( .A1(n1704), .A2(n2564), .ZN(n2444) );
  NAND2_X2 U1900 ( .A1(n3969), .A2(n4099), .ZN(n3970) );
  INV_X4 U1901 ( .A(net331092), .ZN(net331090) );
  XNOR2_X2 U1903 ( .A(n3979), .B(n3891), .ZN(n1328) );
  NOR2_X4 U1904 ( .A1(net328583), .A2(net328919), .ZN(n1545) );
  INV_X8 U1905 ( .A(n3730), .ZN(n1927) );
  INV_X4 U1906 ( .A(n1760), .ZN(n1761) );
  NAND2_X4 U1907 ( .A1(n3504), .A2(n1879), .ZN(n3392) );
  INV_X4 U1908 ( .A(n3101), .ZN(n3026) );
  NAND2_X2 U1909 ( .A1(n2967), .A2(n2881), .ZN(n1636) );
  NAND2_X4 U1910 ( .A1(n3520), .A2(n3686), .ZN(n3612) );
  OAI21_X2 U1911 ( .B1(net328403), .B2(net328404), .A(net332891), .ZN(n4137)
         );
  NAND2_X4 U1912 ( .A1(n2040), .A2(n2046), .ZN(n2033) );
  NAND2_X2 U1913 ( .A1(n2039), .A2(n2040), .ZN(net330110) );
  NAND2_X4 U1914 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  AOI211_X4 U1915 ( .C1(n2360), .C2(n1778), .A(n2651), .B(n2656), .ZN(n2475)
         );
  INV_X8 U1916 ( .A(n3382), .ZN(n3421) );
  INV_X4 U1917 ( .A(n2125), .ZN(n2126) );
  INV_X8 U1918 ( .A(n2058), .ZN(n2072) );
  NAND2_X4 U1919 ( .A1(n3578), .A2(n1907), .ZN(n3404) );
  INV_X8 U1921 ( .A(n1297), .ZN(n3159) );
  INV_X4 U1922 ( .A(net330213), .ZN(net330098) );
  NAND2_X4 U1923 ( .A1(n3558), .A2(n3471), .ZN(n3562) );
  NAND2_X2 U1925 ( .A1(n3657), .A2(n3656), .ZN(n3756) );
  NAND2_X4 U1926 ( .A1(n3849), .A2(n4457), .ZN(n1786) );
  NAND2_X4 U1927 ( .A1(n2877), .A2(n2876), .ZN(net329593) );
  OAI21_X4 U1928 ( .B1(net328576), .B2(n4403), .A(net328853), .ZN(net328851)
         );
  NAND2_X4 U1929 ( .A1(n3159), .A2(n3160), .ZN(n3414) );
  NOR2_X2 U1930 ( .A1(net331614), .A2(n4022), .ZN(n4023) );
  NAND2_X2 U1931 ( .A1(n2941), .A2(n3044), .ZN(n3045) );
  NAND2_X2 U1932 ( .A1(n1457), .A2(n1458), .ZN(net329812) );
  NAND2_X2 U1933 ( .A1(n2747), .A2(n1980), .ZN(n1981) );
  NOR2_X2 U1934 ( .A1(n2269), .A2(n2270), .ZN(n2272) );
  INV_X4 U1935 ( .A(n3022), .ZN(n2908) );
  INV_X4 U1936 ( .A(n3000), .ZN(n1449) );
  INV_X4 U1937 ( .A(n4332), .ZN(n1370) );
  INV_X4 U1939 ( .A(n2982), .ZN(n2974) );
  INV_X2 U1940 ( .A(n2394), .ZN(n1748) );
  NAND3_X2 U1941 ( .A1(n3180), .A2(n3186), .A3(n3181), .ZN(n3184) );
  NAND2_X2 U1942 ( .A1(n3178), .A2(n3179), .ZN(n3180) );
  NAND3_X2 U1943 ( .A1(n4469), .A2(n4245), .A3(n1946), .ZN(n4246) );
  INV_X4 U1944 ( .A(n1945), .ZN(n1946) );
  NAND2_X2 U1945 ( .A1(n4242), .A2(net328272), .ZN(n4247) );
  NOR2_X2 U1947 ( .A1(n4240), .A2(n4239), .ZN(net328274) );
  INV_X4 U1949 ( .A(net331299), .ZN(net331293) );
  INV_X8 U1951 ( .A(net328259), .ZN(net328254) );
  NAND2_X2 U1952 ( .A1(a[6]), .A2(n2032), .ZN(n2278) );
  NAND2_X2 U1953 ( .A1(n2218), .A2(net330834), .ZN(n2574) );
  INV_X4 U1954 ( .A(n2865), .ZN(n3125) );
  INV_X4 U1956 ( .A(net331086), .ZN(net331083) );
  NAND4_X2 U1957 ( .A1(n3056), .A2(n3055), .A3(a[15]), .A4(n2034), .ZN(n3350)
         );
  INV_X4 U1958 ( .A(n1617), .ZN(n1618) );
  INV_X4 U1959 ( .A(n3698), .ZN(n3781) );
  INV_X4 U1960 ( .A(net330457), .ZN(net330458) );
  INV_X4 U1961 ( .A(n3700), .ZN(n1783) );
  OAI211_X2 U1962 ( .C1(net330600), .C2(net330599), .A(net330601), .B(
        net330510), .ZN(net330598) );
  OAI22_X2 U1963 ( .A1(n1104), .A2(net330385), .B1(net330384), .B2(net330386), 
        .ZN(net330383) );
  NOR2_X2 U1964 ( .A1(net331212), .A2(net331213), .ZN(net331211) );
  AOI21_X2 U1965 ( .B1(n2354), .B2(n4436), .A(n2353), .ZN(n2356) );
  NAND2_X2 U1966 ( .A1(n2706), .A2(n2430), .ZN(n2752) );
  NAND2_X2 U1967 ( .A1(n2840), .A2(n2839), .ZN(n2703) );
  NAND2_X2 U1968 ( .A1(n3009), .A2(n3008), .ZN(n2704) );
  NOR2_X2 U1969 ( .A1(net334433), .A2(n3611), .ZN(n3614) );
  INV_X4 U1970 ( .A(n3001), .ZN(n1448) );
  OAI21_X2 U1971 ( .B1(n2883), .B2(n2882), .A(n2881), .ZN(n2884) );
  INV_X4 U1972 ( .A(n2341), .ZN(n2344) );
  NAND2_X2 U1973 ( .A1(n4166), .A2(n4165), .ZN(n4167) );
  INV_X4 U1974 ( .A(n3972), .ZN(n3977) );
  AOI21_X2 U1975 ( .B1(n1681), .B2(n4155), .A(n4153), .ZN(n4158) );
  NAND2_X2 U1976 ( .A1(n2629), .A2(n1905), .ZN(n2829) );
  INV_X8 U1977 ( .A(n3754), .ZN(n3761) );
  INV_X4 U1978 ( .A(n4311), .ZN(n1621) );
  NAND3_X2 U1979 ( .A1(control[1]), .A2(b[2]), .A3(control[0]), .ZN(n2042) );
  INV_X4 U1980 ( .A(net331269), .ZN(net332264) );
  NAND3_X2 U1981 ( .A1(net331221), .A2(n1511), .A3(n1512), .ZN(n1509) );
  NAND3_X2 U1982 ( .A1(net331169), .A2(net331170), .A3(n1566), .ZN(n1565) );
  INV_X4 U1983 ( .A(net331311), .ZN(net331307) );
  NAND2_X2 U1984 ( .A1(n4084), .A2(n4086), .ZN(n4140) );
  INV_X16 U1985 ( .A(n1513), .ZN(net331341) );
  NAND2_X2 U1987 ( .A1(n3674), .A2(control[1]), .ZN(n1841) );
  NAND2_X2 U1988 ( .A1(n3827), .A2(n3963), .ZN(n3828) );
  NOR2_X1 U1989 ( .A1(net331614), .A2(net328250), .ZN(n1613) );
  AOI21_X2 U1990 ( .B1(net328035), .B2(n4110), .A(n4109), .ZN(n4111) );
  NOR2_X1 U1991 ( .A1(net331614), .A2(n4108), .ZN(n4109) );
  OAI21_X2 U1992 ( .B1(n3496), .B2(n3493), .A(n3492), .ZN(n3499) );
  NOR2_X2 U1993 ( .A1(n3495), .A2(n3494), .ZN(n3497) );
  INV_X4 U1994 ( .A(n4226), .ZN(n3742) );
  AOI21_X2 U1995 ( .B1(net328035), .B2(n3818), .A(n3817), .ZN(n3819) );
  NOR2_X2 U1996 ( .A1(n3816), .A2(net331614), .ZN(n3817) );
  INV_X4 U1997 ( .A(n3936), .ZN(n4120) );
  NOR2_X2 U1998 ( .A1(n2626), .A2(n2823), .ZN(n2728) );
  OAI21_X2 U1999 ( .B1(n3503), .B2(n3502), .A(n4209), .ZN(n3841) );
  OAI21_X2 U2000 ( .B1(n3844), .B2(n3927), .A(n3929), .ZN(n3936) );
  NOR2_X1 U2001 ( .A1(n3930), .A2(n3928), .ZN(n3844) );
  OAI21_X2 U2002 ( .B1(n4122), .B2(n4121), .A(n4120), .ZN(n4123) );
  NOR2_X1 U2003 ( .A1(net328254), .A2(n4126), .ZN(n4122) );
  NOR2_X2 U2004 ( .A1(net328254), .A2(n4127), .ZN(n4121) );
  NOR2_X2 U2005 ( .A1(n4201), .A2(n4200), .ZN(n4202) );
  AOI21_X2 U2006 ( .B1(n4199), .B2(n4206), .A(net328118), .ZN(n4201) );
  NOR2_X2 U2007 ( .A1(n4198), .A2(n4197), .ZN(n4199) );
  NAND2_X2 U2008 ( .A1(n1579), .A2(net328110), .ZN(n1578) );
  NAND2_X1 U2009 ( .A1(a[19]), .A2(n2037), .ZN(n3855) );
  AND2_X4 U2010 ( .A1(a[14]), .A2(net331329), .ZN(n1330) );
  AND2_X2 U2011 ( .A1(a[16]), .A2(n2037), .ZN(n1331) );
  AND2_X4 U2012 ( .A1(product_in[28]), .A2(net331295), .ZN(n1332) );
  AND3_X4 U2013 ( .A1(n1640), .A2(net331092), .A3(n1345), .ZN(n1333) );
  AND2_X2 U2014 ( .A1(n2823), .A2(n2822), .ZN(n1334) );
  NAND3_X2 U2015 ( .A1(n2202), .A2(n2201), .A3(n2200), .ZN(net328068) );
  AND3_X4 U2016 ( .A1(n1514), .A2(n1515), .A3(n1516), .ZN(n1335) );
  AND3_X4 U2017 ( .A1(n2150), .A2(n2149), .A3(n2148), .ZN(n1336) );
  NAND2_X1 U2018 ( .A1(a[22]), .A2(net331323), .ZN(net328567) );
  AND2_X4 U2019 ( .A1(product_in[20]), .A2(net331293), .ZN(n1337) );
  AND2_X4 U2020 ( .A1(a[4]), .A2(net331307), .ZN(n1338) );
  AND2_X4 U2021 ( .A1(a[2]), .A2(net331323), .ZN(n1339) );
  AND2_X4 U2022 ( .A1(a[16]), .A2(n2032), .ZN(n1340) );
  INV_X4 U2023 ( .A(net329465), .ZN(net329754) );
  INV_X4 U2024 ( .A(n2975), .ZN(n2978) );
  AND2_X2 U2025 ( .A1(n4239), .A2(n3928), .ZN(n1341) );
  NAND4_X2 U2026 ( .A1(a[23]), .A2(n3789), .A3(n3863), .A4(n2034), .ZN(n3876)
         );
  INV_X2 U2027 ( .A(net331362), .ZN(net331363) );
  INV_X4 U2028 ( .A(net328030), .ZN(net331362) );
  INV_X4 U2029 ( .A(n4090), .ZN(n3814) );
  AND2_X4 U2030 ( .A1(a[24]), .A2(n1719), .ZN(n1342) );
  AND2_X4 U2031 ( .A1(product_in[16]), .A2(net331293), .ZN(n1343) );
  INV_X4 U2032 ( .A(n3745), .ZN(n4233) );
  AND2_X2 U2033 ( .A1(n2703), .A2(n4433), .ZN(n1344) );
  INV_X4 U2034 ( .A(net331299), .ZN(net331295) );
  AND2_X2 U2035 ( .A1(a[2]), .A2(a[3]), .ZN(n1345) );
  INV_X1 U2036 ( .A(net331613), .ZN(net331614) );
  AND2_X2 U2037 ( .A1(n2856), .A2(n2855), .ZN(n1346) );
  AND2_X4 U2038 ( .A1(a[0]), .A2(net331305), .ZN(n1347) );
  AND2_X2 U2039 ( .A1(n2042), .A2(n2041), .ZN(n1348) );
  OR2_X4 U2040 ( .A1(n1513), .A2(net334240), .ZN(n1349) );
  AND2_X4 U2041 ( .A1(net331329), .A2(a[27]), .ZN(n1350) );
  AND2_X2 U2042 ( .A1(n4228), .A2(n4120), .ZN(n1351) );
  INV_X4 U2043 ( .A(n2097), .ZN(n2051) );
  OR2_X2 U2044 ( .A1(n2656), .A2(n2651), .ZN(n1352) );
  AND2_X2 U2045 ( .A1(a[18]), .A2(n1719), .ZN(n1353) );
  NAND2_X2 U2046 ( .A1(a[12]), .A2(net331323), .ZN(n3097) );
  INV_X4 U2047 ( .A(n3901), .ZN(n3894) );
  AND2_X2 U2048 ( .A1(n3490), .A2(n3489), .ZN(n1355) );
  AND2_X2 U2049 ( .A1(a[21]), .A2(n2034), .ZN(n1356) );
  AND2_X2 U2050 ( .A1(n2734), .A2(n2724), .ZN(n1357) );
  NAND2_X2 U2051 ( .A1(a[18]), .A2(net331305), .ZN(n3948) );
  AND2_X2 U2052 ( .A1(n2448), .A2(n1713), .ZN(n1358) );
  NAND3_X2 U2053 ( .A1(n1709), .A2(n2745), .A3(n2531), .ZN(n2747) );
  INV_X8 U2054 ( .A(n1565), .ZN(n1567) );
  INV_X16 U2055 ( .A(n1567), .ZN(net331329) );
  INV_X16 U2056 ( .A(n1335), .ZN(net331323) );
  INV_X16 U2057 ( .A(n1336), .ZN(n2037) );
  INV_X4 U2058 ( .A(net331311), .ZN(net331305) );
  OAI21_X4 U2059 ( .B1(n3084), .B2(n1393), .A(n3186), .ZN(n3085) );
  XNOR2_X1 U2060 ( .A(n3309), .B(n3192), .ZN(product_out[18]) );
  NAND2_X2 U2061 ( .A1(n3501), .A2(n3490), .ZN(n3192) );
  AND2_X2 U2062 ( .A1(n3175), .A2(n3177), .ZN(n1359) );
  XNOR2_X2 U2063 ( .A(n3085), .B(n3086), .ZN(product_out[17]) );
  XNOR2_X2 U2064 ( .A(n3396), .B(n1219), .ZN(product_out[20]) );
  INV_X1 U2068 ( .A(n2903), .ZN(n1362) );
  INV_X2 U2069 ( .A(n3177), .ZN(n3179) );
  NAND3_X2 U2070 ( .A1(n2959), .A2(n3005), .A3(n2834), .ZN(n2835) );
  NAND2_X4 U2071 ( .A1(n2815), .A2(n2816), .ZN(n2819) );
  INV_X8 U2072 ( .A(n3836), .ZN(n3933) );
  AND2_X2 U2073 ( .A1(n2746), .A2(n2531), .ZN(n1363) );
  XNOR2_X2 U2074 ( .A(n3926), .B(n1660), .ZN(product_out[26]) );
  NAND2_X4 U2075 ( .A1(n1750), .A2(n1751), .ZN(n2397) );
  NAND2_X4 U2076 ( .A1(n1748), .A2(n1749), .ZN(n1751) );
  INV_X4 U2077 ( .A(n4365), .ZN(n2896) );
  NAND2_X2 U2078 ( .A1(n2900), .A2(n1247), .ZN(n3181) );
  NAND2_X4 U2079 ( .A1(n1443), .A2(n1444), .ZN(n1446) );
  INV_X2 U2080 ( .A(n2236), .ZN(n2237) );
  NAND2_X4 U2082 ( .A1(n1446), .A2(n1445), .ZN(n3393) );
  INV_X8 U2083 ( .A(n1696), .ZN(n1697) );
  NAND2_X4 U2084 ( .A1(n2317), .A2(n2316), .ZN(n2416) );
  NAND2_X2 U2085 ( .A1(n3020), .A2(n1935), .ZN(n3021) );
  INV_X4 U2086 ( .A(n2315), .ZN(n1882) );
  INV_X4 U2087 ( .A(net334415), .ZN(net333890) );
  NAND2_X4 U2088 ( .A1(n2536), .A2(n2541), .ZN(n2311) );
  XNOR2_X2 U2089 ( .A(n3169), .B(n3168), .ZN(n1365) );
  NAND2_X2 U2090 ( .A1(n1631), .A2(net332977), .ZN(n2204) );
  AOI211_X4 U2091 ( .C1(net332214), .C2(n1623), .A(n3855), .B(net328790), .ZN(
        n3807) );
  BUF_X4 U2092 ( .A(n3859), .Z(n1623) );
  NAND2_X4 U2093 ( .A1(n1628), .A2(n3954), .ZN(n4296) );
  NAND2_X4 U2094 ( .A1(n1804), .A2(n1805), .ZN(n1628) );
  NAND2_X2 U2096 ( .A1(n2944), .A2(n2943), .ZN(n2951) );
  XNOR2_X2 U2097 ( .A(n3716), .B(n3715), .ZN(n1366) );
  NAND2_X4 U2098 ( .A1(n3766), .A2(n3714), .ZN(n3715) );
  NAND2_X4 U2100 ( .A1(n4196), .A2(net331362), .ZN(n4207) );
  NAND2_X4 U2101 ( .A1(n3405), .A2(n3414), .ZN(n3168) );
  INV_X4 U2102 ( .A(n4151), .ZN(n4155) );
  NAND2_X4 U2103 ( .A1(n2486), .A2(n2387), .ZN(n2489) );
  OAI211_X4 U2104 ( .C1(net328576), .C2(n1517), .A(net328578), .B(net328579), 
        .ZN(n1367) );
  OAI211_X2 U2105 ( .C1(net328576), .C2(n1517), .A(net328578), .B(net328579), 
        .ZN(net328230) );
  NAND2_X2 U2106 ( .A1(net328230), .A2(net328568), .ZN(net328562) );
  AOI21_X4 U2107 ( .B1(n2572), .B2(n2571), .A(n2579), .ZN(n2581) );
  INV_X2 U2108 ( .A(n3375), .ZN(n3373) );
  NAND2_X4 U2109 ( .A1(n1682), .A2(n2706), .ZN(n2495) );
  XNOR2_X2 U2111 ( .A(n4049), .B(n4161), .ZN(n4056) );
  NAND2_X4 U2112 ( .A1(n4048), .A2(n4047), .ZN(n4049) );
  NAND2_X4 U2113 ( .A1(n2603), .A2(n2604), .ZN(n2957) );
  INV_X4 U2115 ( .A(n2974), .ZN(n1687) );
  INV_X8 U2116 ( .A(n2472), .ZN(n2785) );
  OAI221_X4 U2117 ( .B1(n3761), .B2(n1735), .C1(n3682), .C2(n3681), .A(n2016), 
        .ZN(n3716) );
  NAND2_X2 U2118 ( .A1(net331273), .A2(net331272), .ZN(net331862) );
  XNOR2_X2 U2119 ( .A(n4333), .B(n1370), .ZN(n1369) );
  NAND2_X2 U2120 ( .A1(net329593), .A2(n3110), .ZN(n3111) );
  INV_X2 U2121 ( .A(net329593), .ZN(net329858) );
  INV_X4 U2123 ( .A(net330033), .ZN(net330029) );
  NAND2_X2 U2124 ( .A1(n3356), .A2(n3439), .ZN(n3357) );
  INV_X2 U2125 ( .A(n3198), .ZN(n1674) );
  XNOR2_X2 U2126 ( .A(n2768), .B(n2767), .ZN(n2857) );
  NAND2_X4 U2127 ( .A1(n1510), .A2(n1371), .ZN(net330955) );
  INV_X4 U2128 ( .A(net331059), .ZN(n1372) );
  NAND2_X4 U2129 ( .A1(n1372), .A2(net331033), .ZN(n1371) );
  NAND2_X2 U2130 ( .A1(net331031), .A2(net331059), .ZN(n1510) );
  NAND2_X2 U2131 ( .A1(n2798), .A2(n4432), .ZN(n2799) );
  INV_X8 U2132 ( .A(net330025), .ZN(net330335) );
  NAND2_X4 U2133 ( .A1(n3618), .A2(n3433), .ZN(n3430) );
  NOR2_X4 U2134 ( .A1(n2701), .A2(n2700), .ZN(n2649) );
  NAND3_X2 U2135 ( .A1(n3617), .A2(n3616), .A3(n3615), .ZN(n1374) );
  NAND2_X2 U2136 ( .A1(n3610), .A2(net328856), .ZN(n3616) );
  INV_X4 U2137 ( .A(n2397), .ZN(n2395) );
  NOR2_X4 U2139 ( .A1(net329556), .A2(n1330), .ZN(net333569) );
  NAND2_X4 U2140 ( .A1(n1141), .A2(n3426), .ZN(n1836) );
  INV_X4 U2142 ( .A(n3339), .ZN(n1439) );
  NAND2_X2 U2143 ( .A1(n3416), .A2(n3683), .ZN(n3381) );
  OAI21_X4 U2144 ( .B1(n2744), .B2(n2743), .A(n2959), .ZN(n2812) );
  OAI22_X4 U2145 ( .A1(n1195), .A2(net331138), .B1(net331017), .B2(net331138), 
        .ZN(net331137) );
  XNOR2_X2 U2146 ( .A(n2768), .B(n2767), .ZN(n1423) );
  INV_X8 U2147 ( .A(n2668), .ZN(n2768) );
  NAND2_X1 U2148 ( .A1(a[13]), .A2(n2032), .ZN(n2669) );
  INV_X4 U2149 ( .A(n2669), .ZN(n2767) );
  NAND2_X2 U2150 ( .A1(n2424), .A2(n2746), .ZN(n2432) );
  NAND2_X4 U2151 ( .A1(n3858), .A2(n3857), .ZN(n3915) );
  INV_X4 U2152 ( .A(net328984), .ZN(n1599) );
  NAND2_X2 U2153 ( .A1(n1773), .A2(n3680), .ZN(n3681) );
  NAND2_X2 U2154 ( .A1(n4432), .A2(n2703), .ZN(n2798) );
  INV_X2 U2155 ( .A(n2555), .ZN(n1760) );
  NAND2_X2 U2156 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  INV_X4 U2157 ( .A(n2852), .ZN(n2688) );
  INV_X16 U2158 ( .A(a[3]), .ZN(net331201) );
  NAND2_X2 U2159 ( .A1(n2043), .A2(n1210), .ZN(n2207) );
  NOR2_X1 U2160 ( .A1(n4311), .A2(n4310), .ZN(n4313) );
  NAND3_X4 U2161 ( .A1(n3370), .A2(a[18]), .A3(n2034), .ZN(n3449) );
  NAND4_X4 U2162 ( .A1(net331192), .A2(n1311), .A3(b[24]), .A4(a[3]), .ZN(
        net331244) );
  NAND2_X4 U2163 ( .A1(n2484), .A2(n2485), .ZN(n2387) );
  XNOR2_X2 U2164 ( .A(n2938), .B(n3135), .ZN(n1375) );
  INV_X4 U2165 ( .A(n1375), .ZN(n2940) );
  NAND3_X4 U2166 ( .A1(n2937), .A2(n1487), .A3(n3132), .ZN(n2938) );
  NAND2_X4 U2168 ( .A1(a[3]), .A2(net331341), .ZN(net331031) );
  NAND2_X4 U2169 ( .A1(n1420), .A2(net330595), .ZN(n2472) );
  NAND2_X4 U2170 ( .A1(net331055), .A2(n2140), .ZN(n2348) );
  INV_X8 U2171 ( .A(n2217), .ZN(n2291) );
  NAND2_X4 U2172 ( .A1(net331017), .A2(n1563), .ZN(n1376) );
  INV_X4 U2173 ( .A(net334298), .ZN(net329558) );
  NAND2_X4 U2174 ( .A1(a[9]), .A2(net331343), .ZN(net330457) );
  INV_X4 U2175 ( .A(net331127), .ZN(n1597) );
  OAI221_X4 U2176 ( .B1(n2560), .B2(n2788), .C1(n2558), .C2(n2559), .A(n2919), 
        .ZN(n2591) );
  NAND2_X4 U2178 ( .A1(net331261), .A2(n2043), .ZN(n1377) );
  INV_X8 U2179 ( .A(n1377), .ZN(n2040) );
  OAI22_X4 U2180 ( .A1(n1568), .A2(net330850), .B1(net331359), .B2(net331091), 
        .ZN(net330834) );
  INV_X4 U2181 ( .A(a[6]), .ZN(net330850) );
  OAI21_X4 U2182 ( .B1(n1356), .B2(n1218), .A(n3775), .ZN(n3769) );
  AOI22_X4 U2183 ( .A1(net328035), .A2(b[18]), .B1(net331613), .B2(b[26]), 
        .ZN(n2069) );
  INV_X4 U2184 ( .A(n2573), .ZN(n2577) );
  NAND3_X4 U2185 ( .A1(n4005), .A2(a[23]), .A3(n1565), .ZN(net328385) );
  NAND2_X4 U2186 ( .A1(net331254), .A2(net331194), .ZN(n2076) );
  INV_X32 U2187 ( .A(b[25]), .ZN(net331194) );
  OAI22_X4 U2188 ( .A1(n3228), .A2(n1940), .B1(n3027), .B2(n4442), .ZN(n3068)
         );
  NOR2_X2 U2189 ( .A1(n1378), .A2(n1718), .ZN(n1379) );
  INV_X4 U2190 ( .A(a[14]), .ZN(n1378) );
  INV_X2 U2191 ( .A(n1379), .ZN(n2762) );
  OAI221_X4 U2192 ( .B1(n3776), .B2(n3775), .C1(n3774), .C2(n3773), .A(n3772), 
        .ZN(n3777) );
  NAND2_X1 U2193 ( .A1(net328385), .A2(n4147), .ZN(n4149) );
  AOI21_X2 U2194 ( .B1(n1840), .B2(n1839), .A(n1211), .ZN(n1380) );
  INV_X4 U2195 ( .A(n1380), .ZN(n3110) );
  NAND2_X4 U2196 ( .A1(n1381), .A2(n3044), .ZN(n3117) );
  INV_X4 U2197 ( .A(n2941), .ZN(n1381) );
  AOI21_X4 U2198 ( .B1(n3276), .B2(n3275), .A(net329552), .ZN(n3278) );
  INV_X4 U2199 ( .A(n3107), .ZN(n3276) );
  NAND3_X2 U2200 ( .A1(net330998), .A2(n1809), .A3(n1808), .ZN(net331127) );
  NAND2_X4 U2201 ( .A1(net331860), .A2(net331861), .ZN(net331863) );
  NAND3_X4 U2202 ( .A1(n4426), .A2(n1312), .A3(b[25]), .ZN(net331284) );
  INV_X8 U2203 ( .A(control[0]), .ZN(n1382) );
  INV_X16 U2204 ( .A(control[1]), .ZN(n1383) );
  NAND2_X4 U2205 ( .A1(net328860), .A2(net328861), .ZN(n1384) );
  NAND2_X2 U2206 ( .A1(n2003), .A2(net332018), .ZN(n2005) );
  INV_X2 U2207 ( .A(net328740), .ZN(n1385) );
  INV_X4 U2208 ( .A(n1385), .ZN(n1386) );
  INV_X4 U2209 ( .A(n3055), .ZN(n3053) );
  NAND2_X2 U2210 ( .A1(n1771), .A2(n3680), .ZN(n3476) );
  INV_X4 U2211 ( .A(net328871), .ZN(n1387) );
  NAND2_X4 U2212 ( .A1(net334298), .A2(net329340), .ZN(net329463) );
  NAND2_X2 U2213 ( .A1(net332946), .A2(net332947), .ZN(n1852) );
  OAI21_X2 U2214 ( .B1(n1606), .B2(net330039), .A(n4390), .ZN(n1389) );
  NAND2_X4 U2215 ( .A1(n3074), .A2(n1442), .ZN(n3087) );
  CLKBUF_X3 U2216 ( .A(n3200), .Z(n1442) );
  INV_X8 U2218 ( .A(n1439), .ZN(n1390) );
  NAND2_X4 U2219 ( .A1(n1977), .A2(n1978), .ZN(n3555) );
  NAND2_X2 U2220 ( .A1(n1978), .A2(n1977), .ZN(n1403) );
  INV_X8 U2221 ( .A(n2205), .ZN(n1881) );
  XNOR2_X2 U2222 ( .A(n1681), .B(n4155), .ZN(n1391) );
  INV_X4 U2223 ( .A(n1391), .ZN(n3999) );
  NAND2_X4 U2224 ( .A1(net328740), .A2(net328871), .ZN(n1392) );
  INV_X2 U2225 ( .A(n3082), .ZN(n1393) );
  INV_X4 U2226 ( .A(n1394), .ZN(n1395) );
  INV_X4 U2227 ( .A(n3956), .ZN(n1396) );
  INV_X4 U2229 ( .A(net328235), .ZN(net328229) );
  INV_X4 U2230 ( .A(n1398), .ZN(n1399) );
  NAND2_X2 U2231 ( .A1(net328921), .A2(net328922), .ZN(net328919) );
  XNOR2_X2 U2233 ( .A(n3482), .B(n1401), .ZN(n1400) );
  INV_X1 U2235 ( .A(n1423), .ZN(n2672) );
  NAND2_X4 U2236 ( .A1(net331478), .A2(net331479), .ZN(n2031) );
  INV_X4 U2237 ( .A(n4189), .ZN(n1832) );
  XNOR2_X2 U2238 ( .A(net328912), .B(net328751), .ZN(n1402) );
  NAND2_X1 U2239 ( .A1(a[19]), .A2(net331323), .ZN(net328916) );
  OAI21_X4 U2240 ( .B1(n3947), .B2(n3856), .A(n4086), .ZN(n3858) );
  NAND2_X2 U2243 ( .A1(n3601), .A2(n3678), .ZN(n3563) );
  INV_X1 U2244 ( .A(n1133), .ZN(n3818) );
  NAND2_X4 U2246 ( .A1(n1208), .A2(net331238), .ZN(n2057) );
  NAND4_X4 U2247 ( .A1(n4426), .A2(net331254), .A3(b[25]), .A4(a[2]), .ZN(
        net331238) );
  NAND2_X4 U2248 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  NOR3_X2 U2249 ( .A1(n3761), .A2(n1955), .A3(n3760), .ZN(n1408) );
  INV_X2 U2250 ( .A(net328869), .ZN(n1409) );
  NAND2_X2 U2251 ( .A1(n4438), .A2(n2188), .ZN(n2144) );
  NAND4_X2 U2252 ( .A1(net331238), .A2(net331237), .A3(n1176), .A4(n1202), 
        .ZN(n2050) );
  INV_X4 U2253 ( .A(n2644), .ZN(n1410) );
  NAND2_X2 U2254 ( .A1(n1604), .A2(n1603), .ZN(n1485) );
  BUF_X4 U2256 ( .A(n2168), .Z(n1724) );
  NAND2_X2 U2257 ( .A1(n2653), .A2(n2652), .ZN(n1416) );
  NAND2_X4 U2259 ( .A1(n2232), .A2(n2233), .ZN(n2355) );
  NAND2_X1 U2260 ( .A1(n2233), .A2(n2232), .ZN(n1912) );
  INV_X4 U2261 ( .A(n3889), .ZN(n1413) );
  INV_X8 U2262 ( .A(n1413), .ZN(n1414) );
  INV_X4 U2263 ( .A(n2788), .ZN(n1460) );
  NAND2_X1 U2264 ( .A1(a[7]), .A2(n2035), .ZN(n2440) );
  XNOR2_X2 U2265 ( .A(n2269), .B(n2203), .ZN(n2248) );
  INV_X8 U2266 ( .A(n2246), .ZN(n2269) );
  INV_X8 U2267 ( .A(n2247), .ZN(n2203) );
  NAND2_X2 U2268 ( .A1(net333530), .A2(net333531), .ZN(net328555) );
  INV_X2 U2269 ( .A(n3902), .ZN(n3903) );
  AOI21_X4 U2270 ( .B1(net328734), .B2(n3894), .A(net328736), .ZN(n3906) );
  NAND2_X2 U2271 ( .A1(n1254), .A2(n1126), .ZN(net332820) );
  INV_X4 U2273 ( .A(n2655), .ZN(n1816) );
  NAND2_X4 U2274 ( .A1(net330238), .A2(n1643), .ZN(n2655) );
  BUF_X4 U2275 ( .A(n2746), .Z(n1709) );
  INV_X4 U2276 ( .A(n2314), .ZN(n1883) );
  INV_X2 U2277 ( .A(n3899), .ZN(net328605) );
  INV_X2 U2278 ( .A(n2595), .ZN(n2593) );
  NAND2_X4 U2279 ( .A1(n2595), .A2(n2640), .ZN(n2698) );
  NAND2_X2 U2280 ( .A1(n2182), .A2(n1420), .ZN(net332855) );
  OAI21_X4 U2281 ( .B1(n1544), .B2(n1545), .A(net328582), .ZN(net328579) );
  INV_X8 U2283 ( .A(n2845), .ZN(n2844) );
  INV_X8 U2284 ( .A(n2468), .ZN(n2002) );
  XNOR2_X2 U2286 ( .A(n2955), .B(n3026), .ZN(n1419) );
  NAND3_X1 U2287 ( .A1(net328235), .A2(net328473), .A3(net328236), .ZN(
        net328563) );
  NAND2_X1 U2288 ( .A1(net328562), .A2(net328563), .ZN(n1851) );
  NAND2_X1 U2289 ( .A1(n3737), .A2(n3736), .ZN(n1421) );
  NAND2_X1 U2290 ( .A1(n2394), .A2(n2393), .ZN(n1750) );
  INV_X4 U2291 ( .A(n2365), .ZN(n1617) );
  NAND2_X4 U2293 ( .A1(n2692), .A2(n2691), .ZN(n2693) );
  INV_X1 U2294 ( .A(n1606), .ZN(net333944) );
  BUF_X4 U2295 ( .A(n3350), .Z(n1655) );
  NAND2_X4 U2296 ( .A1(n2122), .A2(n2121), .ZN(n2244) );
  INV_X2 U2297 ( .A(n2430), .ZN(n2533) );
  AOI22_X4 U2298 ( .A1(n2647), .A2(n2702), .B1(n2547), .B2(n1428), .ZN(n2598)
         );
  NAND2_X4 U2299 ( .A1(n2647), .A2(n4486), .ZN(n2648) );
  NAND2_X4 U2300 ( .A1(n2336), .A2(n2331), .ZN(n2337) );
  NAND2_X4 U2301 ( .A1(n2327), .A2(n2328), .ZN(n2331) );
  NAND2_X2 U2302 ( .A1(n3100), .A2(net329750), .ZN(n1831) );
  CLKBUF_X3 U2303 ( .A(net328149), .Z(net332378) );
  NAND2_X4 U2304 ( .A1(n2797), .A2(n2796), .ZN(net330043) );
  AOI21_X4 U2305 ( .B1(n3208), .B2(n1677), .A(n3206), .ZN(n3210) );
  NAND2_X4 U2306 ( .A1(n1732), .A2(n2827), .ZN(n2959) );
  NAND2_X4 U2307 ( .A1(n1440), .A2(n1441), .ZN(n1739) );
  NAND2_X4 U2309 ( .A1(n1424), .A2(n3805), .ZN(n1426) );
  NAND2_X4 U2310 ( .A1(n1425), .A2(n1426), .ZN(n4012) );
  INV_X4 U2311 ( .A(net328851), .ZN(n1424) );
  NAND2_X4 U2312 ( .A1(n4012), .A2(n4013), .ZN(n4086) );
  NAND2_X2 U2313 ( .A1(n3155), .A2(n3156), .ZN(n1859) );
  AOI22_X4 U2314 ( .A1(n3278), .A2(net329547), .B1(n3277), .B2(net333678), 
        .ZN(n3279) );
  NAND2_X4 U2315 ( .A1(n1477), .A2(n1478), .ZN(n1480) );
  INV_X8 U2316 ( .A(n3925), .ZN(n4130) );
  INV_X4 U2317 ( .A(n3580), .ZN(n3582) );
  INV_X2 U2319 ( .A(n2393), .ZN(n1749) );
  NAND2_X2 U2320 ( .A1(n1358), .A2(n2449), .ZN(n2455) );
  INV_X1 U2321 ( .A(n2684), .ZN(n2448) );
  INV_X2 U2322 ( .A(n2455), .ZN(n2451) );
  NAND2_X2 U2323 ( .A1(n1429), .A2(n3528), .ZN(n1431) );
  INV_X4 U2324 ( .A(n3467), .ZN(n1429) );
  INV_X4 U2325 ( .A(net329017), .ZN(n1432) );
  NAND2_X2 U2326 ( .A1(n3623), .A2(n3434), .ZN(n3436) );
  NAND2_X2 U2327 ( .A1(n4075), .A2(n1822), .ZN(n1436) );
  NAND2_X4 U2328 ( .A1(n1434), .A2(n1435), .ZN(n1437) );
  NAND2_X4 U2329 ( .A1(n1436), .A2(n1437), .ZN(n1700) );
  INV_X4 U2330 ( .A(n4075), .ZN(n1434) );
  INV_X4 U2331 ( .A(n1822), .ZN(n1435) );
  INV_X8 U2332 ( .A(net328741), .ZN(net329017) );
  NAND2_X4 U2333 ( .A1(n3375), .A2(n3376), .ZN(n3433) );
  INV_X4 U2334 ( .A(net330456), .ZN(net330459) );
  NAND2_X2 U2335 ( .A1(n4057), .A2(n4056), .ZN(n4156) );
  NAND2_X4 U2337 ( .A1(n3223), .A2(n3222), .ZN(n3327) );
  XNOR2_X2 U2338 ( .A(n3221), .B(n4386), .ZN(n3223) );
  OAI21_X4 U2339 ( .B1(n3247), .B2(n1447), .A(n1633), .ZN(n3268) );
  NOR2_X2 U2340 ( .A1(net331353), .A2(n2763), .ZN(n2764) );
  NAND2_X4 U2341 ( .A1(n1488), .A2(n1489), .ZN(n1491) );
  INV_X4 U2342 ( .A(net329472), .ZN(net329751) );
  INV_X2 U2343 ( .A(n3404), .ZN(n1444) );
  NAND3_X2 U2344 ( .A1(n3942), .A2(n3941), .A3(n1351), .ZN(n1639) );
  NOR2_X4 U2345 ( .A1(net329297), .A2(n1349), .ZN(net334239) );
  INV_X4 U2346 ( .A(a[18]), .ZN(net334240) );
  NAND2_X2 U2347 ( .A1(n3354), .A2(n3148), .ZN(n3355) );
  NAND2_X2 U2348 ( .A1(n3001), .A2(n3000), .ZN(n1450) );
  NAND2_X4 U2349 ( .A1(n1448), .A2(n1449), .ZN(n1451) );
  NAND2_X4 U2350 ( .A1(n1450), .A2(n1451), .ZN(n3003) );
  NAND2_X4 U2351 ( .A1(n2890), .A2(n2000), .ZN(n3001) );
  NAND2_X4 U2352 ( .A1(n2768), .A2(n2767), .ZN(n2856) );
  NAND2_X1 U2353 ( .A1(n1412), .A2(net328125), .ZN(n1454) );
  NAND2_X2 U2354 ( .A1(n1452), .A2(n1453), .ZN(n1455) );
  NAND2_X2 U2355 ( .A1(n1454), .A2(n1455), .ZN(product_out[30]) );
  INV_X4 U2356 ( .A(n4308), .ZN(n1452) );
  INV_X2 U2357 ( .A(net328125), .ZN(n1453) );
  NAND2_X4 U2358 ( .A1(n2223), .A2(n2222), .ZN(n2224) );
  OAI21_X2 U2359 ( .B1(n1217), .B2(n2436), .A(n2437), .ZN(n2368) );
  INV_X2 U2360 ( .A(n2782), .ZN(n1778) );
  OAI21_X4 U2361 ( .B1(n1400), .B2(net331295), .A(n4222), .ZN(n1657) );
  NAND2_X2 U2362 ( .A1(n3092), .A2(n3007), .ZN(n2975) );
  NAND2_X1 U2363 ( .A1(net331799), .A2(net329813), .ZN(n1457) );
  INV_X4 U2364 ( .A(net329813), .ZN(n1456) );
  INV_X4 U2365 ( .A(n1771), .ZN(n1459) );
  NAND2_X2 U2367 ( .A1(n3380), .A2(n3381), .ZN(n1463) );
  NAND2_X4 U2368 ( .A1(n1461), .A2(n1462), .ZN(n1464) );
  NAND2_X4 U2369 ( .A1(n1463), .A2(n1464), .ZN(n3593) );
  INV_X4 U2370 ( .A(n3381), .ZN(n1461) );
  INV_X4 U2371 ( .A(n3380), .ZN(n1462) );
  INV_X2 U2372 ( .A(n3612), .ZN(n3613) );
  INV_X8 U2373 ( .A(n2600), .ZN(n2749) );
  NAND2_X4 U2375 ( .A1(net333795), .A2(net331113), .ZN(net331032) );
  NAND2_X2 U2376 ( .A1(n1913), .A2(n3203), .ZN(n1915) );
  NAND2_X2 U2377 ( .A1(n2958), .A2(n2957), .ZN(n2743) );
  OAI21_X4 U2378 ( .B1(net329821), .B2(net332231), .A(net329737), .ZN(n1555)
         );
  NAND2_X4 U2379 ( .A1(net329592), .A2(net329593), .ZN(n3344) );
  NAND2_X4 U2380 ( .A1(n1781), .A2(n1782), .ZN(n3924) );
  INV_X4 U2381 ( .A(n2720), .ZN(n2718) );
  NAND2_X4 U2382 ( .A1(net329334), .A2(net329073), .ZN(net329398) );
  INV_X2 U2383 ( .A(net329545), .ZN(net329352) );
  NAND2_X4 U2384 ( .A1(n3161), .A2(n3297), .ZN(n3162) );
  AOI22_X4 U2386 ( .A1(n1954), .A2(n2523), .B1(n2523), .B2(net331293), .ZN(
        n2513) );
  NAND2_X4 U2387 ( .A1(n4137), .A2(net334167), .ZN(n4138) );
  NAND2_X1 U2388 ( .A1(n3195), .A2(n3408), .ZN(n1465) );
  BUF_X8 U2389 ( .A(n3195), .Z(n1678) );
  NAND2_X2 U2390 ( .A1(net331031), .A2(net333862), .ZN(net331029) );
  INV_X4 U2391 ( .A(n1715), .ZN(n3104) );
  NAND2_X1 U2392 ( .A1(n1331), .A2(n3471), .ZN(n1466) );
  NAND2_X2 U2393 ( .A1(n1467), .A2(n3558), .ZN(n3557) );
  INV_X4 U2394 ( .A(n1466), .ZN(n1467) );
  NAND2_X2 U2395 ( .A1(n3557), .A2(n3556), .ZN(n1470) );
  NAND2_X4 U2396 ( .A1(n1468), .A2(n1469), .ZN(n1471) );
  NAND2_X4 U2397 ( .A1(n1470), .A2(n1471), .ZN(n3601) );
  INV_X4 U2398 ( .A(n3557), .ZN(n1468) );
  INV_X4 U2399 ( .A(n3556), .ZN(n1469) );
  NAND2_X1 U2400 ( .A1(n3610), .A2(n1331), .ZN(n3556) );
  INV_X8 U2401 ( .A(n3601), .ZN(n3760) );
  OAI21_X2 U2402 ( .B1(net328254), .B2(n4252), .A(net328414), .ZN(n4132) );
  INV_X1 U2403 ( .A(n4252), .ZN(n4113) );
  INV_X4 U2404 ( .A(net328981), .ZN(net328983) );
  INV_X1 U2405 ( .A(net328254), .ZN(n1584) );
  INV_X4 U2406 ( .A(n2748), .ZN(n1472) );
  NAND2_X4 U2407 ( .A1(n1909), .A2(n4455), .ZN(n3512) );
  OAI21_X4 U2408 ( .B1(n1606), .B2(net330039), .A(net330142), .ZN(net329467)
         );
  INV_X1 U2409 ( .A(n2820), .ZN(n2730) );
  NAND2_X4 U2411 ( .A1(n4374), .A2(n4375), .ZN(net327996) );
  NAND2_X2 U2412 ( .A1(n4355), .A2(n4294), .ZN(net333311) );
  NAND2_X2 U2413 ( .A1(n2363), .A2(n1143), .ZN(n2364) );
  NAND2_X4 U2414 ( .A1(n2838), .A2(n4458), .ZN(n1926) );
  NAND2_X4 U2415 ( .A1(n2997), .A2(n2996), .ZN(n3194) );
  NAND2_X4 U2416 ( .A1(n1823), .A2(n1824), .ZN(n2996) );
  NAND2_X2 U2417 ( .A1(n2995), .A2(n1669), .ZN(n1823) );
  NOR2_X2 U2418 ( .A1(net329972), .A2(net329592), .ZN(net329981) );
  XOR2_X2 U2419 ( .A(n1678), .B(n1675), .Z(n1708) );
  INV_X4 U2420 ( .A(n1674), .ZN(n1675) );
  INV_X8 U2421 ( .A(net330512), .ZN(net330385) );
  NAND3_X1 U2422 ( .A1(n3666), .A2(n3665), .A3(net329055), .ZN(n4229) );
  INV_X2 U2423 ( .A(n3665), .ZN(n3668) );
  NAND2_X4 U2424 ( .A1(n4146), .A2(n1149), .ZN(n4269) );
  NAND2_X2 U2425 ( .A1(n4116), .A2(n4115), .ZN(n1475) );
  INV_X2 U2426 ( .A(n3940), .ZN(n3575) );
  NAND2_X1 U2427 ( .A1(n2891), .A2(n2975), .ZN(n1949) );
  INV_X2 U2428 ( .A(n2891), .ZN(n1948) );
  NAND2_X1 U2429 ( .A1(n2086), .A2(n4463), .ZN(n2090) );
  INV_X2 U2430 ( .A(n2831), .ZN(n2742) );
  OAI22_X2 U2431 ( .A1(n2344), .A2(n2343), .B1(n2342), .B2(n2344), .ZN(n2345)
         );
  NAND2_X4 U2432 ( .A1(n3592), .A2(n3593), .ZN(n3509) );
  OAI21_X2 U2434 ( .B1(n3764), .B2(n3603), .A(n3602), .ZN(n3660) );
  INV_X2 U2435 ( .A(net328109), .ZN(net328125) );
  INV_X16 U2437 ( .A(n2036), .ZN(n2035) );
  NAND2_X4 U2438 ( .A1(n1473), .A2(n1474), .ZN(n1476) );
  NAND2_X2 U2439 ( .A1(n1476), .A2(n1475), .ZN(product_out[28]) );
  INV_X4 U2440 ( .A(n4116), .ZN(n1473) );
  INV_X4 U2441 ( .A(n4115), .ZN(n1474) );
  NAND2_X4 U2442 ( .A1(net328855), .A2(net328856), .ZN(net328854) );
  NOR3_X2 U2443 ( .A1(n3957), .A2(n3956), .A3(n3814), .ZN(n3969) );
  NAND2_X2 U2444 ( .A1(n2500), .A2(n2499), .ZN(n1905) );
  NAND2_X4 U2445 ( .A1(n3559), .A2(n3560), .ZN(n3606) );
  AOI21_X4 U2446 ( .B1(n3924), .B2(net331299), .A(n4243), .ZN(n3925) );
  NAND2_X2 U2447 ( .A1(n1480), .A2(n1479), .ZN(product_out[31]) );
  INV_X4 U2448 ( .A(net327991), .ZN(n1477) );
  INV_X4 U2450 ( .A(n1303), .ZN(n1982) );
  NAND2_X4 U2451 ( .A1(n1949), .A2(n1950), .ZN(n2892) );
  INV_X8 U2452 ( .A(n4036), .ZN(n4037) );
  NAND3_X2 U2453 ( .A1(n3326), .A2(n3591), .A3(n3327), .ZN(n3328) );
  NAND2_X4 U2454 ( .A1(n3239), .A2(net329598), .ZN(n3240) );
  NAND2_X4 U2455 ( .A1(n2528), .A2(n1338), .ZN(n2724) );
  NOR2_X4 U2456 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  INV_X2 U2457 ( .A(n3333), .ZN(n1481) );
  INV_X4 U2458 ( .A(n1481), .ZN(n1482) );
  NAND2_X4 U2459 ( .A1(n1483), .A2(n1484), .ZN(n1486) );
  NAND2_X4 U2460 ( .A1(n1485), .A2(n1486), .ZN(n1602) );
  INV_X4 U2461 ( .A(n1603), .ZN(n1483) );
  INV_X4 U2462 ( .A(n1604), .ZN(n1484) );
  INV_X8 U2463 ( .A(n1602), .ZN(n1601) );
  NAND2_X2 U2464 ( .A1(n1772), .A2(net328856), .ZN(n3561) );
  INV_X4 U2466 ( .A(n1622), .ZN(n3213) );
  OAI211_X4 U2467 ( .C1(n1874), .C2(n2350), .A(n2349), .B(n2348), .ZN(n2352)
         );
  INV_X4 U2468 ( .A(n1588), .ZN(n1585) );
  AND2_X4 U2469 ( .A1(n3471), .A2(n3605), .ZN(n1959) );
  INV_X4 U2470 ( .A(n2972), .ZN(n2973) );
  INV_X8 U2471 ( .A(n4092), .ZN(n3826) );
  NAND2_X4 U2472 ( .A1(n3720), .A2(n3721), .ZN(n1630) );
  AND2_X2 U2474 ( .A1(n2032), .A2(a[9]), .ZN(n2284) );
  NAND2_X2 U2475 ( .A1(a[11]), .A2(n2032), .ZN(n2563) );
  NAND2_X2 U2476 ( .A1(n1706), .A2(n2611), .ZN(n2615) );
  INV_X8 U2477 ( .A(n2084), .ZN(n2092) );
  NAND2_X4 U2478 ( .A1(n4175), .A2(n4283), .ZN(n4284) );
  INV_X2 U2480 ( .A(n3476), .ZN(n1489) );
  NAND2_X2 U2481 ( .A1(n2222), .A2(n2362), .ZN(n1492) );
  NAND2_X2 U2482 ( .A1(n2205), .A2(n1493), .ZN(n2214) );
  INV_X4 U2483 ( .A(n1492), .ZN(n1493) );
  INV_X2 U2484 ( .A(n2214), .ZN(n1928) );
  NAND2_X1 U2485 ( .A1(n2213), .A2(n2214), .ZN(n1929) );
  NAND2_X2 U2486 ( .A1(n3919), .A2(n3918), .ZN(n1781) );
  NOR2_X2 U2487 ( .A1(n3956), .A2(n3847), .ZN(n3851) );
  NAND2_X2 U2488 ( .A1(n2958), .A2(n2959), .ZN(n2716) );
  NAND2_X4 U2489 ( .A1(n2546), .A2(n2644), .ZN(n2486) );
  NAND3_X4 U2490 ( .A1(net330752), .A2(net330863), .A3(n2354), .ZN(n2185) );
  NAND2_X2 U2492 ( .A1(net333045), .A2(net328168), .ZN(n4104) );
  XNOR2_X2 U2493 ( .A(n2952), .B(n4445), .ZN(n3230) );
  NAND2_X1 U2494 ( .A1(net329069), .A2(net329068), .ZN(n1494) );
  NAND2_X2 U2495 ( .A1(net328126), .A2(net328123), .ZN(n1497) );
  NAND2_X4 U2496 ( .A1(n1495), .A2(n1496), .ZN(n1498) );
  NAND2_X4 U2497 ( .A1(n1498), .A2(n1497), .ZN(net328109) );
  INV_X4 U2498 ( .A(net328126), .ZN(n1495) );
  INV_X4 U2499 ( .A(net328123), .ZN(n1496) );
  NAND2_X4 U2500 ( .A1(n1499), .A2(net329014), .ZN(n1501) );
  NAND2_X4 U2501 ( .A1(n1500), .A2(n1501), .ZN(net328922) );
  INV_X4 U2502 ( .A(net329070), .ZN(n1499) );
  NAND2_X4 U2503 ( .A1(net329071), .A2(n1388), .ZN(net329070) );
  NAND3_X2 U2504 ( .A1(net328742), .A2(net328741), .A3(n1386), .ZN(net329071)
         );
  NAND2_X4 U2505 ( .A1(n1108), .A2(n1502), .ZN(net328871) );
  INV_X4 U2506 ( .A(net329194), .ZN(n1502) );
  NAND2_X4 U2507 ( .A1(net329020), .A2(net329021), .ZN(net328742) );
  NAND3_X2 U2508 ( .A1(n1432), .A2(net328742), .A3(net328869), .ZN(net328752)
         );
  NAND3_X2 U2509 ( .A1(n1386), .A2(net328742), .A3(net328741), .ZN(net328734)
         );
  INV_X8 U2510 ( .A(net329072), .ZN(net329021) );
  NAND3_X2 U2511 ( .A1(net329020), .A2(n1388), .A3(net329021), .ZN(net329015)
         );
  NAND2_X4 U2512 ( .A1(net329073), .A2(net329019), .ZN(net329072) );
  NAND2_X4 U2513 ( .A1(net329018), .A2(net329019), .ZN(net328741) );
  NAND2_X4 U2514 ( .A1(n1503), .A2(net329194), .ZN(net328740) );
  INV_X4 U2515 ( .A(net329020), .ZN(net329225) );
  XNOR2_X2 U2516 ( .A(net329291), .B(n1433), .ZN(net329230) );
  NAND2_X4 U2517 ( .A1(net331284), .A2(n1200), .ZN(net331282) );
  NOR2_X4 U2518 ( .A1(net328173), .A2(net328174), .ZN(net328169) );
  XNOR2_X2 U2519 ( .A(net328169), .B(net328170), .ZN(net328149) );
  NAND2_X4 U2520 ( .A1(net328176), .A2(net331479), .ZN(net328174) );
  NAND2_X4 U2521 ( .A1(net328408), .A2(net331479), .ZN(net328147) );
  INV_X4 U2522 ( .A(net328177), .ZN(net328173) );
  NAND2_X4 U2524 ( .A1(net328177), .A2(net328176), .ZN(net331520) );
  INV_X2 U2526 ( .A(net328474), .ZN(net332891) );
  NAND2_X4 U2527 ( .A1(net328474), .A2(net328473), .ZN(net328470) );
  OAI21_X4 U2528 ( .B1(net328474), .B2(net328473), .A(net328406), .ZN(
        net328472) );
  XNOR2_X2 U2529 ( .A(net328570), .B(net328569), .ZN(net328405) );
  XOR2_X2 U2530 ( .A(net328608), .B(n1505), .Z(n1504) );
  NAND2_X4 U2531 ( .A1(net328597), .A2(n1507), .ZN(net328491) );
  NAND2_X1 U2532 ( .A1(net328385), .A2(n1507), .ZN(net328484) );
  NAND3_X1 U2533 ( .A1(net328485), .A2(net328564), .A3(net328385), .ZN(
        net328608) );
  INV_X4 U2534 ( .A(net328404), .ZN(net328473) );
  NAND2_X2 U2535 ( .A1(a[21]), .A2(net331305), .ZN(net328171) );
  INV_X2 U2536 ( .A(net328171), .ZN(net331479) );
  NAND2_X4 U2537 ( .A1(net332264), .A2(net332265), .ZN(n1508) );
  NAND2_X4 U2538 ( .A1(n1508), .A2(net332266), .ZN(net331263) );
  INV_X4 U2539 ( .A(net331270), .ZN(net332265) );
  NOR2_X4 U2540 ( .A1(net331143), .A2(net331271), .ZN(net331270) );
  NAND2_X2 U2541 ( .A1(net331269), .A2(net331270), .ZN(net332266) );
  NAND2_X4 U2542 ( .A1(net331862), .A2(net331863), .ZN(net331269) );
  OAI22_X4 U2543 ( .A1(net331086), .A2(net331143), .B1(net331145), .B2(
        net331144), .ZN(net331028) );
  NOR2_X2 U2544 ( .A1(net331245), .A2(net331143), .ZN(net331247) );
  INV_X1 U2545 ( .A(net331271), .ZN(net331277) );
  INV_X4 U2546 ( .A(net328472), .ZN(net332028) );
  NAND2_X4 U2547 ( .A1(net332820), .A2(net332821), .ZN(net329816) );
  INV_X2 U2548 ( .A(net329981), .ZN(net332819) );
  INV_X8 U2549 ( .A(net329859), .ZN(net329592) );
  NOR2_X4 U2550 ( .A1(net334441), .A2(net329815), .ZN(net329813) );
  OAI21_X2 U2551 ( .B1(net329819), .B2(net329456), .A(net329972), .ZN(
        net329971) );
  INV_X4 U2552 ( .A(net329972), .ZN(net329811) );
  XNOR2_X2 U2553 ( .A(net331072), .B(net331061), .ZN(net331059) );
  INV_X4 U2554 ( .A(net331031), .ZN(net331033) );
  INV_X16 U2555 ( .A(n1509), .ZN(n1513) );
  INV_X32 U2556 ( .A(n1513), .ZN(net331343) );
  INV_X16 U2557 ( .A(net328712), .ZN(net328035) );
  NAND4_X4 U2558 ( .A1(net331193), .A2(b[9]), .A3(control[1]), .A4(a[2]), .ZN(
        net331235) );
  INV_X32 U2559 ( .A(control[1]), .ZN(net331253) );
  AOI21_X1 U2560 ( .B1(net329043), .B2(n1383), .A(n1382), .ZN(net329918) );
  NAND4_X4 U2561 ( .A1(a[2]), .A2(b[17]), .A3(control[0]), .A4(net331200), 
        .ZN(net331237) );
  NAND2_X2 U2562 ( .A1(b[3]), .A2(net331299), .ZN(n1511) );
  NAND2_X4 U2564 ( .A1(control[0]), .A2(control[1]), .ZN(net328006) );
  NAND2_X2 U2565 ( .A1(n1494), .A2(net328584), .ZN(net329033) );
  INV_X4 U2566 ( .A(net328922), .ZN(net329069) );
  NAND2_X2 U2567 ( .A1(a[18]), .A2(net331323), .ZN(net329068) );
  INV_X4 U2568 ( .A(net329068), .ZN(net328921) );
  AOI22_X2 U2569 ( .A1(b[29]), .A2(net331613), .B1(b[21]), .B2(net328035), 
        .ZN(n1516) );
  NAND2_X2 U2570 ( .A1(b[5]), .A2(net331299), .ZN(n1515) );
  NAND2_X2 U2571 ( .A1(b[13]), .A2(net331362), .ZN(n1514) );
  NAND2_X4 U2572 ( .A1(net328593), .A2(n1384), .ZN(n1517) );
  NAND2_X4 U2575 ( .A1(n1518), .A2(net328861), .ZN(net328582) );
  XNOR2_X2 U2577 ( .A(net328864), .B(net328865), .ZN(net328860) );
  NAND2_X2 U2579 ( .A1(net328917), .A2(net328918), .ZN(net328911) );
  NAND3_X2 U2580 ( .A1(n1282), .A2(net328980), .A3(net328981), .ZN(net328937)
         );
  OAI211_X4 U2581 ( .C1(net331063), .C2(net331062), .A(net331064), .B(
        net333853), .ZN(net331061) );
  NAND3_X4 U2583 ( .A1(n1151), .A2(net331069), .A3(n1519), .ZN(net330650) );
  INV_X4 U2584 ( .A(net331132), .ZN(n1519) );
  NAND3_X2 U2585 ( .A1(net331069), .A2(net331070), .A3(n1519), .ZN(net331066)
         );
  NOR2_X4 U2586 ( .A1(net331263), .A2(net331264), .ZN(net331499) );
  INV_X4 U2587 ( .A(net331499), .ZN(net331131) );
  NAND2_X1 U2588 ( .A1(net330994), .A2(net331499), .ZN(net333915) );
  NAND2_X4 U2590 ( .A1(net331128), .A2(net331129), .ZN(net330994) );
  INV_X2 U2591 ( .A(net331130), .ZN(net331128) );
  INV_X4 U2592 ( .A(net331070), .ZN(n1520) );
  OAI21_X4 U2593 ( .B1(n1520), .B2(n1521), .A(net331132), .ZN(net330653) );
  OAI21_X4 U2594 ( .B1(n1520), .B2(n1521), .A(net331132), .ZN(net333853) );
  NAND2_X1 U2595 ( .A1(net334464), .A2(net331264), .ZN(net331262) );
  INV_X2 U2596 ( .A(net331264), .ZN(net331180) );
  NAND2_X2 U2597 ( .A1(n1522), .A2(net331129), .ZN(net331226) );
  AOI22_X2 U2598 ( .A1(net331178), .A2(net330991), .B1(n1522), .B2(net331129), 
        .ZN(net331177) );
  NAND4_X4 U2599 ( .A1(net331130), .A2(net331227), .A3(n4325), .A4(a[1]), .ZN(
        net330991) );
  NAND2_X2 U2600 ( .A1(net331227), .A2(net331130), .ZN(n1522) );
  NAND2_X4 U2601 ( .A1(net329337), .A2(n4462), .ZN(net329336) );
  NAND3_X4 U2602 ( .A1(net329336), .A2(net329334), .A3(n1523), .ZN(net329020)
         );
  OAI21_X4 U2603 ( .B1(net329461), .B2(net329462), .A(net329463), .ZN(
        net329337) );
  INV_X2 U2604 ( .A(net329337), .ZN(net329457) );
  NAND3_X2 U2605 ( .A1(net329466), .A2(net329465), .A3(net329464), .ZN(
        net329462) );
  AOI211_X4 U2606 ( .C1(n1389), .C2(n4485), .A(net329469), .B(net329470), .ZN(
        net329461) );
  INV_X4 U2607 ( .A(net329469), .ZN(net333577) );
  NAND2_X4 U2608 ( .A1(net329558), .A2(net329557), .ZN(net329338) );
  AOI21_X2 U2609 ( .B1(net329399), .B2(n4462), .A(net329397), .ZN(net329395)
         );
  NAND2_X4 U2610 ( .A1(net329399), .A2(n4462), .ZN(net329407) );
  NAND2_X4 U2611 ( .A1(net329463), .A2(net329338), .ZN(net329545) );
  INV_X4 U2612 ( .A(net329340), .ZN(net329557) );
  NAND2_X2 U2613 ( .A1(net329465), .A2(n4448), .ZN(net329549) );
  NAND2_X4 U2614 ( .A1(net329345), .A2(net329464), .ZN(net329750) );
  NAND3_X2 U2615 ( .A1(net334227), .A2(net329808), .A3(net329751), .ZN(
        net329803) );
  INV_X8 U2617 ( .A(net331282), .ZN(net331017) );
  NAND3_X4 U2618 ( .A1(control[0]), .A2(net331251), .A3(b[17]), .ZN(net331283)
         );
  INV_X32 U2619 ( .A(control[1]), .ZN(net329919) );
  NAND4_X4 U2620 ( .A1(a[3]), .A2(b[16]), .A3(control[0]), .A4(n1383), .ZN(
        net331243) );
  INV_X4 U2621 ( .A(b[17]), .ZN(net331195) );
  NAND2_X4 U2622 ( .A1(n1524), .A2(n1525), .ZN(net327992) );
  NAND2_X2 U2623 ( .A1(n1526), .A2(net327996), .ZN(n1525) );
  NOR2_X2 U2624 ( .A1(net327997), .A2(net327998), .ZN(n1526) );
  AOI21_X4 U2625 ( .B1(net327999), .B2(net328000), .A(n1527), .ZN(n1524) );
  AOI22_X2 U2626 ( .A1(n1534), .A2(net328003), .B1(n1529), .B2(n1530), .ZN(
        n1527) );
  NAND2_X2 U2627 ( .A1(net328003), .A2(net331293), .ZN(n1530) );
  INV_X4 U2628 ( .A(n1528), .ZN(n1529) );
  INV_X2 U2629 ( .A(n1529), .ZN(n1534) );
  NAND2_X2 U2630 ( .A1(net328003), .A2(n1529), .ZN(net327998) );
  OAI211_X1 U2631 ( .C1(net328029), .C2(net331363), .A(net328031), .B(n1531), 
        .ZN(n1528) );
  NAND2_X2 U2632 ( .A1(net331613), .A2(n1532), .ZN(n1531) );
  INV_X4 U2633 ( .A(n1533), .ZN(n1532) );
  MUX2_X2 U2634 ( .A(product_in[7]), .B(n1532), .S(net331299), .Z(
        product_out[7]) );
  NAND2_X2 U2635 ( .A1(net331362), .A2(n1532), .ZN(net330067) );
  NAND2_X2 U2636 ( .A1(net328035), .A2(n1532), .ZN(net329055) );
  XNOR2_X2 U2637 ( .A(net330876), .B(n1347), .ZN(n1533) );
  NAND2_X2 U2638 ( .A1(n1347), .A2(net330876), .ZN(net330786) );
  NAND2_X4 U2639 ( .A1(net329980), .A2(net329872), .ZN(net329455) );
  INV_X8 U2641 ( .A(n1535), .ZN(net329980) );
  INV_X2 U2642 ( .A(net329980), .ZN(net333802) );
  NAND2_X4 U2643 ( .A1(net329980), .A2(net329872), .ZN(net329990) );
  OAI211_X4 U2644 ( .C1(n1539), .C2(net334211), .A(n1536), .B(n4468), .ZN(
        n1535) );
  NAND2_X4 U2645 ( .A1(net330237), .A2(net330238), .ZN(n1537) );
  NOR2_X4 U2646 ( .A1(n4388), .A2(net329994), .ZN(net330379) );
  OAI22_X2 U2647 ( .A1(net330385), .A2(n1104), .B1(net330384), .B2(net330386), 
        .ZN(n1541) );
  INV_X4 U2648 ( .A(net330513), .ZN(net330386) );
  NAND2_X4 U2649 ( .A1(net330385), .A2(net330386), .ZN(net333621) );
  NAND2_X4 U2650 ( .A1(net330385), .A2(net330386), .ZN(net330510) );
  INV_X4 U2651 ( .A(net329872), .ZN(net329860) );
  NAND2_X4 U2652 ( .A1(n1540), .A2(net330330), .ZN(net329989) );
  NAND2_X4 U2653 ( .A1(net329988), .A2(net329989), .ZN(net332761) );
  NAND2_X2 U2654 ( .A1(net332668), .A2(n4468), .ZN(net330327) );
  XNOR2_X2 U2655 ( .A(net330331), .B(n1538), .ZN(n1540) );
  BUF_X8 U2656 ( .A(net330026), .Z(n1538) );
  INV_X8 U2657 ( .A(net330332), .ZN(net330026) );
  OAI21_X2 U2658 ( .B1(net330026), .B2(net333079), .A(net333315), .ZN(
        net330213) );
  NOR2_X4 U2659 ( .A1(n1156), .A2(net330026), .ZN(net330197) );
  OAI211_X2 U2660 ( .C1(net328230), .C2(net328229), .A(net328232), .B(
        net328231), .ZN(net328222) );
  NAND2_X4 U2661 ( .A1(n1367), .A2(net331477), .ZN(net328388) );
  OAI21_X4 U2662 ( .B1(net328983), .B2(net328982), .A(net328583), .ZN(
        net328936) );
  NOR2_X4 U2663 ( .A1(n1546), .A2(n1307), .ZN(net328578) );
  OAI21_X4 U2665 ( .B1(n1542), .B2(n1543), .A(net328573), .ZN(net328524) );
  INV_X4 U2666 ( .A(net328574), .ZN(n1543) );
  INV_X4 U2667 ( .A(net328575), .ZN(n1542) );
  NAND2_X2 U2668 ( .A1(net329033), .A2(net328919), .ZN(net328980) );
  NAND3_X2 U2669 ( .A1(net328855), .A2(net328856), .A3(net328919), .ZN(
        net328981) );
  NAND3_X4 U2670 ( .A1(net330246), .A2(net330247), .A3(net330245), .ZN(
        net330244) );
  OAI22_X4 U2671 ( .A1(n1551), .A2(net330741), .B1(net334385), .B2(net330247), 
        .ZN(net330705) );
  NAND3_X1 U2672 ( .A1(net330245), .A2(n1162), .A3(net330246), .ZN(net330406)
         );
  NAND2_X4 U2673 ( .A1(n1547), .A2(net333890), .ZN(net330246) );
  NAND2_X4 U2674 ( .A1(net330858), .A2(net333890), .ZN(net330808) );
  OAI21_X4 U2675 ( .B1(net333519), .B2(n1548), .A(net330614), .ZN(n1547) );
  NOR2_X4 U2676 ( .A1(n1549), .A2(n1550), .ZN(n1548) );
  INV_X4 U2677 ( .A(n1552), .ZN(n1550) );
  OAI21_X4 U2678 ( .B1(n1549), .B2(n1550), .A(net330746), .ZN(net330745) );
  NAND2_X2 U2679 ( .A1(net330748), .A2(n1553), .ZN(n1552) );
  NAND2_X2 U2680 ( .A1(net331033), .A2(net331034), .ZN(n1553) );
  INV_X1 U2681 ( .A(net331034), .ZN(net333862) );
  NAND2_X4 U2682 ( .A1(net331034), .A2(net331033), .ZN(net332977) );
  INV_X4 U2684 ( .A(n1554), .ZN(n1549) );
  NAND2_X2 U2685 ( .A1(net332977), .A2(net330751), .ZN(n1554) );
  INV_X4 U2686 ( .A(net333275), .ZN(net333519) );
  NAND2_X2 U2687 ( .A1(net330599), .A2(net334044), .ZN(net330245) );
  INV_X4 U2688 ( .A(net330752), .ZN(net330599) );
  NAND2_X4 U2689 ( .A1(net329816), .A2(net329817), .ZN(net329470) );
  NAND3_X2 U2690 ( .A1(net329966), .A2(net329968), .A3(net329967), .ZN(
        net329817) );
  NAND2_X4 U2691 ( .A1(net329816), .A2(net333894), .ZN(net329965) );
  NAND2_X4 U2692 ( .A1(n1456), .A2(net332819), .ZN(net332821) );
  NAND2_X2 U2693 ( .A1(net329978), .A2(n1557), .ZN(net329966) );
  NAND3_X2 U2694 ( .A1(net329966), .A2(net329967), .A3(net329968), .ZN(
        net333894) );
  INV_X4 U2695 ( .A(n1558), .ZN(n1557) );
  NAND2_X1 U2697 ( .A1(net329592), .A2(net329456), .ZN(n1558) );
  NAND3_X2 U2698 ( .A1(net332231), .A2(net329973), .A3(net329974), .ZN(
        net329967) );
  INV_X4 U2699 ( .A(n1556), .ZN(net332230) );
  OAI21_X4 U2700 ( .B1(net329452), .B2(net329453), .A(n1556), .ZN(net329985)
         );
  INV_X4 U2701 ( .A(net329973), .ZN(net329819) );
  NOR2_X4 U2702 ( .A1(net330861), .A2(net330912), .ZN(net334415) );
  INV_X4 U2703 ( .A(net330912), .ZN(net330859) );
  NAND3_X1 U2704 ( .A1(net330854), .A2(n4451), .A3(net330859), .ZN(net330917)
         );
  NAND2_X1 U2705 ( .A1(net330856), .A2(net330859), .ZN(net330916) );
  NAND2_X4 U2706 ( .A1(net334334), .A2(net330912), .ZN(net330614) );
  NAND2_X4 U2707 ( .A1(net330745), .A2(net330614), .ZN(net330600) );
  NAND2_X2 U2708 ( .A1(a[1]), .A2(n1376), .ZN(net331273) );
  NAND2_X4 U2709 ( .A1(net331017), .A2(n1194), .ZN(net330839) );
  NOR2_X4 U2710 ( .A1(n1560), .A2(n1559), .ZN(n1564) );
  INV_X8 U2711 ( .A(n1562), .ZN(n1559) );
  NOR2_X4 U2712 ( .A1(n1560), .A2(n1559), .ZN(n1563) );
  NAND3_X4 U2713 ( .A1(control[0]), .A2(control[1]), .A3(b[1]), .ZN(n1562) );
  NAND3_X4 U2714 ( .A1(net331583), .A2(b[9]), .A3(control[1]), .ZN(n1561) );
  NAND3_X4 U2715 ( .A1(net332836), .A2(n1326), .A3(b[24]), .ZN(net331261) );
  NAND2_X4 U2716 ( .A1(net331017), .A2(n1564), .ZN(net331092) );
  NAND4_X4 U2717 ( .A1(control[1]), .A2(b[1]), .A3(control[0]), .A4(a[2]), 
        .ZN(net331234) );
  NOR2_X4 U2718 ( .A1(b[9]), .A2(control[0]), .ZN(net331199) );
  NAND3_X4 U2719 ( .A1(net329410), .A2(a[16]), .A3(net331329), .ZN(net329073)
         );
  NOR2_X4 U2720 ( .A1(n1568), .A2(net331212), .ZN(net331272) );
  INV_X4 U2721 ( .A(a[2]), .ZN(net331212) );
  INV_X8 U2722 ( .A(n2033), .ZN(n1568) );
  NAND2_X4 U2723 ( .A1(net330110), .A2(a[7]), .ZN(net330843) );
  OAI21_X4 U2724 ( .B1(net328128), .B2(net328127), .A(net328129), .ZN(
        net328126) );
  OAI221_X4 U2725 ( .B1(net328130), .B2(net328131), .C1(net328132), .C2(n1569), 
        .A(net328134), .ZN(net328129) );
  NOR3_X4 U2726 ( .A1(n1570), .A2(net328137), .A3(n1571), .ZN(net328134) );
  XNOR2_X2 U2727 ( .A(net328025), .B(net328024), .ZN(n1571) );
  NOR3_X4 U2728 ( .A1(net332747), .A2(n1572), .A3(net332583), .ZN(n1570) );
  INV_X8 U2729 ( .A(net328147), .ZN(net332583) );
  INV_X1 U2730 ( .A(net332583), .ZN(net332584) );
  INV_X4 U2731 ( .A(net328158), .ZN(n1572) );
  INV_X2 U2732 ( .A(n1572), .ZN(net331895) );
  AOI21_X4 U2733 ( .B1(net328148), .B2(net332378), .A(n1573), .ZN(n1569) );
  NOR3_X4 U2734 ( .A1(net328151), .A2(net333044), .A3(net328130), .ZN(n1573)
         );
  INV_X8 U2735 ( .A(net328167), .ZN(net333044) );
  INV_X4 U2736 ( .A(net328027), .ZN(net328130) );
  INV_X4 U2737 ( .A(net328149), .ZN(net328151) );
  NOR2_X2 U2738 ( .A1(net328151), .A2(net333044), .ZN(net328162) );
  NAND3_X2 U2739 ( .A1(net328168), .A2(net332378), .A3(net333045), .ZN(
        net328013) );
  INV_X4 U2740 ( .A(net332287), .ZN(net328132) );
  INV_X4 U2741 ( .A(net328026), .ZN(net328131) );
  NOR3_X2 U2742 ( .A1(net328137), .A2(net332747), .A3(net328182), .ZN(
        net328181) );
  XNOR2_X2 U2743 ( .A(net328183), .B(n1574), .ZN(net328182) );
  INV_X4 U2746 ( .A(net328083), .ZN(net328047) );
  XNOR2_X2 U2747 ( .A(net328046), .B(net328047), .ZN(net328019) );
  NAND2_X4 U2748 ( .A1(n1576), .A2(net329409), .ZN(net329334) );
  INV_X4 U2749 ( .A(n1373), .ZN(net329409) );
  NAND2_X2 U2750 ( .A1(a[16]), .A2(net331329), .ZN(n1576) );
  NAND2_X2 U2751 ( .A1(b[4]), .A2(net331299), .ZN(net331170) );
  NAND3_X2 U2752 ( .A1(net330862), .A2(net330614), .A3(net330752), .ZN(
        net330858) );
  XNOR2_X2 U2753 ( .A(net330913), .B(net330856), .ZN(net334334) );
  INV_X4 U2754 ( .A(net330925), .ZN(net330856) );
  NAND3_X2 U2755 ( .A1(net330854), .A2(n4451), .A3(net330856), .ZN(net330853)
         );
  XNOR2_X2 U2756 ( .A(net330913), .B(net330856), .ZN(net330861) );
  NAND2_X2 U2757 ( .A1(net330738), .A2(net330595), .ZN(net330925) );
  NAND2_X4 U2758 ( .A1(net332856), .A2(net332855), .ZN(net330748) );
  INV_X4 U2759 ( .A(net330748), .ZN(net330987) );
  NAND2_X4 U2760 ( .A1(n4450), .A2(net330751), .ZN(net330752) );
  NAND2_X2 U2761 ( .A1(net329811), .A2(net329456), .ZN(net329815) );
  NAND2_X4 U2762 ( .A1(net329818), .A2(net329811), .ZN(net329465) );
  OAI21_X4 U2763 ( .B1(net329452), .B2(net329453), .A(net333532), .ZN(
        net329451) );
  NAND2_X4 U2764 ( .A1(n1577), .A2(net328525), .ZN(net328167) );
  INV_X4 U2765 ( .A(net328528), .ZN(net328525) );
  XNOR2_X2 U2766 ( .A(net328527), .B(net332028), .ZN(n1577) );
  NAND2_X4 U2767 ( .A1(net332028), .A2(net328525), .ZN(net333531) );
  NAND2_X2 U2768 ( .A1(a[22]), .A2(net331305), .ZN(net328027) );
  NAND2_X2 U2769 ( .A1(net328026), .A2(net328027), .ZN(net328021) );
  NAND2_X1 U2770 ( .A1(net328528), .A2(net328472), .ZN(net333530) );
  XNOR2_X2 U2771 ( .A(net328555), .B(net328527), .ZN(net328160) );
  AOI21_X4 U2772 ( .B1(net328109), .B2(net328110), .A(net328111), .ZN(
        net327991) );
  AOI21_X4 U2773 ( .B1(net328113), .B2(net331938), .A(n1578), .ZN(net328111)
         );
  NAND2_X2 U2774 ( .A1(n1580), .A2(net328117), .ZN(n1579) );
  INV_X4 U2775 ( .A(net328118), .ZN(n1580) );
  INV_X4 U2776 ( .A(n1582), .ZN(n1581) );
  NAND2_X1 U2777 ( .A1(n1583), .A2(net328259), .ZN(n1582) );
  NAND3_X2 U2778 ( .A1(net328272), .A2(net328259), .A3(net328274), .ZN(
        net328264) );
  NAND3_X4 U2780 ( .A1(n1129), .A2(net332761), .A3(net332668), .ZN(net329453)
         );
  NAND3_X2 U2782 ( .A1(n1129), .A2(net332668), .A3(net330131), .ZN(net330128)
         );
  INV_X8 U2783 ( .A(net329868), .ZN(net332666) );
  OAI21_X4 U2784 ( .B1(n1585), .B2(n1586), .A(net330954), .ZN(net330746) );
  NAND3_X2 U2785 ( .A1(net330746), .A2(net334437), .A3(net330863), .ZN(
        net330862) );
  INV_X8 U2786 ( .A(net330955), .ZN(net330954) );
  OAI21_X4 U2787 ( .B1(n1585), .B2(n1586), .A(net330954), .ZN(net333275) );
  INV_X4 U2788 ( .A(n1587), .ZN(n1586) );
  NAND2_X4 U2789 ( .A1(n1589), .A2(n1590), .ZN(n1587) );
  NAND3_X2 U2790 ( .A1(net331032), .A2(n1587), .A3(net332977), .ZN(net330983)
         );
  XNOR2_X2 U2791 ( .A(net333618), .B(net331096), .ZN(n1590) );
  INV_X4 U2792 ( .A(net331098), .ZN(n1589) );
  NAND2_X4 U2793 ( .A1(net331113), .A2(n1591), .ZN(n1588) );
  XNOR2_X2 U2794 ( .A(n1593), .B(net331096), .ZN(n1591) );
  XNOR2_X2 U2795 ( .A(net331097), .B(net331098), .ZN(n1593) );
  XNOR2_X2 U2796 ( .A(n1592), .B(net331096), .ZN(net333795) );
  XNOR2_X2 U2797 ( .A(net331097), .B(net331098), .ZN(n1592) );
  XNOR2_X2 U2798 ( .A(net329690), .B(net329441), .ZN(n1594) );
  NAND2_X4 U2799 ( .A1(n1595), .A2(net328567), .ZN(net328236) );
  XNOR2_X2 U2800 ( .A(net328595), .B(net328596), .ZN(n1595) );
  OAI21_X4 U2801 ( .B1(net328612), .B2(n1596), .A(net328614), .ZN(net328487)
         );
  NAND2_X2 U2802 ( .A1(net328599), .A2(net328607), .ZN(n1596) );
  INV_X4 U2803 ( .A(net328617), .ZN(net328612) );
  NAND3_X2 U2804 ( .A1(net328601), .A2(net328603), .A3(net328602), .ZN(
        net328617) );
  XNOR2_X2 U2805 ( .A(net328331), .B(n4303), .ZN(net332558) );
  NAND2_X2 U2806 ( .A1(a[0]), .A2(n4325), .ZN(net331264) );
  NAND2_X2 U2807 ( .A1(a[1]), .A2(net331228), .ZN(net331129) );
  NOR2_X4 U2808 ( .A1(n1597), .A2(net331182), .ZN(net331176) );
  NAND2_X2 U2809 ( .A1(net330990), .A2(net333879), .ZN(net331063) );
  NAND3_X2 U2810 ( .A1(net330654), .A2(net330652), .A3(net333853), .ZN(
        net330730) );
  NAND2_X4 U2811 ( .A1(net331066), .A2(net330653), .ZN(net331097) );
  NAND2_X2 U2812 ( .A1(net331126), .A2(net331127), .ZN(net331123) );
  NAND3_X2 U2813 ( .A1(net330026), .A2(net333315), .A3(net330024), .ZN(
        net330021) );
  AOI21_X4 U2814 ( .B1(n1598), .B2(net330334), .A(net330335), .ZN(net330332)
         );
  NAND2_X4 U2815 ( .A1(net330459), .A2(net330458), .ZN(net330237) );
  INV_X4 U2816 ( .A(net330237), .ZN(net329988) );
  NAND2_X2 U2817 ( .A1(net334167), .A2(net328142), .ZN(net328475) );
  INV_X4 U2819 ( .A(net328567), .ZN(net328564) );
  NAND2_X2 U2820 ( .A1(a[25]), .A2(net331323), .ZN(net328051) );
  NAND2_X2 U2821 ( .A1(a[24]), .A2(net331323), .ZN(net328338) );
  NAND2_X2 U2822 ( .A1(a[23]), .A2(net331323), .ZN(net328392) );
  NAND2_X4 U2823 ( .A1(net328922), .A2(net328921), .ZN(net328584) );
  NAND2_X4 U2824 ( .A1(net332894), .A2(net332895), .ZN(net328918) );
  NAND2_X4 U2825 ( .A1(n1599), .A2(n1402), .ZN(net332895) );
  NAND2_X2 U2826 ( .A1(net328984), .A2(n1600), .ZN(net332894) );
  INV_X4 U2827 ( .A(net328916), .ZN(net328912) );
  OAI21_X1 U2828 ( .B1(net328750), .B2(net328751), .A(net328616), .ZN(
        net328748) );
  INV_X8 U2829 ( .A(net330037), .ZN(n1606) );
  NAND2_X4 U2830 ( .A1(n1601), .A2(net330044), .ZN(net329810) );
  NAND2_X2 U2831 ( .A1(net329876), .A2(net329593), .ZN(n1604) );
  AOI22_X4 U2832 ( .A1(net330127), .A2(net330126), .B1(net330128), .B2(n1605), 
        .ZN(n1603) );
  INV_X2 U2833 ( .A(net330130), .ZN(n1605) );
  NAND2_X4 U2835 ( .A1(net334039), .A2(n1610), .ZN(net331072) );
  INV_X8 U2837 ( .A(net330822), .ZN(n1611) );
  NAND3_X2 U2839 ( .A1(net330651), .A2(n1610), .A3(net330650), .ZN(net330204)
         );
  NAND2_X2 U2840 ( .A1(n1610), .A2(net330650), .ZN(net333614) );
  INV_X2 U2841 ( .A(n1610), .ZN(net330999) );
  INV_X4 U2842 ( .A(net331073), .ZN(n1609) );
  NAND2_X2 U2843 ( .A1(net330822), .A2(n1609), .ZN(net330649) );
  NAND2_X4 U2844 ( .A1(net330822), .A2(n1609), .ZN(n1610) );
  NAND2_X4 U2845 ( .A1(net328872), .A2(net328738), .ZN(net328873) );
  NAND3_X2 U2846 ( .A1(n1131), .A2(net328616), .A3(net328873), .ZN(net328866)
         );
  INV_X1 U2847 ( .A(net328738), .ZN(net328750) );
  OAI21_X4 U2848 ( .B1(net328245), .B2(net331363), .A(n1612), .ZN(net328137)
         );
  AOI21_X1 U2849 ( .B1(net328035), .B2(net328247), .A(n1613), .ZN(n1612) );
  XNOR2_X1 U2850 ( .A(n2129), .B(net331277), .ZN(n3816) );
  XOR2_X2 U2852 ( .A(n2312), .B(n2311), .Z(n1614) );
  OAI21_X4 U2853 ( .B1(n2271), .B2(n2272), .A(n1912), .ZN(n2312) );
  OAI21_X4 U2854 ( .B1(n2584), .B2(n1616), .A(n2855), .ZN(n1615) );
  NOR2_X1 U2855 ( .A1(net330942), .A2(n2583), .ZN(n1616) );
  NAND3_X4 U2857 ( .A1(n2075), .A2(net331196), .A3(net331198), .ZN(n2079) );
  XNOR2_X2 U2858 ( .A(n2490), .B(n2547), .ZN(n2494) );
  NAND3_X1 U2859 ( .A1(net331204), .A2(n2074), .A3(n2129), .ZN(n1620) );
  INV_X8 U2860 ( .A(n2784), .ZN(n2556) );
  CLKBUF_X3 U2861 ( .A(n3038), .Z(n1661) );
  INV_X4 U2862 ( .A(net330028), .ZN(net330377) );
  NOR2_X2 U2863 ( .A1(n1881), .A2(n2228), .ZN(n1960) );
  INV_X2 U2864 ( .A(n2562), .ZN(n2570) );
  XNOR2_X2 U2865 ( .A(n4310), .B(n1621), .ZN(n4321) );
  INV_X4 U2866 ( .A(n4309), .ZN(n4310) );
  NAND2_X4 U2867 ( .A1(n1423), .A2(n2856), .ZN(n3124) );
  INV_X1 U2868 ( .A(net331181), .ZN(net334464) );
  NAND2_X4 U2869 ( .A1(n1861), .A2(n1862), .ZN(n1864) );
  NOR2_X2 U2870 ( .A1(net331353), .A2(n2927), .ZN(n2928) );
  NOR2_X1 U2872 ( .A1(n4483), .A2(n3142), .ZN(n3143) );
  NOR2_X1 U2873 ( .A1(n4483), .A2(net329006), .ZN(n3699) );
  NAND2_X1 U2874 ( .A1(a[19]), .A2(net331349), .ZN(n3364) );
  NAND2_X1 U2875 ( .A1(a[21]), .A2(net331349), .ZN(n3538) );
  NAND2_X1 U2876 ( .A1(a[27]), .A2(net331349), .ZN(n4050) );
  NAND3_X2 U2877 ( .A1(n1342), .A2(a[23]), .A3(net331349), .ZN(n3779) );
  NAND3_X2 U2878 ( .A1(a[21]), .A2(n3540), .A3(net331349), .ZN(n3631) );
  NAND3_X2 U2879 ( .A1(a[19]), .A2(n3366), .A3(net331349), .ZN(n3453) );
  NAND3_X1 U2880 ( .A1(n1353), .A2(a[17]), .A3(net331349), .ZN(n3256) );
  OAI21_X2 U2881 ( .B1(n1353), .B2(n3143), .A(n3256), .ZN(n3251) );
  NAND2_X1 U2882 ( .A1(n3364), .A2(n3365), .ZN(n3367) );
  NAND2_X1 U2883 ( .A1(n3538), .A2(n3539), .ZN(n3541) );
  NAND2_X1 U2884 ( .A1(n4050), .A2(n4051), .ZN(n4053) );
  INV_X4 U2885 ( .A(n3047), .ZN(n3140) );
  INV_X2 U2886 ( .A(n3631), .ZN(n3634) );
  OAI21_X4 U2887 ( .B1(n3904), .B2(n3903), .A(net328616), .ZN(n3905) );
  NAND2_X1 U2888 ( .A1(a[17]), .A2(net331323), .ZN(n3554) );
  NAND2_X2 U2889 ( .A1(net330042), .A2(n2011), .ZN(n2914) );
  CLKBUF_X3 U2891 ( .A(n2341), .Z(n1626) );
  NAND2_X4 U2892 ( .A1(n2248), .A2(n1339), .ZN(n2341) );
  INV_X1 U2895 ( .A(n2656), .ZN(n1629) );
  INV_X4 U2896 ( .A(n2585), .ZN(n1766) );
  NAND2_X4 U2897 ( .A1(n2366), .A2(n1618), .ZN(n2367) );
  NAND2_X2 U2898 ( .A1(n2011), .A2(n3065), .ZN(n2802) );
  NAND2_X4 U2899 ( .A1(net330987), .A2(net330986), .ZN(n1631) );
  INV_X2 U2900 ( .A(net329033), .ZN(net333237) );
  INV_X4 U2901 ( .A(n1166), .ZN(n1632) );
  BUF_X16 U2902 ( .A(n3354), .Z(n1633) );
  NOR2_X4 U2903 ( .A1(n1635), .A2(n1333), .ZN(n1634) );
  AND3_X4 U2904 ( .A1(net331357), .A2(n2125), .A3(net331211), .ZN(n1635) );
  INV_X2 U2905 ( .A(n2797), .ZN(n2794) );
  INV_X4 U2906 ( .A(net332364), .ZN(net334385) );
  INV_X8 U2907 ( .A(n1104), .ZN(net332364) );
  INV_X4 U2908 ( .A(n2766), .ZN(n2850) );
  INV_X2 U2909 ( .A(n1637), .ZN(n1638) );
  NAND2_X2 U2910 ( .A1(n2002), .A2(n2757), .ZN(net333659) );
  NAND2_X4 U2911 ( .A1(n2939), .A2(n1375), .ZN(n2941) );
  NAND2_X4 U2913 ( .A1(n3706), .A2(n1237), .ZN(n3653) );
  INV_X8 U2915 ( .A(n2665), .ZN(n1736) );
  INV_X8 U2916 ( .A(n1615), .ZN(n2933) );
  INV_X8 U2917 ( .A(n2582), .ZN(n2584) );
  NAND2_X4 U2918 ( .A1(a[12]), .A2(n1719), .ZN(n2582) );
  OAI21_X4 U2919 ( .B1(n2830), .B2(n2829), .A(n2828), .ZN(n2831) );
  INV_X4 U2920 ( .A(n3505), .ZN(n3402) );
  NAND4_X2 U2921 ( .A1(n4120), .A2(n3942), .A3(n4228), .A4(n3941), .ZN(n4039)
         );
  INV_X2 U2922 ( .A(n2778), .ZN(n1664) );
  NAND2_X4 U2923 ( .A1(n2047), .A2(n2046), .ZN(n1640) );
  INV_X8 U2924 ( .A(n2080), .ZN(n2047) );
  CLKBUF_X2 U2926 ( .A(n3347), .Z(n1641) );
  INV_X1 U2927 ( .A(n4251), .ZN(n4200) );
  NAND2_X2 U2928 ( .A1(n3327), .A2(n3591), .ZN(n3330) );
  NAND2_X2 U2930 ( .A1(n3766), .A2(n1957), .ZN(n1642) );
  NAND2_X2 U2931 ( .A1(net329598), .A2(n2951), .ZN(net329973) );
  NAND2_X4 U2932 ( .A1(net330459), .A2(net330458), .ZN(n1643) );
  INV_X1 U2933 ( .A(n4164), .ZN(n4166) );
  NAND2_X2 U2934 ( .A1(n3265), .A2(n3266), .ZN(n3440) );
  INV_X2 U2935 ( .A(n3266), .ZN(n3267) );
  NAND2_X2 U2936 ( .A1(n3264), .A2(n3361), .ZN(n3266) );
  XNOR2_X2 U2937 ( .A(net329559), .B(net329560), .ZN(net334298) );
  NAND2_X2 U2938 ( .A1(n3435), .A2(n3341), .ZN(net329560) );
  XNOR2_X2 U2939 ( .A(n3363), .B(n3454), .ZN(n3370) );
  NAND2_X4 U2940 ( .A1(n3367), .A2(n3453), .ZN(n3454) );
  NAND2_X4 U2942 ( .A1(n3826), .A2(n1666), .ZN(n3850) );
  NAND2_X2 U2943 ( .A1(net328388), .A2(n1397), .ZN(n1645) );
  INV_X16 U2944 ( .A(a[9]), .ZN(n2377) );
  OAI21_X4 U2945 ( .B1(n3088), .B2(n3087), .A(n1442), .ZN(n3171) );
  XNOR2_X2 U2947 ( .A(n2955), .B(n3101), .ZN(n1646) );
  INV_X4 U2949 ( .A(n2548), .ZN(n2551) );
  XNOR2_X2 U2950 ( .A(n2845), .B(n2842), .ZN(n1648) );
  INV_X2 U2951 ( .A(n3237), .ZN(n3238) );
  AOI21_X2 U2952 ( .B1(n3352), .B2(n3351), .A(n3246), .ZN(n3247) );
  CLKBUF_X2 U2953 ( .A(n3433), .Z(n1649) );
  INV_X8 U2954 ( .A(n2781), .ZN(n2656) );
  INV_X4 U2955 ( .A(n3694), .ZN(n3774) );
  NAND3_X2 U2956 ( .A1(n2129), .A2(n2074), .A3(net331204), .ZN(n2180) );
  NOR2_X2 U2957 ( .A1(n2660), .A2(n2788), .ZN(n1651) );
  INV_X4 U2958 ( .A(n1651), .ZN(n2650) );
  INV_X2 U2959 ( .A(n2918), .ZN(n2660) );
  NAND2_X2 U2960 ( .A1(net331084), .A2(net331204), .ZN(n2099) );
  NAND3_X2 U2961 ( .A1(n2790), .A2(n2552), .A3(n2789), .ZN(n1652) );
  INV_X8 U2962 ( .A(net334239), .ZN(net329112) );
  INV_X4 U2963 ( .A(net329295), .ZN(net329297) );
  XNOR2_X2 U2964 ( .A(n3283), .B(n3282), .ZN(n1653) );
  NAND2_X2 U2965 ( .A1(n3383), .A2(n3426), .ZN(n3282) );
  NAND2_X4 U2966 ( .A1(n4144), .A2(net328392), .ZN(net328231) );
  XNOR2_X2 U2967 ( .A(n4001), .B(n4002), .ZN(n1654) );
  INV_X8 U2968 ( .A(n2620), .ZN(n2623) );
  NAND2_X4 U2969 ( .A1(n2817), .A2(n2818), .ZN(n3177) );
  INV_X4 U2970 ( .A(n2817), .ZN(n2815) );
  OAI22_X4 U2971 ( .A1(net331363), .A2(net328250), .B1(net333424), .B2(
        net331293), .ZN(n2817) );
  NAND2_X4 U2972 ( .A1(n1664), .A2(n2776), .ZN(n2924) );
  XNOR2_X2 U2973 ( .A(n2186), .B(n2185), .ZN(n1694) );
  NAND2_X4 U2974 ( .A1(net328385), .A2(net328485), .ZN(net328596) );
  AOI21_X1 U2975 ( .B1(n3302), .B2(n4020), .A(n3491), .ZN(n3303) );
  NAND3_X2 U2976 ( .A1(n1363), .A2(n2745), .A3(n1682), .ZN(n2535) );
  NAND2_X4 U2977 ( .A1(n4460), .A2(n2492), .ZN(n2748) );
  INV_X2 U2978 ( .A(net328563), .ZN(net332947) );
  NAND2_X4 U2979 ( .A1(n3159), .A2(n3160), .ZN(n1656) );
  INV_X1 U2981 ( .A(n2540), .ZN(n2542) );
  OAI21_X2 U2982 ( .B1(n2270), .B2(n2247), .A(n2540), .ZN(n2271) );
  NAND2_X4 U2983 ( .A1(n1956), .A2(n3855), .ZN(n1957) );
  AOI21_X2 U2984 ( .B1(net328748), .B2(n3896), .A(n3895), .ZN(n3897) );
  NAND2_X4 U2986 ( .A1(product_in[21]), .A2(n3487), .ZN(n4209) );
  NAND2_X4 U2987 ( .A1(n3193), .A2(n1680), .ZN(n3672) );
  INV_X2 U2988 ( .A(n3934), .ZN(n1660) );
  NAND2_X4 U2989 ( .A1(n3216), .A2(n3222), .ZN(n3405) );
  NAND2_X4 U2990 ( .A1(n4487), .A2(n4080), .ZN(net334167) );
  INV_X4 U2991 ( .A(n3605), .ZN(n3688) );
  NAND2_X2 U2992 ( .A1(n1171), .A2(n2226), .ZN(n1900) );
  NAND2_X2 U2993 ( .A1(n3094), .A2(n3093), .ZN(n3407) );
  NAND2_X1 U2995 ( .A1(n2307), .A2(n2306), .ZN(n1663) );
  INV_X8 U2996 ( .A(n2358), .ZN(n2306) );
  AOI21_X2 U2997 ( .B1(n3578), .B2(n3402), .A(n1906), .ZN(n3403) );
  INV_X4 U2998 ( .A(n1665), .ZN(n1666) );
  AOI21_X4 U2999 ( .B1(n2908), .B2(n2910), .A(n2883), .ZN(n2913) );
  INV_X8 U3000 ( .A(n1630), .ZN(n3960) );
  NAND2_X4 U3001 ( .A1(n2807), .A2(n2808), .ZN(n1668) );
  NAND2_X2 U3002 ( .A1(n2016), .A2(n1773), .ZN(n3659) );
  NAND2_X2 U3003 ( .A1(n3658), .A2(n1979), .ZN(n1773) );
  INV_X2 U3004 ( .A(n1106), .ZN(n1669) );
  NAND2_X4 U3005 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  NAND4_X1 U3006 ( .A1(n4208), .A2(net328118), .A3(n4206), .A4(n4207), .ZN(
        n1670) );
  INV_X4 U3007 ( .A(net329343), .ZN(net329552) );
  XNOR2_X2 U3008 ( .A(n3195), .B(n3196), .ZN(n3199) );
  NAND2_X4 U3009 ( .A1(n2740), .A2(n2739), .ZN(n1671) );
  NAND2_X2 U3010 ( .A1(n2721), .A2(n2720), .ZN(n2739) );
  NAND2_X2 U3011 ( .A1(n1608), .A2(n2471), .ZN(n2438) );
  INV_X1 U3012 ( .A(n3933), .ZN(n1672) );
  XNOR2_X1 U3013 ( .A(n2616), .B(n1917), .ZN(n1733) );
  NAND2_X4 U3014 ( .A1(n2965), .A2(n1668), .ZN(n3205) );
  INV_X4 U3015 ( .A(n3027), .ZN(n1673) );
  INV_X2 U3016 ( .A(net328117), .ZN(net328309) );
  NAND2_X4 U3017 ( .A1(n2413), .A2(n1697), .ZN(n2399) );
  NAND2_X4 U3018 ( .A1(n1714), .A2(n3069), .ZN(n3406) );
  NAND2_X4 U3020 ( .A1(n3910), .A2(n3911), .ZN(n4139) );
  OAI22_X4 U3023 ( .A1(n3816), .A2(net331363), .B1(n3815), .B2(net331293), 
        .ZN(n2329) );
  INV_X4 U3024 ( .A(n2463), .ZN(n1844) );
  OAI21_X4 U3025 ( .B1(n3997), .B2(n1198), .A(n3995), .ZN(n1681) );
  NAND2_X4 U3026 ( .A1(n3874), .A2(n3873), .ZN(n3995) );
  INV_X1 U3027 ( .A(n1705), .ZN(n3082) );
  NAND2_X4 U3028 ( .A1(n3167), .A2(n3166), .ZN(n3169) );
  NAND2_X4 U3029 ( .A1(n4460), .A2(n2492), .ZN(n1682) );
  NAND2_X1 U3031 ( .A1(net328179), .A2(net331506), .ZN(n4192) );
  INV_X8 U3032 ( .A(n2459), .ZN(n2659) );
  NAND2_X2 U3033 ( .A1(net331181), .A2(net331180), .ZN(net331178) );
  INV_X4 U3034 ( .A(n3586), .ZN(n1684) );
  XNOR2_X2 U3035 ( .A(n4290), .B(n4344), .ZN(n1685) );
  INV_X4 U3036 ( .A(n1685), .ZN(n4293) );
  INV_X2 U3037 ( .A(n4258), .ZN(n1686) );
  INV_X2 U3038 ( .A(n4363), .ZN(n4258) );
  INV_X4 U3039 ( .A(net328172), .ZN(net331478) );
  INV_X1 U3041 ( .A(n2425), .ZN(n2427) );
  INV_X8 U3043 ( .A(n3686), .ZN(n3515) );
  INV_X8 U3045 ( .A(n2979), .ZN(n2825) );
  XNOR2_X1 U3046 ( .A(n2905), .B(n2904), .ZN(product_out[15]) );
  OAI21_X1 U3047 ( .B1(n1118), .B2(net331363), .A(n3301), .ZN(n3491) );
  AOI21_X2 U3048 ( .B1(n3495), .B2(n3494), .A(n3491), .ZN(n3492) );
  INV_X2 U3049 ( .A(n1733), .ZN(n4110) );
  XOR2_X2 U3051 ( .A(net328020), .B(net328083), .Z(n1690) );
  BUF_X4 U3052 ( .A(n3019), .Z(n1935) );
  NAND2_X4 U3053 ( .A1(n3479), .A2(n3478), .ZN(n3579) );
  OAI21_X2 U3054 ( .B1(n1359), .B2(n2905), .A(n3181), .ZN(n2906) );
  NAND2_X1 U3055 ( .A1(n2798), .A2(n2755), .ZN(n2696) );
  NAND2_X4 U3056 ( .A1(n2745), .A2(n1709), .ZN(n2390) );
  NAND2_X2 U3057 ( .A1(net329112), .A2(n3623), .ZN(n2029) );
  NAND2_X4 U3058 ( .A1(n3428), .A2(n3429), .ZN(n3472) );
  OAI22_X1 U3059 ( .A1(n2823), .A2(n2822), .B1(n1984), .B2(n2820), .ZN(n1693)
         );
  OAI211_X4 U3060 ( .C1(n2729), .C2(n2728), .A(n2727), .B(n2726), .ZN(n2820)
         );
  INV_X1 U3061 ( .A(net328616), .ZN(net328615) );
  NAND2_X2 U3062 ( .A1(net328737), .A2(net328866), .ZN(n2022) );
  INV_X8 U3063 ( .A(n2908), .ZN(n1695) );
  INV_X4 U3064 ( .A(n2414), .ZN(n1696) );
  XNOR2_X2 U3065 ( .A(n4187), .B(n4186), .ZN(n1723) );
  OAI21_X2 U3066 ( .B1(n2676), .B2(n2288), .A(n2665), .ZN(n2445) );
  NAND2_X4 U3067 ( .A1(net329344), .A2(net329345), .ZN(n3277) );
  BUF_X32 U3068 ( .A(n2515), .Z(n1699) );
  NAND2_X2 U3069 ( .A1(net333915), .A2(net333879), .ZN(net331126) );
  INV_X4 U3070 ( .A(n1988), .ZN(n1822) );
  NAND2_X4 U3071 ( .A1(n3089), .A2(n3090), .ZN(n3071) );
  NOR2_X2 U3072 ( .A1(n1899), .A2(n2435), .ZN(n1701) );
  INV_X4 U3073 ( .A(n1701), .ZN(n2213) );
  NAND2_X4 U3074 ( .A1(a[6]), .A2(n4325), .ZN(n2435) );
  OAI211_X4 U3075 ( .C1(n3245), .C2(n3244), .A(n3243), .B(n3242), .ZN(
        net329559) );
  NAND2_X1 U3076 ( .A1(n2068), .A2(n2091), .ZN(n4022) );
  INV_X8 U3077 ( .A(n2048), .ZN(n2129) );
  INV_X1 U3079 ( .A(n2066), .ZN(n1703) );
  NAND2_X2 U3080 ( .A1(n1812), .A2(n1813), .ZN(n1704) );
  NAND2_X4 U3081 ( .A1(n1810), .A2(n1811), .ZN(n1813) );
  XNOR2_X2 U3082 ( .A(n3083), .B(n1343), .ZN(n1705) );
  NAND2_X2 U3083 ( .A1(n1630), .A2(n3732), .ZN(n1971) );
  INV_X4 U3084 ( .A(n3213), .ZN(n1707) );
  NAND3_X4 U3086 ( .A1(n2646), .A2(n1411), .A3(n2645), .ZN(n2647) );
  OAI21_X4 U3087 ( .B1(net329459), .B2(n3339), .A(net333678), .ZN(n3340) );
  XNOR2_X2 U3088 ( .A(n4465), .B(n2723), .ZN(n1954) );
  OAI21_X4 U3089 ( .B1(n2528), .B2(n1338), .A(n2506), .ZN(n2527) );
  INV_X8 U3090 ( .A(n2527), .ZN(n2723) );
  OAI22_X1 U3091 ( .A1(n2518), .A2(n2517), .B1(n1880), .B2(n1699), .ZN(n1710)
         );
  XNOR2_X1 U3092 ( .A(n2297), .B(n2296), .ZN(n1712) );
  OAI21_X4 U3093 ( .B1(n3358), .B2(n3357), .A(n3445), .ZN(n3372) );
  AOI21_X2 U3094 ( .B1(n3352), .B2(n3351), .A(n3444), .ZN(n3358) );
  INV_X1 U3095 ( .A(n2683), .ZN(n1713) );
  INV_X4 U3096 ( .A(n2450), .ZN(n2683) );
  INV_X4 U3097 ( .A(net330918), .ZN(net333869) );
  INV_X4 U3098 ( .A(net334039), .ZN(net330918) );
  XNOR2_X2 U3099 ( .A(n3068), .B(n3217), .ZN(n1714) );
  NAND2_X2 U3100 ( .A1(n3331), .A2(n1715), .ZN(n3217) );
  XNOR2_X2 U3101 ( .A(n3066), .B(n1831), .ZN(n1715) );
  NAND2_X4 U3102 ( .A1(a[3]), .A2(n4325), .ZN(net331132) );
  NAND2_X2 U3103 ( .A1(n2355), .A2(n2540), .ZN(n2236) );
  NAND2_X2 U3104 ( .A1(n1903), .A2(n1904), .ZN(n1717) );
  OAI21_X4 U3105 ( .B1(net328254), .B2(n4252), .A(n4251), .ZN(net328120) );
  OAI21_X4 U3106 ( .B1(n3609), .B2(n3688), .A(n3608), .ZN(n3617) );
  NAND4_X2 U3107 ( .A1(net331244), .A2(net331243), .A3(n1170), .A4(n2055), 
        .ZN(n2049) );
  INV_X4 U3108 ( .A(n2033), .ZN(n1718) );
  INV_X16 U3109 ( .A(n1718), .ZN(n1719) );
  OAI211_X4 U3110 ( .C1(n2439), .C2(n2438), .A(n2555), .B(n2556), .ZN(n1720)
         );
  NAND2_X4 U3111 ( .A1(n2276), .A2(n1354), .ZN(n1721) );
  NAND2_X2 U3114 ( .A1(n3662), .A2(n3661), .ZN(n3961) );
  NAND3_X2 U3116 ( .A1(net332364), .A2(net333621), .A3(n2548), .ZN(n1722) );
  OAI22_X4 U3117 ( .A1(n4150), .A2(n4149), .B1(n4270), .B2(n4268), .ZN(n4187)
         );
  XOR2_X2 U3119 ( .A(net330808), .B(n2469), .Z(n1726) );
  NAND2_X2 U3120 ( .A1(n1663), .A2(n1712), .ZN(n2469) );
  XNOR2_X2 U3121 ( .A(n3467), .B(n3527), .ZN(n1727) );
  OAI21_X4 U3122 ( .B1(n3764), .B2(n1459), .A(n3762), .ZN(n1729) );
  OAI21_X2 U3123 ( .B1(n3764), .B2(n1459), .A(n1408), .ZN(n4087) );
  INV_X1 U3124 ( .A(n3133), .ZN(n1731) );
  INV_X4 U3125 ( .A(n3050), .ZN(n3133) );
  XNOR2_X2 U3126 ( .A(n2712), .B(n2713), .ZN(n1732) );
  NAND2_X4 U3127 ( .A1(n2705), .A2(n2886), .ZN(n2713) );
  NAND2_X2 U3128 ( .A1(net328607), .A2(net328601), .ZN(net328864) );
  NAND2_X4 U3129 ( .A1(n2329), .A2(n2330), .ZN(n2336) );
  INV_X4 U3130 ( .A(n2329), .ZN(n2327) );
  INV_X8 U3131 ( .A(n1734), .ZN(n1735) );
  XNOR2_X2 U3133 ( .A(n2806), .B(n2805), .ZN(n1737) );
  XNOR2_X2 U3134 ( .A(n1231), .B(n4395), .ZN(n1740) );
  XNOR2_X2 U3135 ( .A(n2095), .B(n2134), .ZN(n1741) );
  NAND2_X2 U3136 ( .A1(n2731), .A2(n2615), .ZN(n2732) );
  NAND3_X2 U3137 ( .A1(n3101), .A2(n1673), .A3(n1850), .ZN(n3220) );
  INV_X1 U3138 ( .A(n4037), .ZN(n1742) );
  NAND2_X4 U3140 ( .A1(n3292), .A2(n3291), .ZN(n3325) );
  NAND2_X2 U3141 ( .A1(net330456), .A2(net330457), .ZN(net330238) );
  NAND2_X2 U3142 ( .A1(n2383), .A2(n2382), .ZN(n1746) );
  NAND2_X4 U3143 ( .A1(n1744), .A2(n1745), .ZN(n1747) );
  NAND2_X4 U3144 ( .A1(n1746), .A2(n1747), .ZN(net330512) );
  INV_X4 U3145 ( .A(n2383), .ZN(n1744) );
  INV_X8 U3148 ( .A(n2780), .ZN(n2788) );
  INV_X8 U3149 ( .A(n2773), .ZN(n2671) );
  AOI21_X2 U3150 ( .B1(n3899), .B2(n3900), .A(n4009), .ZN(n3898) );
  NAND2_X4 U3151 ( .A1(n3296), .A2(n3297), .ZN(n3321) );
  INV_X4 U3152 ( .A(n2353), .ZN(n1874) );
  OAI211_X2 U3153 ( .C1(n2836), .C2(n4424), .A(n2881), .B(n1695), .ZN(n2885)
         );
  NAND2_X4 U3154 ( .A1(net330853), .A2(n2274), .ZN(n2297) );
  INV_X2 U3155 ( .A(net330738), .ZN(net330737) );
  NAND2_X4 U3156 ( .A1(n3049), .A2(n1731), .ZN(n3056) );
  NAND2_X4 U3157 ( .A1(n2912), .A2(n2913), .ZN(n2955) );
  NAND2_X4 U3158 ( .A1(n3098), .A2(n3097), .ZN(n3331) );
  NAND2_X4 U3159 ( .A1(net329344), .A2(n4482), .ZN(n3339) );
  NAND2_X2 U3160 ( .A1(n2144), .A2(n2145), .ZN(n1754) );
  NAND2_X4 U3161 ( .A1(n1752), .A2(n1753), .ZN(n1755) );
  NAND2_X4 U3162 ( .A1(n1754), .A2(n1755), .ZN(n2192) );
  INV_X4 U3163 ( .A(n2145), .ZN(n1752) );
  INV_X4 U3164 ( .A(n2144), .ZN(n1753) );
  NOR2_X2 U3165 ( .A1(n4102), .A2(net331895), .ZN(n4103) );
  INV_X1 U3167 ( .A(n4391), .ZN(net328393) );
  NAND2_X4 U3168 ( .A1(n1212), .A2(n2940), .ZN(n3044) );
  XNOR2_X1 U3170 ( .A(n1416), .B(n2461), .ZN(n1756) );
  XNOR2_X2 U3171 ( .A(n4358), .B(n4357), .ZN(n1757) );
  AND2_X2 U3172 ( .A1(net328039), .A2(n4367), .ZN(n1758) );
  NAND2_X2 U3173 ( .A1(n2682), .A2(n2685), .ZN(n2687) );
  NAND2_X4 U3174 ( .A1(n2569), .A2(n2570), .ZN(n2769) );
  NAND4_X1 U3175 ( .A1(n1620), .A2(net330998), .A3(n2178), .A4(n1207), .ZN(
        net330654) );
  NAND2_X4 U3176 ( .A1(n3435), .A2(n3433), .ZN(n3524) );
  INV_X8 U3177 ( .A(n3524), .ZN(n3623) );
  INV_X4 U3178 ( .A(n3553), .ZN(n1976) );
  INV_X4 U3179 ( .A(n3471), .ZN(n3611) );
  NAND2_X4 U3180 ( .A1(n1308), .A2(net330239), .ZN(net329868) );
  NAND2_X2 U3181 ( .A1(n2560), .A2(n2477), .ZN(n2478) );
  NAND2_X2 U3182 ( .A1(n2479), .A2(n2478), .ZN(n1791) );
  INV_X8 U3183 ( .A(n2467), .ZN(n2468) );
  NAND2_X2 U3184 ( .A1(net328013), .A2(n4370), .ZN(n4372) );
  NAND2_X4 U3185 ( .A1(n1791), .A2(n1792), .ZN(n2480) );
  NAND2_X2 U3186 ( .A1(n3706), .A2(n1237), .ZN(n3650) );
  XNOR2_X1 U3187 ( .A(n4354), .B(n4353), .ZN(n4356) );
  INV_X4 U3189 ( .A(net330377), .ZN(net333079) );
  NAND2_X4 U3190 ( .A1(net330512), .A2(net330513), .ZN(n2467) );
  INV_X4 U3192 ( .A(n2379), .ZN(n1861) );
  NAND2_X2 U3193 ( .A1(n2379), .A2(n1827), .ZN(n1863) );
  XNOR2_X2 U3194 ( .A(n2704), .B(n1406), .ZN(n3011) );
  INV_X4 U3195 ( .A(net333614), .ZN(net333615) );
  INV_X8 U3197 ( .A(n4083), .ZN(n4142) );
  INV_X4 U3198 ( .A(n3205), .ZN(n3208) );
  NAND2_X2 U3199 ( .A1(n3811), .A2(n3810), .ZN(n1764) );
  NAND2_X4 U3200 ( .A1(n1762), .A2(n1763), .ZN(n1765) );
  NAND2_X4 U3201 ( .A1(n1764), .A2(n1765), .ZN(n4092) );
  INV_X4 U3202 ( .A(n3811), .ZN(n1762) );
  INV_X4 U3203 ( .A(n3810), .ZN(n1763) );
  INV_X1 U3204 ( .A(n3950), .ZN(n3810) );
  OAI21_X4 U3205 ( .B1(n4203), .B2(n1670), .A(n4202), .ZN(n4204) );
  NAND2_X2 U3206 ( .A1(n2933), .A2(n2585), .ZN(n1768) );
  NAND2_X4 U3207 ( .A1(n1766), .A2(n1767), .ZN(n1769) );
  NAND2_X4 U3208 ( .A1(n1768), .A2(n1769), .ZN(n2587) );
  INV_X8 U3209 ( .A(n2933), .ZN(n1767) );
  INV_X8 U3210 ( .A(n2386), .ZN(n2484) );
  INV_X8 U3211 ( .A(net333569), .ZN(net329344) );
  INV_X4 U3212 ( .A(n2826), .ZN(n2714) );
  INV_X4 U3213 ( .A(n2553), .ZN(n2380) );
  INV_X2 U3214 ( .A(n1699), .ZN(n2410) );
  NAND2_X4 U3215 ( .A1(n3999), .A2(n4000), .ZN(n4176) );
  OAI211_X4 U3216 ( .C1(n3448), .C2(n1793), .A(n3446), .B(n3445), .ZN(n3451)
         );
  INV_X4 U3217 ( .A(net327996), .ZN(net328000) );
  INV_X1 U3218 ( .A(n3986), .ZN(n3988) );
  INV_X1 U3219 ( .A(net331032), .ZN(net331115) );
  INV_X1 U3220 ( .A(n1420), .ZN(n1876) );
  INV_X4 U3222 ( .A(n4292), .ZN(n4291) );
  INV_X2 U3223 ( .A(n3051), .ZN(n3049) );
  NAND2_X2 U3224 ( .A1(n2627), .A2(n2629), .ZN(n2501) );
  INV_X8 U3225 ( .A(net329873), .ZN(net333532) );
  NAND2_X4 U3226 ( .A1(n4433), .A2(n4458), .ZN(net330039) );
  NAND2_X4 U3227 ( .A1(n3322), .A2(n1999), .ZN(n3323) );
  NAND2_X4 U3229 ( .A1(n2416), .A2(n2417), .ZN(n2400) );
  NAND2_X2 U3230 ( .A1(n4174), .A2(n4173), .ZN(n4283) );
  NAND2_X4 U3231 ( .A1(n4275), .A2(n4171), .ZN(n4276) );
  OAI211_X4 U3232 ( .C1(n3761), .C2(n1735), .A(n3757), .B(n3756), .ZN(n3759)
         );
  INV_X1 U3233 ( .A(n3689), .ZN(n1772) );
  XNOR2_X2 U3234 ( .A(n2562), .B(n2563), .ZN(n2450) );
  INV_X4 U3235 ( .A(net333500), .ZN(net333501) );
  INV_X8 U3236 ( .A(n2679), .ZN(n2561) );
  NAND2_X1 U3237 ( .A1(n2255), .A2(n2320), .ZN(n2199) );
  AND3_X4 U3238 ( .A1(n3490), .A2(n3489), .A3(n3488), .ZN(n1774) );
  NAND2_X4 U3239 ( .A1(n3183), .A2(n3080), .ZN(n3490) );
  OAI21_X4 U3240 ( .B1(n2337), .B2(n2338), .A(n1189), .ZN(n2339) );
  NAND2_X4 U3241 ( .A1(n2754), .A2(n2755), .ZN(n3023) );
  NAND3_X2 U3242 ( .A1(n2198), .A2(a[1]), .A3(n2037), .ZN(n2320) );
  INV_X4 U3243 ( .A(n2197), .ZN(n2198) );
  CLKBUF_X2 U3244 ( .A(n4271), .Z(n1775) );
  NAND2_X4 U3245 ( .A1(n3426), .A2(n3337), .ZN(n3514) );
  AND3_X4 U3246 ( .A1(n1153), .A2(n4464), .A3(n2780), .ZN(n2657) );
  INV_X4 U3247 ( .A(n3234), .ZN(n2027) );
  INV_X2 U3248 ( .A(n2454), .ZN(n2452) );
  NAND2_X2 U3249 ( .A1(n3638), .A2(n3637), .ZN(n3537) );
  NAND2_X4 U3250 ( .A1(net331123), .A2(n2138), .ZN(net331096) );
  OAI21_X2 U3251 ( .B1(n3952), .B2(n3956), .A(n4296), .ZN(n3953) );
  OAI21_X4 U3252 ( .B1(n2671), .B2(n2670), .A(n1395), .ZN(net330337) );
  INV_X2 U3253 ( .A(n3016), .ZN(n2879) );
  INV_X32 U3254 ( .A(control[0]), .ZN(net331193) );
  NAND3_X2 U3255 ( .A1(n3004), .A2(n1636), .A3(n3005), .ZN(n3006) );
  NAND2_X4 U3257 ( .A1(n3466), .A2(net329297), .ZN(n3619) );
  INV_X8 U3258 ( .A(n3865), .ZN(n3984) );
  OAI211_X4 U3259 ( .C1(n2688), .C2(n2687), .A(n2933), .B(n2932), .ZN(n2689)
         );
  NAND2_X4 U3260 ( .A1(n2413), .A2(n1697), .ZN(n2415) );
  NAND2_X4 U3261 ( .A1(n1711), .A2(n4009), .ZN(net328575) );
  AOI21_X2 U3262 ( .B1(n1337), .B2(n4211), .A(n4210), .ZN(n4220) );
  NAND2_X4 U3263 ( .A1(n3065), .A2(net329810), .ZN(net329472) );
  INV_X4 U3264 ( .A(net331938), .ZN(net331939) );
  INV_X8 U3265 ( .A(n3172), .ZN(n3922) );
  INV_X4 U3266 ( .A(n3005), .ZN(n3206) );
  NAND2_X4 U3267 ( .A1(n2395), .A2(n2396), .ZN(n2508) );
  NAND2_X4 U3268 ( .A1(n2146), .A2(n2193), .ZN(n2242) );
  OAI22_X4 U3269 ( .A1(n2618), .A2(n2617), .B1(n2621), .B2(n2622), .ZN(n2619)
         );
  XNOR2_X2 U3270 ( .A(n2825), .B(n2824), .ZN(net333424) );
  XNOR2_X2 U3271 ( .A(n3629), .B(n3547), .ZN(n3550) );
  INV_X2 U3272 ( .A(n3147), .ZN(n3145) );
  NAND3_X1 U3273 ( .A1(n4208), .A2(n4207), .A3(n4206), .ZN(net328117) );
  NAND2_X4 U3274 ( .A1(n3879), .A2(n3880), .ZN(n3883) );
  INV_X8 U3275 ( .A(n2637), .ZN(n2757) );
  NAND2_X4 U3277 ( .A1(n1779), .A2(n1780), .ZN(n1782) );
  INV_X4 U3278 ( .A(n3919), .ZN(n1779) );
  INV_X4 U3279 ( .A(n3918), .ZN(n1780) );
  XNOR2_X2 U3280 ( .A(n3698), .B(n1783), .ZN(n3702) );
  NAND2_X4 U3281 ( .A1(n2322), .A2(n2012), .ZN(n2413) );
  NAND2_X4 U3282 ( .A1(n2250), .A2(n2251), .ZN(n2012) );
  INV_X1 U3283 ( .A(n2923), .ZN(n1785) );
  NAND2_X4 U3284 ( .A1(n3978), .A2(n3883), .ZN(n3979) );
  NAND2_X4 U3285 ( .A1(n1654), .A2(n4003), .ZN(net328485) );
  NAND2_X1 U3287 ( .A1(net334044), .A2(net330509), .ZN(net330741) );
  NOR2_X4 U3288 ( .A1(n2473), .A2(n1352), .ZN(n2474) );
  NAND2_X4 U3289 ( .A1(n1789), .A2(n1790), .ZN(n1792) );
  INV_X4 U3290 ( .A(n2479), .ZN(n1789) );
  INV_X4 U3291 ( .A(n2478), .ZN(n1790) );
  NAND3_X2 U3292 ( .A1(a[22]), .A2(n3702), .A3(n2034), .ZN(n3772) );
  NAND2_X2 U3293 ( .A1(n3427), .A2(n3426), .ZN(n3519) );
  NAND2_X2 U3294 ( .A1(n3118), .A2(n3117), .ZN(n1793) );
  NAND2_X4 U3295 ( .A1(n3590), .A2(n3589), .ZN(n3592) );
  NAND2_X4 U3296 ( .A1(n3707), .A2(n3711), .ZN(n3705) );
  NAND2_X4 U3297 ( .A1(n3649), .A2(n3648), .ZN(n3711) );
  INV_X4 U3298 ( .A(n2612), .ZN(n2613) );
  NAND3_X4 U3299 ( .A1(n1420), .A2(n2364), .A3(net333869), .ZN(n2366) );
  INV_X2 U3300 ( .A(net333795), .ZN(net331119) );
  NAND3_X4 U3301 ( .A1(n2917), .A2(n2916), .A3(n2915), .ZN(n2952) );
  NAND4_X2 U3302 ( .A1(net330037), .A2(n3065), .A3(net329810), .A4(net330038), 
        .ZN(n2915) );
  NAND2_X2 U3303 ( .A1(n1132), .A2(n2644), .ZN(n2019) );
  NAND2_X4 U3304 ( .A1(n3108), .A2(n3109), .ZN(n3154) );
  NAND2_X2 U3305 ( .A1(n2191), .A2(n1196), .ZN(n1877) );
  INV_X4 U3306 ( .A(n2638), .ZN(n2639) );
  INV_X4 U3307 ( .A(n1120), .ZN(n1819) );
  INV_X1 U3308 ( .A(n4267), .ZN(n4273) );
  AOI21_X4 U3309 ( .B1(n2774), .B2(n2773), .A(n2772), .ZN(n2775) );
  INV_X2 U3310 ( .A(net332088), .ZN(net333336) );
  INV_X2 U3311 ( .A(net330040), .ZN(net332088) );
  NAND2_X4 U3313 ( .A1(n2840), .A2(n2839), .ZN(net330042) );
  NAND2_X4 U3314 ( .A1(a[14]), .A2(net331349), .ZN(n2862) );
  NAND2_X4 U3315 ( .A1(n2136), .A2(n1724), .ZN(n2137) );
  AOI21_X4 U3316 ( .B1(net334005), .B2(net332364), .A(n2468), .ZN(n2470) );
  INV_X8 U3317 ( .A(n2849), .ZN(n2665) );
  CLKBUF_X3 U3318 ( .A(net330025), .Z(net333315) );
  NAND2_X4 U3319 ( .A1(n2175), .A2(n2229), .ZN(n1828) );
  NAND2_X2 U3320 ( .A1(net331176), .A2(net331177), .ZN(n1796) );
  NAND2_X4 U3321 ( .A1(net333276), .A2(net333277), .ZN(n1797) );
  NAND2_X4 U3322 ( .A1(n1796), .A2(n1797), .ZN(n2084) );
  INV_X4 U3323 ( .A(net331176), .ZN(net333276) );
  INV_X4 U3324 ( .A(net331177), .ZN(net333277) );
  NAND2_X2 U3325 ( .A1(n2384), .A2(net330705), .ZN(n1799) );
  NAND2_X4 U3326 ( .A1(net333280), .A2(n1798), .ZN(n1800) );
  NAND2_X4 U3327 ( .A1(n1799), .A2(n1800), .ZN(n2386) );
  INV_X4 U3328 ( .A(net330705), .ZN(net333280) );
  INV_X4 U3329 ( .A(n2384), .ZN(n1798) );
  XNOR2_X2 U3330 ( .A(n4443), .B(n3385), .ZN(n1801) );
  NAND2_X2 U3331 ( .A1(n3915), .A2(n3914), .ZN(n1804) );
  NAND2_X4 U3332 ( .A1(n1802), .A2(n1803), .ZN(n1805) );
  INV_X4 U3333 ( .A(n3915), .ZN(n1802) );
  INV_X4 U3334 ( .A(n3914), .ZN(n1803) );
  NAND2_X4 U3336 ( .A1(n1806), .A2(n1807), .ZN(n1809) );
  NAND2_X4 U3337 ( .A1(n1809), .A2(n1808), .ZN(net331125) );
  INV_X4 U3338 ( .A(n2082), .ZN(n1806) );
  INV_X4 U3339 ( .A(n2178), .ZN(n1807) );
  NAND2_X4 U3340 ( .A1(n2386), .A2(n2385), .ZN(n2644) );
  NAND2_X2 U3341 ( .A1(n1138), .A2(n3517), .ZN(n3385) );
  NAND2_X4 U3342 ( .A1(net331125), .A2(net331124), .ZN(n2138) );
  NAND2_X4 U3343 ( .A1(net330131), .A2(net332668), .ZN(n2759) );
  NAND2_X4 U3344 ( .A1(n1318), .A2(net331351), .ZN(n2567) );
  NAND2_X4 U3345 ( .A1(n2373), .A2(n2372), .ZN(n2568) );
  AOI21_X1 U3346 ( .B1(n3276), .B2(n3275), .A(net329549), .ZN(n3273) );
  INV_X2 U3348 ( .A(n1692), .ZN(n3475) );
  CLKBUF_X3 U3349 ( .A(n2683), .Z(n1814) );
  OAI21_X4 U3350 ( .B1(n2447), .B2(n2684), .A(n1814), .ZN(n2454) );
  OAI211_X4 U3351 ( .C1(net333770), .C2(n2156), .A(n1145), .B(n2216), .ZN(
        net331069) );
  NAND2_X2 U3352 ( .A1(n2372), .A2(n2284), .ZN(n1812) );
  NAND2_X4 U3353 ( .A1(n1812), .A2(n1813), .ZN(n2443) );
  INV_X2 U3354 ( .A(n2372), .ZN(n1810) );
  INV_X4 U3355 ( .A(n2284), .ZN(n1811) );
  NAND2_X4 U3356 ( .A1(n2216), .A2(n2215), .ZN(n2217) );
  INV_X4 U3357 ( .A(n3628), .ZN(n3547) );
  NAND2_X4 U3358 ( .A1(n1815), .A2(n1816), .ZN(n1818) );
  NAND2_X4 U3359 ( .A1(n1817), .A2(n1818), .ZN(n2595) );
  INV_X4 U3360 ( .A(n2592), .ZN(n1815) );
  OAI221_X4 U3361 ( .B1(n2551), .B2(n2002), .C1(n4388), .C2(n1722), .A(n2550), 
        .ZN(n2592) );
  NOR2_X2 U3362 ( .A1(n2784), .A2(n2783), .ZN(n2790) );
  NAND2_X2 U3364 ( .A1(n1374), .A2(net329033), .ZN(n1820) );
  NAND2_X4 U3365 ( .A1(n1819), .A2(net333237), .ZN(n1821) );
  NAND2_X4 U3366 ( .A1(n1821), .A2(n1820), .ZN(n1979) );
  INV_X1 U3367 ( .A(net330942), .ZN(net333222) );
  NAND2_X4 U3368 ( .A1(n3619), .A2(net329112), .ZN(n3527) );
  INV_X4 U3369 ( .A(n4274), .ZN(n4277) );
  NAND3_X2 U3370 ( .A1(a[25]), .A2(n3868), .A3(net331351), .ZN(n3982) );
  INV_X4 U3371 ( .A(n2868), .ZN(n2870) );
  INV_X8 U3372 ( .A(n2275), .ZN(n2276) );
  NAND2_X2 U3373 ( .A1(n2292), .A2(n2572), .ZN(n2294) );
  INV_X2 U3375 ( .A(n4056), .ZN(n4054) );
  INV_X1 U3376 ( .A(n3783), .ZN(n3785) );
  NAND2_X4 U3377 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  NAND2_X4 U3378 ( .A1(n3195), .A2(n3408), .ZN(n3166) );
  NAND2_X4 U3379 ( .A1(net331235), .A2(net331234), .ZN(n2058) );
  INV_X8 U3380 ( .A(n2783), .ZN(n2555) );
  NAND2_X4 U3382 ( .A1(n2349), .A2(n2348), .ZN(n2247) );
  OAI21_X4 U3383 ( .B1(n2340), .B2(n2001), .A(n1983), .ZN(n2394) );
  NOR2_X4 U3384 ( .A1(n3016), .A2(n3015), .ZN(n3017) );
  NOR3_X4 U3385 ( .A1(n2579), .A2(n2578), .A3(n1736), .ZN(n2580) );
  NAND2_X2 U3386 ( .A1(n3058), .A2(n3116), .ZN(n1839) );
  NAND2_X2 U3387 ( .A1(n2164), .A2(net330843), .ZN(n1903) );
  OAI21_X4 U3388 ( .B1(n2289), .B2(n1736), .A(n2566), .ZN(n2374) );
  NAND2_X2 U3389 ( .A1(a[3]), .A2(n1376), .ZN(n2159) );
  NAND2_X2 U3390 ( .A1(n1698), .A2(n1106), .ZN(n1824) );
  NAND2_X4 U3391 ( .A1(n2529), .A2(n2530), .ZN(n2531) );
  INV_X2 U3392 ( .A(n4352), .ZN(n4353) );
  NAND2_X4 U3393 ( .A1(n3155), .A2(n3156), .ZN(n3335) );
  INV_X4 U3394 ( .A(n3406), .ZN(n1825) );
  INV_X4 U3395 ( .A(n1825), .ZN(n1826) );
  INV_X8 U3396 ( .A(net331028), .ZN(net331025) );
  NOR2_X1 U3397 ( .A1(n2681), .A2(n2849), .ZN(n2682) );
  INV_X2 U3398 ( .A(n2464), .ZN(n1843) );
  NAND2_X2 U3400 ( .A1(n2847), .A2(net329992), .ZN(net330127) );
  NAND2_X2 U3401 ( .A1(n2607), .A2(n1338), .ZN(n2504) );
  INV_X1 U3402 ( .A(n1862), .ZN(n1827) );
  XNOR2_X2 U3404 ( .A(n3066), .B(n1831), .ZN(n1830) );
  NAND2_X4 U3405 ( .A1(n2949), .A2(n2950), .ZN(n3028) );
  NAND2_X4 U3406 ( .A1(n3516), .A2(n3422), .ZN(n3429) );
  NAND2_X2 U3407 ( .A1(n3516), .A2(n3422), .ZN(n3604) );
  OAI21_X4 U3408 ( .B1(n2889), .B2(n2756), .A(n3023), .ZN(n2806) );
  NAND2_X4 U3409 ( .A1(n3150), .A2(n1655), .ZN(n3151) );
  NAND2_X4 U3410 ( .A1(n3236), .A2(n3235), .ZN(n3431) );
  OAI21_X2 U3411 ( .B1(n4218), .B2(n4217), .A(n4216), .ZN(n4219) );
  NAND2_X4 U3412 ( .A1(n3137), .A2(n3136), .ZN(n3138) );
  NAND2_X4 U3413 ( .A1(n3272), .A2(n3271), .ZN(n3341) );
  NAND2_X4 U3414 ( .A1(n3237), .A2(n3153), .ZN(net329445) );
  NAND3_X2 U3415 ( .A1(n1695), .A2(n2889), .A3(n3023), .ZN(n2890) );
  NAND3_X4 U3416 ( .A1(n1702), .A2(n2666), .A3(n2571), .ZN(n2773) );
  NAND2_X2 U3417 ( .A1(n4189), .A2(n1952), .ZN(n1834) );
  NAND2_X4 U3418 ( .A1(n1832), .A2(n4461), .ZN(n1835) );
  NAND2_X4 U3419 ( .A1(n1834), .A2(n1835), .ZN(n1951) );
  INV_X8 U3421 ( .A(n1951), .ZN(n4305) );
  NOR2_X4 U3422 ( .A1(n2474), .A2(n2475), .ZN(n2479) );
  NAND2_X2 U3424 ( .A1(n2287), .A2(net330834), .ZN(n2288) );
  NAND2_X4 U3425 ( .A1(n1625), .A2(n2665), .ZN(n2666) );
  NAND2_X4 U3426 ( .A1(n1837), .A2(n1838), .ZN(n1840) );
  NAND2_X4 U3427 ( .A1(n1839), .A2(n1840), .ZN(n3059) );
  INV_X4 U3428 ( .A(n3058), .ZN(n1837) );
  INV_X1 U3429 ( .A(n3116), .ZN(n1838) );
  INV_X8 U3430 ( .A(n3059), .ZN(n3112) );
  NAND2_X4 U3431 ( .A1(n1914), .A2(n1915), .ZN(n3172) );
  NAND2_X2 U3432 ( .A1(net329043), .A2(n4427), .ZN(n1842) );
  NAND2_X4 U3433 ( .A1(n1841), .A2(n1842), .ZN(n3677) );
  NAND2_X4 U3434 ( .A1(n3902), .A2(n3800), .ZN(net328607) );
  XNOR2_X2 U3435 ( .A(n3972), .B(n3976), .ZN(n3902) );
  NAND2_X4 U3436 ( .A1(n2932), .A2(n2933), .ZN(n3120) );
  INV_X2 U3437 ( .A(n3449), .ZN(n3450) );
  NAND2_X2 U3438 ( .A1(n2650), .A2(n2457), .ZN(n1986) );
  INV_X4 U3439 ( .A(n2457), .ZN(n1985) );
  NAND2_X4 U3440 ( .A1(n2430), .A2(n2531), .ZN(n2389) );
  NAND2_X4 U3441 ( .A1(n2957), .A2(n1186), .ZN(n2630) );
  NAND3_X4 U3442 ( .A1(n1830), .A2(n3331), .A3(n3332), .ZN(n3231) );
  INV_X2 U3443 ( .A(n4027), .ZN(n4119) );
  NAND2_X2 U3444 ( .A1(a[1]), .A2(n2104), .ZN(net331086) );
  INV_X8 U3445 ( .A(n3116), .ZN(n3118) );
  NAND2_X4 U3446 ( .A1(n2934), .A2(n3255), .ZN(n2937) );
  NAND2_X4 U3447 ( .A1(n1723), .A2(net328338), .ZN(n4263) );
  NAND2_X4 U3448 ( .A1(n2950), .A2(n2949), .ZN(net329598) );
  NAND2_X4 U3449 ( .A1(n1967), .A2(n1637), .ZN(n1969) );
  NAND2_X4 U3450 ( .A1(n3730), .A2(n3731), .ZN(n3958) );
  NAND2_X2 U3451 ( .A1(n2464), .A2(n2463), .ZN(n1845) );
  NAND2_X4 U3452 ( .A1(n1843), .A2(n1844), .ZN(n1846) );
  NAND2_X4 U3453 ( .A1(n1845), .A2(n1846), .ZN(n2632) );
  OAI211_X1 U3454 ( .C1(n2651), .C2(n2549), .A(n1756), .B(n2545), .ZN(n2464)
         );
  INV_X8 U3455 ( .A(n2543), .ZN(n2544) );
  AOI21_X4 U3456 ( .B1(n1259), .B2(n2014), .A(n3417), .ZN(n3418) );
  INV_X2 U3457 ( .A(n2752), .ZN(n1980) );
  OAI21_X4 U3458 ( .B1(n1927), .B2(n1418), .A(n4435), .ZN(n3567) );
  NAND2_X2 U3460 ( .A1(net333621), .A2(net332364), .ZN(n2758) );
  NAND2_X2 U3461 ( .A1(a[5]), .A2(net331137), .ZN(n1847) );
  INV_X4 U3463 ( .A(net331137), .ZN(net332987) );
  INV_X4 U3464 ( .A(a[5]), .ZN(net332988) );
  NAND2_X2 U3466 ( .A1(net331125), .A2(net331124), .ZN(net330990) );
  NAND2_X4 U3467 ( .A1(n3933), .A2(n1627), .ZN(n4034) );
  NAND2_X2 U3468 ( .A1(net331083), .A2(n2129), .ZN(n2131) );
  NAND2_X4 U3469 ( .A1(n2494), .A2(n2493), .ZN(n2706) );
  NAND2_X2 U3470 ( .A1(n4431), .A2(n3669), .ZN(n2991) );
  INV_X4 U3471 ( .A(n1940), .ZN(n1849) );
  NAND2_X1 U3473 ( .A1(n2745), .A2(n1709), .ZN(n2709) );
  INV_X8 U3474 ( .A(n2564), .ZN(n1862) );
  NAND2_X4 U3475 ( .A1(n3099), .A2(n3100), .ZN(n1850) );
  NAND2_X2 U3477 ( .A1(n3659), .A2(n3660), .ZN(n1855) );
  NAND2_X4 U3478 ( .A1(n1853), .A2(n1854), .ZN(n1856) );
  NAND2_X4 U3479 ( .A1(n1855), .A2(n1856), .ZN(n3662) );
  INV_X4 U3480 ( .A(n3660), .ZN(n1853) );
  INV_X2 U3481 ( .A(n3659), .ZN(n1854) );
  NAND2_X2 U3482 ( .A1(n3678), .A2(n1857), .ZN(n1858) );
  NAND2_X2 U3483 ( .A1(n1858), .A2(n1735), .ZN(n3602) );
  INV_X2 U3484 ( .A(n3760), .ZN(n1857) );
  NAND2_X2 U3485 ( .A1(net328268), .A2(n4245), .ZN(net328533) );
  INV_X16 U3486 ( .A(control[1]), .ZN(net331251) );
  NAND2_X2 U3487 ( .A1(n4386), .A2(n3158), .ZN(n1896) );
  XNOR2_X2 U3488 ( .A(net329545), .B(n3281), .ZN(n3425) );
  NAND2_X4 U3489 ( .A1(n4292), .A2(n4293), .ZN(n4355) );
  NOR2_X4 U3490 ( .A1(n4188), .A2(net328338), .ZN(n1860) );
  NAND2_X4 U3491 ( .A1(n3881), .A2(n3882), .ZN(n3978) );
  NAND2_X4 U3492 ( .A1(n3809), .A2(n3854), .ZN(n3950) );
  NAND2_X4 U3493 ( .A1(n3549), .A2(n3548), .ZN(n3625) );
  INV_X2 U3494 ( .A(n3550), .ZN(n3548) );
  NAND2_X4 U3495 ( .A1(n2549), .A2(n2651), .ZN(n2548) );
  NAND2_X4 U3496 ( .A1(n4097), .A2(n4105), .ZN(net332287) );
  INV_X1 U3498 ( .A(n3963), .ZN(n3725) );
  NAND2_X1 U3499 ( .A1(n2129), .A2(net331204), .ZN(n2062) );
  OAI21_X2 U3500 ( .B1(n2630), .B2(n2831), .A(n1286), .ZN(n2717) );
  NOR2_X4 U3501 ( .A1(n2108), .A2(n2109), .ZN(n2132) );
  NOR2_X4 U3502 ( .A1(n2051), .A2(n1333), .ZN(n2020) );
  NAND2_X1 U3504 ( .A1(n3031), .A2(n2841), .ZN(n2846) );
  NAND2_X4 U3506 ( .A1(n1205), .A2(n2179), .ZN(n2156) );
  NAND3_X2 U3507 ( .A1(net331092), .A2(n2104), .A3(n1345), .ZN(n2179) );
  NAND2_X2 U3508 ( .A1(n2258), .A2(n2257), .ZN(n1868) );
  NAND2_X4 U3509 ( .A1(n1866), .A2(n1867), .ZN(n1869) );
  NAND2_X4 U3510 ( .A1(n1868), .A2(n1869), .ZN(n2261) );
  INV_X4 U3511 ( .A(n2258), .ZN(n1866) );
  INV_X4 U3512 ( .A(n2257), .ZN(n1867) );
  NAND2_X2 U3513 ( .A1(n2137), .A2(n1650), .ZN(n1872) );
  NAND2_X4 U3514 ( .A1(n1870), .A2(n1871), .ZN(n1873) );
  NAND2_X4 U3515 ( .A1(n1872), .A2(n1873), .ZN(net330822) );
  INV_X4 U3516 ( .A(n2137), .ZN(n1870) );
  INV_X4 U3517 ( .A(n1650), .ZN(n1871) );
  NAND2_X4 U3518 ( .A1(n1624), .A2(n2203), .ZN(n1878) );
  NAND2_X4 U3519 ( .A1(n1878), .A2(n1877), .ZN(n2343) );
  NAND2_X1 U3520 ( .A1(n2321), .A2(n2320), .ZN(n2257) );
  NAND2_X2 U3521 ( .A1(n2752), .A2(n4493), .ZN(n2707) );
  AOI21_X2 U3523 ( .B1(n4261), .B2(n4360), .A(n4260), .ZN(net328183) );
  NAND2_X4 U3524 ( .A1(net328177), .A2(n4259), .ZN(n4360) );
  NAND2_X4 U3525 ( .A1(n1902), .A2(net332690), .ZN(n1904) );
  NOR2_X4 U3526 ( .A1(n3515), .A2(n1836), .ZN(n3422) );
  NAND2_X1 U3527 ( .A1(n2324), .A2(n2325), .ZN(n2263) );
  NOR2_X2 U3528 ( .A1(n3164), .A2(n2024), .ZN(n3095) );
  INV_X8 U3529 ( .A(n2156), .ZN(n2157) );
  XNOR2_X1 U3530 ( .A(n3569), .B(n1725), .ZN(product_out[22]) );
  INV_X8 U3531 ( .A(n2370), .ZN(n2375) );
  NAND2_X1 U3533 ( .A1(n3350), .A2(n3354), .ZN(n3444) );
  NAND2_X4 U3534 ( .A1(n4465), .A2(n2723), .ZN(n2734) );
  NOR2_X4 U3535 ( .A1(net331359), .A2(net331138), .ZN(n2095) );
  BUF_X32 U3536 ( .A(n2516), .Z(n1880) );
  INV_X4 U3537 ( .A(n2658), .ZN(n2460) );
  NAND2_X4 U3538 ( .A1(net328142), .A2(n4136), .ZN(net328172) );
  OAI211_X4 U3539 ( .C1(n2303), .C2(n2302), .A(n2300), .B(n2301), .ZN(n2305)
         );
  OAI21_X2 U3540 ( .B1(n3774), .B2(n3769), .A(n3775), .ZN(n3797) );
  NAND2_X2 U3541 ( .A1(n4086), .A2(n4082), .ZN(n4015) );
  NAND3_X2 U3542 ( .A1(n3124), .A2(n2932), .A3(n2933), .ZN(n2858) );
  INV_X1 U3543 ( .A(n3545), .ZN(n3543) );
  NAND2_X4 U3544 ( .A1(n3546), .A2(n3627), .ZN(n3628) );
  INV_X4 U3545 ( .A(n2305), .ZN(n1890) );
  NAND2_X2 U3546 ( .A1(net332668), .A2(n1201), .ZN(n3033) );
  INV_X4 U3547 ( .A(n2777), .ZN(n2778) );
  NAND2_X2 U3548 ( .A1(n1638), .A2(n2793), .ZN(n1968) );
  NOR2_X4 U3549 ( .A1(n4191), .A2(net328027), .ZN(net332747) );
  NAND2_X4 U3550 ( .A1(n2227), .A2(n1420), .ZN(n2230) );
  NAND2_X2 U3551 ( .A1(n2315), .A2(n2314), .ZN(n1884) );
  NAND2_X4 U3552 ( .A1(n1882), .A2(n1883), .ZN(n1885) );
  NAND2_X4 U3553 ( .A1(n1885), .A2(n1884), .ZN(n2317) );
  XNOR2_X2 U3554 ( .A(n2231), .B(net330910), .ZN(n1886) );
  NAND2_X2 U3555 ( .A1(n2237), .A2(n2238), .ZN(n1888) );
  NAND2_X4 U3556 ( .A1(n1887), .A2(n2236), .ZN(n1889) );
  NAND2_X4 U3557 ( .A1(n1888), .A2(n1889), .ZN(n2240) );
  INV_X4 U3558 ( .A(n2238), .ZN(n1887) );
  INV_X4 U3559 ( .A(n3443), .ZN(n3448) );
  NAND2_X4 U3560 ( .A1(n2229), .A2(n1960), .ZN(n2365) );
  NAND2_X4 U3561 ( .A1(n2766), .A2(n2769), .ZN(n2579) );
  INV_X2 U3562 ( .A(n1417), .ZN(n2518) );
  NAND2_X4 U3563 ( .A1(n3368), .A2(n3369), .ZN(n3371) );
  NAND2_X2 U3564 ( .A1(n3770), .A2(n3772), .ZN(n3796) );
  INV_X4 U3565 ( .A(n3702), .ZN(n3701) );
  NAND2_X2 U3566 ( .A1(n2304), .A2(n2305), .ZN(n1892) );
  NAND2_X4 U3567 ( .A1(n1890), .A2(n1891), .ZN(n1893) );
  NAND2_X4 U3568 ( .A1(n1892), .A2(n1893), .ZN(n2358) );
  INV_X4 U3569 ( .A(n2304), .ZN(n1891) );
  NAND2_X4 U3570 ( .A1(n1894), .A2(n1895), .ZN(n1897) );
  NAND2_X4 U3572 ( .A1(n1898), .A2(n1899), .ZN(n1901) );
  NAND2_X4 U3573 ( .A1(n1904), .A2(n1903), .ZN(n2174) );
  NAND2_X2 U3574 ( .A1(a[6]), .A2(net331357), .ZN(n2164) );
  NAND2_X1 U3575 ( .A1(n4322), .A2(n4321), .ZN(n4324) );
  NAND2_X2 U3576 ( .A1(n2500), .A2(n2499), .ZN(n2628) );
  NAND2_X4 U3577 ( .A1(n2860), .A2(n2859), .ZN(n2861) );
  NOR2_X4 U3578 ( .A1(n2931), .A2(n3121), .ZN(n2860) );
  OAI21_X4 U3579 ( .B1(n3906), .B2(n3905), .A(net328601), .ZN(n3907) );
  NAND2_X4 U3580 ( .A1(n2819), .A2(n3177), .ZN(n2901) );
  INV_X1 U3581 ( .A(n1954), .ZN(n4024) );
  NAND2_X2 U3582 ( .A1(n2837), .A2(n2698), .ZN(n2596) );
  NAND3_X2 U3583 ( .A1(n1192), .A2(n1246), .A3(n1355), .ZN(n3398) );
  NAND2_X2 U3585 ( .A1(n1259), .A2(n3387), .ZN(n1910) );
  NAND2_X4 U3586 ( .A1(n1908), .A2(n1909), .ZN(n1911) );
  NAND2_X4 U3587 ( .A1(n1910), .A2(n1911), .ZN(n3390) );
  INV_X2 U3589 ( .A(n1134), .ZN(n4260) );
  NAND2_X2 U3590 ( .A1(n4190), .A2(n1951), .ZN(n4363) );
  NAND2_X2 U3591 ( .A1(net329992), .A2(n2637), .ZN(n2550) );
  OAI21_X4 U3592 ( .B1(net328483), .B2(net328484), .A(net328485), .ZN(n4075)
         );
  XNOR2_X2 U3593 ( .A(n3972), .B(n3801), .ZN(n3802) );
  INV_X4 U3594 ( .A(n3429), .ZN(n3609) );
  NAND2_X2 U3595 ( .A1(n2018), .A2(n3171), .ZN(n1914) );
  INV_X1 U3597 ( .A(net329549), .ZN(net329547) );
  NAND2_X1 U3598 ( .A1(n3181), .A2(n3178), .ZN(n2905) );
  INV_X2 U3599 ( .A(n3178), .ZN(n3176) );
  INV_X4 U3600 ( .A(n2732), .ZN(n1916) );
  INV_X8 U3601 ( .A(n1916), .ZN(n1917) );
  OAI211_X2 U3602 ( .C1(net329860), .C2(net333802), .A(n3035), .B(n3034), .ZN(
        n3036) );
  INV_X1 U3603 ( .A(n3262), .ZN(n3260) );
  NAND3_X2 U3604 ( .A1(n4041), .A2(n4042), .A3(n4043), .ZN(n1918) );
  INV_X4 U3605 ( .A(n4177), .ZN(n4178) );
  INV_X4 U3606 ( .A(n2866), .ZN(n2864) );
  NAND2_X2 U3607 ( .A1(n3555), .A2(n3554), .ZN(n3687) );
  OAI21_X4 U3608 ( .B1(n2659), .B2(n2658), .A(n2657), .ZN(n2662) );
  NAND2_X1 U3609 ( .A1(n4296), .A2(n4094), .ZN(n3918) );
  NAND2_X2 U3610 ( .A1(net331520), .A2(net328409), .ZN(n1919) );
  NAND2_X4 U3611 ( .A1(net332585), .A2(net332586), .ZN(n1920) );
  NAND2_X4 U3612 ( .A1(n1920), .A2(n1919), .ZN(net328408) );
  INV_X4 U3613 ( .A(net331520), .ZN(net332585) );
  INV_X4 U3614 ( .A(net328409), .ZN(net332586) );
  NAND3_X2 U3615 ( .A1(n3193), .A2(n1680), .A3(control[1]), .ZN(n2989) );
  NAND2_X4 U3616 ( .A1(n3475), .A2(n3474), .ZN(n3680) );
  NAND2_X2 U3617 ( .A1(n2021), .A2(n2482), .ZN(n1923) );
  NAND2_X4 U3618 ( .A1(n1921), .A2(n1922), .ZN(n1924) );
  NAND2_X4 U3619 ( .A1(n1923), .A2(n1924), .ZN(n2543) );
  INV_X2 U3620 ( .A(n2021), .ZN(n1922) );
  NAND2_X4 U3621 ( .A1(n2543), .A2(n2483), .ZN(n2631) );
  INV_X8 U3622 ( .A(n3678), .ZN(n1955) );
  INV_X4 U3623 ( .A(n2499), .ZN(n2497) );
  INV_X2 U3624 ( .A(n3710), .ZN(n3704) );
  INV_X2 U3625 ( .A(n1657), .ZN(n3503) );
  NAND2_X2 U3626 ( .A1(net330037), .A2(net330038), .ZN(n2800) );
  XNOR2_X2 U3627 ( .A(n4367), .B(net328019), .ZN(n4368) );
  INV_X8 U3628 ( .A(n3507), .ZN(n3586) );
  NAND2_X4 U3629 ( .A1(n1928), .A2(n1701), .ZN(n1930) );
  NAND2_X4 U3630 ( .A1(n1929), .A2(n1930), .ZN(net330738) );
  INV_X32 U3631 ( .A(control[1]), .ZN(net331200) );
  INV_X32 U3632 ( .A(control[1]), .ZN(net331192) );
  NAND2_X4 U3634 ( .A1(n1634), .A2(n2180), .ZN(n2082) );
  NAND3_X2 U3635 ( .A1(n2537), .A2(n2536), .A3(n2540), .ZN(n2487) );
  NAND3_X2 U3636 ( .A1(n2963), .A2(n2831), .A3(n1286), .ZN(n2965) );
  AOI21_X4 U3637 ( .B1(n2181), .B2(net330819), .A(net330918), .ZN(n2182) );
  NAND2_X1 U3638 ( .A1(n2069), .A2(n1348), .ZN(net331228) );
  NAND2_X4 U3639 ( .A1(n2160), .A2(n2159), .ZN(n2218) );
  NAND2_X4 U3640 ( .A1(n4271), .A2(n4267), .ZN(n4186) );
  NAND2_X4 U3641 ( .A1(n1932), .A2(n2596), .ZN(n1934) );
  NAND2_X4 U3642 ( .A1(n1933), .A2(n1934), .ZN(n2600) );
  INV_X4 U3643 ( .A(n2598), .ZN(n1932) );
  NAND2_X4 U3644 ( .A1(net331025), .A2(n2157), .ZN(n1936) );
  NAND2_X2 U3645 ( .A1(net329407), .A2(net329398), .ZN(n1937) );
  NAND2_X4 U3646 ( .A1(net332462), .A2(net332463), .ZN(n1938) );
  NAND2_X4 U3647 ( .A1(n1938), .A2(n1937), .ZN(n3379) );
  INV_X4 U3648 ( .A(net329407), .ZN(net332462) );
  INV_X2 U3649 ( .A(net329398), .ZN(net332463) );
  NAND2_X4 U3650 ( .A1(n4067), .A2(n4068), .ZN(n4071) );
  NAND2_X4 U3651 ( .A1(n3335), .A2(n3157), .ZN(n3227) );
  NAND2_X4 U3652 ( .A1(n2561), .A2(n2222), .ZN(n2225) );
  NAND2_X2 U3653 ( .A1(n2496), .A2(n2495), .ZN(n1943) );
  NAND2_X4 U3654 ( .A1(n1941), .A2(n1942), .ZN(n1944) );
  NAND2_X4 U3655 ( .A1(n1943), .A2(n1944), .ZN(n2499) );
  INV_X4 U3656 ( .A(n2496), .ZN(n1941) );
  INV_X4 U3657 ( .A(n2495), .ZN(n1942) );
  INV_X8 U3658 ( .A(n2167), .ZN(n2096) );
  NAND2_X4 U3659 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  INV_X4 U3660 ( .A(n3938), .ZN(n3576) );
  NAND2_X4 U3661 ( .A1(n3585), .A2(n3411), .ZN(n3412) );
  NAND4_X4 U3662 ( .A1(n1794), .A2(n1114), .A3(n3408), .A4(n2025), .ZN(n3585)
         );
  NAND2_X4 U3663 ( .A1(n4184), .A2(n4185), .ZN(n4267) );
  NAND2_X4 U3664 ( .A1(n1140), .A2(n3944), .ZN(n4245) );
  NAND2_X4 U3665 ( .A1(n3332), .A2(n3103), .ZN(n3101) );
  NAND2_X4 U3666 ( .A1(n1826), .A2(n3405), .ZN(n3587) );
  NAND2_X1 U3668 ( .A1(n4360), .A2(n4484), .ZN(n4362) );
  INV_X2 U3669 ( .A(n3337), .ZN(n3234) );
  NAND2_X4 U3670 ( .A1(n3225), .A2(n3226), .ZN(n3337) );
  NAND2_X4 U3671 ( .A1(n1948), .A2(n2978), .ZN(n1950) );
  AND2_X2 U3672 ( .A1(n4262), .A2(n4263), .ZN(n1952) );
  INV_X2 U3673 ( .A(n3912), .ZN(n3910) );
  INV_X4 U3674 ( .A(n3854), .ZN(n3856) );
  NAND2_X4 U3675 ( .A1(n2544), .A2(n2545), .ZN(n1953) );
  NAND2_X4 U3676 ( .A1(n2071), .A2(n2070), .ZN(n2060) );
  INV_X4 U3677 ( .A(n1740), .ZN(n4011) );
  NAND2_X2 U3678 ( .A1(n2412), .A2(n2411), .ZN(n2629) );
  NAND3_X4 U3679 ( .A1(n4072), .A2(net328485), .A3(net328491), .ZN(n4146) );
  NAND2_X2 U3680 ( .A1(n3562), .A2(n3561), .ZN(n1994) );
  NAND2_X2 U3681 ( .A1(n2265), .A2(n2264), .ZN(n2241) );
  NAND2_X2 U3682 ( .A1(n3813), .A2(n1366), .ZN(n3719) );
  NAND2_X4 U3684 ( .A1(n2044), .A2(n1327), .ZN(n2206) );
  OAI21_X1 U3685 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(n4334) );
  INV_X1 U3686 ( .A(n3637), .ZN(n3458) );
  NAND3_X1 U3687 ( .A1(n4458), .A2(n2647), .A3(n2702), .ZN(n3008) );
  NAND2_X4 U3688 ( .A1(n2346), .A2(n2746), .ZN(n2314) );
  NAND2_X4 U3689 ( .A1(n3853), .A2(n3852), .ZN(n3766) );
  XNOR2_X2 U3690 ( .A(n3472), .B(n1959), .ZN(n1958) );
  NAND2_X4 U3692 ( .A1(n2947), .A2(n2948), .ZN(net329876) );
  NAND3_X1 U3693 ( .A1(n2503), .A2(n2629), .A3(n1338), .ZN(n2505) );
  INV_X2 U3694 ( .A(n4245), .ZN(n3945) );
  NAND2_X1 U3695 ( .A1(n4118), .A2(n4245), .ZN(n4126) );
  NAND2_X1 U3696 ( .A1(n4119), .A2(n4245), .ZN(n4127) );
  NAND3_X2 U3697 ( .A1(n3604), .A2(n3612), .A3(n3605), .ZN(n3558) );
  NAND2_X4 U3698 ( .A1(n1119), .A2(n3521), .ZN(n3471) );
  NAND2_X2 U3699 ( .A1(n4364), .A2(n1686), .ZN(n4367) );
  NAND2_X1 U3700 ( .A1(net330738), .A2(n1608), .ZN(n2303) );
  NAND2_X4 U3702 ( .A1(n1343), .A2(n3083), .ZN(n3186) );
  NAND2_X4 U3703 ( .A1(n3896), .A2(n2023), .ZN(net328865) );
  NOR2_X4 U3704 ( .A1(n3599), .A2(n1331), .ZN(n1963) );
  NAND2_X2 U3705 ( .A1(net333078), .A2(n2591), .ZN(n1965) );
  NAND2_X4 U3706 ( .A1(n1964), .A2(net332292), .ZN(n1966) );
  NAND2_X4 U3707 ( .A1(n1965), .A2(n1966), .ZN(net330456) );
  NAND2_X4 U3708 ( .A1(n1968), .A2(n1969), .ZN(n2797) );
  INV_X4 U3709 ( .A(n2793), .ZN(n1967) );
  NAND2_X1 U3710 ( .A1(a[30]), .A2(net333222), .ZN(n4312) );
  NAND2_X1 U3711 ( .A1(a[29]), .A2(n4488), .ZN(n4281) );
  NAND3_X2 U3712 ( .A1(a[4]), .A2(n4488), .A3(n2135), .ZN(n2168) );
  NAND2_X2 U3713 ( .A1(a[6]), .A2(net331357), .ZN(n2281) );
  INV_X2 U3714 ( .A(n2847), .ZN(n2761) );
  NAND2_X4 U3715 ( .A1(n1691), .A2(n2391), .ZN(n2420) );
  NAND3_X2 U3716 ( .A1(net330652), .A2(net330653), .A3(net330654), .ZN(
        net330651) );
  NAND2_X4 U3717 ( .A1(n3900), .A2(n3899), .ZN(net328597) );
  NAND3_X4 U3718 ( .A1(n3133), .A2(n3134), .A3(n3135), .ZN(n3137) );
  NAND2_X2 U3719 ( .A1(n3132), .A2(n3131), .ZN(n3134) );
  NAND2_X4 U3720 ( .A1(n2718), .A2(n2719), .ZN(n2736) );
  INV_X1 U3721 ( .A(net328025), .ZN(net328023) );
  NAND2_X4 U3722 ( .A1(n2633), .A2(n1132), .ZN(n2643) );
  NAND2_X4 U3723 ( .A1(n2266), .A2(n1626), .ZN(n2425) );
  NAND2_X4 U3724 ( .A1(net330983), .A2(net331029), .ZN(n2184) );
  NAND2_X4 U3725 ( .A1(net328615), .A2(net328601), .ZN(net328599) );
  NAND2_X4 U3726 ( .A1(n3904), .A2(n3802), .ZN(net328601) );
  OAI21_X4 U3727 ( .B1(net332050), .B2(net329453), .A(net333532), .ZN(n3241)
         );
  NAND2_X4 U3728 ( .A1(a[5]), .A2(net331349), .ZN(n2128) );
  NAND2_X4 U3729 ( .A1(n1973), .A2(n1972), .ZN(n1975) );
  NAND2_X4 U3730 ( .A1(n1975), .A2(n1974), .ZN(n4069) );
  INV_X4 U3731 ( .A(n4066), .ZN(n1972) );
  INV_X4 U3732 ( .A(n4065), .ZN(n1973) );
  INV_X4 U3733 ( .A(n4069), .ZN(n4067) );
  NAND3_X1 U3734 ( .A1(a[27]), .A2(n4052), .A3(net331351), .ZN(n4160) );
  NAND2_X1 U3735 ( .A1(a[26]), .A2(net331351), .ZN(n3980) );
  NAND2_X4 U3736 ( .A1(a[12]), .A2(net331351), .ZN(n2668) );
  INV_X4 U3737 ( .A(n3729), .ZN(n3731) );
  NAND2_X4 U3738 ( .A1(n3846), .A2(n1280), .ZN(n4093) );
  OAI21_X4 U3739 ( .B1(n2635), .B2(n2634), .A(n1953), .ZN(n2636) );
  NAND2_X2 U3740 ( .A1(n4176), .A2(n1918), .ZN(n4179) );
  INV_X1 U3741 ( .A(n3642), .ZN(n3644) );
  NAND2_X4 U3742 ( .A1(n3464), .A2(n3531), .ZN(n3532) );
  NOR2_X2 U3743 ( .A1(n2273), .A2(n2307), .ZN(n2274) );
  NOR2_X2 U3744 ( .A1(n2377), .A2(n2126), .ZN(n2373) );
  NAND2_X2 U3745 ( .A1(n3553), .A2(n1409), .ZN(n1977) );
  NAND2_X4 U3746 ( .A1(n1976), .A2(net328869), .ZN(n1978) );
  NAND3_X2 U3747 ( .A1(n1643), .A2(net329992), .A3(net333659), .ZN(n2691) );
  NAND2_X4 U3748 ( .A1(n3696), .A2(n3697), .ZN(n3698) );
  NAND2_X4 U3749 ( .A1(n3345), .A2(n3344), .ZN(n3349) );
  NAND2_X4 U3750 ( .A1(n3371), .A2(n3449), .ZN(n3441) );
  NAND2_X4 U3752 ( .A1(n2073), .A2(n2072), .ZN(n2059) );
  NAND2_X4 U3753 ( .A1(n1981), .A2(n2751), .ZN(n3020) );
  INV_X8 U3754 ( .A(n2833), .ZN(n2976) );
  INV_X8 U3755 ( .A(n3138), .ZN(n3249) );
  INV_X8 U3756 ( .A(n2922), .ZN(n2923) );
  NAND2_X4 U3757 ( .A1(net328470), .A2(n4082), .ZN(n4083) );
  INV_X8 U3758 ( .A(n1982), .ZN(n1983) );
  AOI22_X1 U3759 ( .A1(n2624), .A2(n2623), .B1(n2622), .B2(n2621), .ZN(n1984)
         );
  NAND2_X1 U3760 ( .A1(net328035), .A2(n1716), .ZN(net328031) );
  NAND2_X1 U3761 ( .A1(net331362), .A2(n4365), .ZN(n3665) );
  INV_X4 U3763 ( .A(n3003), .ZN(n2967) );
  NAND2_X4 U3764 ( .A1(n2753), .A2(n3010), .ZN(n2886) );
  NAND3_X2 U3766 ( .A1(n2295), .A2(n2294), .A3(n2293), .ZN(n2437) );
  NAND2_X2 U3767 ( .A1(a[1]), .A2(n2032), .ZN(net331245) );
  INV_X4 U3768 ( .A(net331245), .ZN(net331154) );
  NAND2_X4 U3769 ( .A1(n1985), .A2(n1651), .ZN(n1987) );
  NAND2_X4 U3770 ( .A1(n1986), .A2(n1987), .ZN(n2549) );
  NAND2_X4 U3771 ( .A1(n2549), .A2(n2651), .ZN(net329992) );
  NAND2_X1 U3772 ( .A1(n2958), .A2(n2957), .ZN(n2834) );
  INV_X4 U3773 ( .A(n2958), .ZN(n2960) );
  NAND2_X4 U3774 ( .A1(n1640), .A2(a[5]), .ZN(n2134) );
  NAND2_X2 U3775 ( .A1(n1388), .A2(net328872), .ZN(n3901) );
  NAND2_X4 U3776 ( .A1(n3720), .A2(n3721), .ZN(n3962) );
  NAND2_X4 U3777 ( .A1(n4180), .A2(n4177), .ZN(n4065) );
  NAND2_X4 U3778 ( .A1(n3233), .A2(n2028), .ZN(n3283) );
  NAND2_X4 U3779 ( .A1(net328388), .A2(n1397), .ZN(n4079) );
  NAND2_X4 U3780 ( .A1(n2832), .A2(n2964), .ZN(n2833) );
  INV_X1 U3781 ( .A(n2337), .ZN(n2335) );
  NAND3_X1 U3782 ( .A1(n2117), .A2(n2116), .A3(net331032), .ZN(n2187) );
  NAND3_X2 U3783 ( .A1(net331119), .A2(n1221), .A3(n2113), .ZN(n2117) );
  NAND3_X1 U3784 ( .A1(n3686), .A2(n3518), .A3(n3416), .ZN(n3380) );
  AOI21_X4 U3785 ( .B1(n4179), .B2(n4180), .A(n4178), .ZN(n4285) );
  NAND2_X4 U3786 ( .A1(control[0]), .A2(net329919), .ZN(net328712) );
  AOI22_X4 U3787 ( .A1(n1786), .A2(n3851), .B1(n3850), .B2(n1396), .ZN(n3919)
         );
  NAND2_X4 U3788 ( .A1(n1989), .A2(n1990), .ZN(n1991) );
  INV_X4 U3790 ( .A(n2170), .ZN(n1989) );
  INV_X4 U3791 ( .A(n2577), .ZN(n1990) );
  NAND2_X4 U3792 ( .A1(n1992), .A2(n1993), .ZN(n1995) );
  NAND2_X4 U3793 ( .A1(n1995), .A2(n1994), .ZN(n3599) );
  INV_X4 U3794 ( .A(n3561), .ZN(n1993) );
  NAND2_X2 U3795 ( .A1(n2878), .A2(net333336), .ZN(n1997) );
  NAND2_X4 U3796 ( .A1(n1996), .A2(net332088), .ZN(n1998) );
  NAND2_X4 U3797 ( .A1(n2267), .A2(n2421), .ZN(n2315) );
  NAND2_X2 U3798 ( .A1(n1131), .A2(n3767), .ZN(net328984) );
  INV_X4 U3799 ( .A(n3606), .ZN(n3607) );
  NAND2_X1 U3800 ( .A1(net328855), .A2(net328856), .ZN(n3859) );
  NAND2_X4 U3801 ( .A1(n3639), .A2(n3640), .ZN(n3642) );
  NAND2_X4 U3802 ( .A1(n3641), .A2(n3642), .ZN(n3696) );
  NAND2_X4 U3803 ( .A1(n3296), .A2(n3297), .ZN(n1999) );
  NAND2_X2 U3804 ( .A1(n1695), .A2(n2888), .ZN(n2000) );
  NAND2_X4 U3805 ( .A1(n2259), .A2(n2260), .ZN(n2324) );
  NAND2_X2 U3806 ( .A1(n1303), .A2(n2416), .ZN(n2001) );
  OAI21_X2 U3807 ( .B1(n2533), .B2(n2532), .A(n4493), .ZN(n2534) );
  NOR3_X2 U3808 ( .A1(n3738), .A2(n3960), .A3(net331295), .ZN(n3740) );
  INV_X8 U3809 ( .A(n3240), .ZN(n3345) );
  NOR2_X2 U3810 ( .A1(net329398), .A2(net329397), .ZN(n3384) );
  INV_X4 U3811 ( .A(n2536), .ZN(n2539) );
  INV_X4 U3812 ( .A(n3318), .ZN(n3193) );
  OAI21_X1 U3813 ( .B1(n4356), .B2(net328051), .A(n4481), .ZN(n4357) );
  NAND2_X4 U3815 ( .A1(n2004), .A2(n2005), .ZN(n2840) );
  NAND2_X4 U3816 ( .A1(net332007), .A2(net332006), .ZN(n2006) );
  NAND2_X4 U3817 ( .A1(n2006), .A2(net329988), .ZN(net330131) );
  INV_X4 U3818 ( .A(net330239), .ZN(net332006) );
  INV_X4 U3819 ( .A(n1308), .ZN(net332007) );
  INV_X1 U3820 ( .A(net330330), .ZN(net330239) );
  NAND2_X2 U3821 ( .A1(n2602), .A2(n2601), .ZN(n2009) );
  NAND2_X4 U3822 ( .A1(n2007), .A2(n2008), .ZN(n2010) );
  NAND2_X4 U3823 ( .A1(n2010), .A2(n2009), .ZN(n2604) );
  INV_X4 U3824 ( .A(n2602), .ZN(n2007) );
  INV_X4 U3825 ( .A(n2601), .ZN(n2008) );
  NOR2_X4 U3826 ( .A1(n1881), .A2(n2228), .ZN(n2175) );
  NAND2_X4 U3827 ( .A1(n4072), .A2(net328491), .ZN(net328595) );
  NAND2_X4 U3828 ( .A1(n1728), .A2(n3152), .ZN(n3237) );
  NAND2_X1 U3829 ( .A1(a[31]), .A2(n1719), .ZN(n4318) );
  NAND2_X1 U3830 ( .A1(a[0]), .A2(n1719), .ZN(net329043) );
  NAND2_X1 U3831 ( .A1(a[29]), .A2(n1719), .ZN(n4159) );
  NAND2_X1 U3832 ( .A1(a[28]), .A2(n1719), .ZN(n4051) );
  NAND2_X1 U3833 ( .A1(a[27]), .A2(n1719), .ZN(n3981) );
  NAND2_X1 U3834 ( .A1(a[26]), .A2(n1719), .ZN(n3867) );
  NAND2_X1 U3835 ( .A1(a[25]), .A2(n1719), .ZN(n3778) );
  NAND2_X1 U3836 ( .A1(a[23]), .A2(n1719), .ZN(n3630) );
  NAND2_X1 U3837 ( .A1(a[22]), .A2(n1719), .ZN(n3539) );
  NAND2_X1 U3838 ( .A1(a[21]), .A2(n1719), .ZN(n3457) );
  NAND2_X1 U3839 ( .A1(a[20]), .A2(n1719), .ZN(n3365) );
  NAND2_X1 U3840 ( .A1(a[19]), .A2(n1719), .ZN(n3259) );
  NAND2_X4 U3842 ( .A1(n2188), .A2(n4438), .ZN(n2190) );
  NAND2_X4 U3843 ( .A1(n2142), .A2(n2143), .ZN(n2188) );
  NAND2_X1 U3844 ( .A1(n2796), .A2(n2797), .ZN(n2011) );
  XNOR2_X2 U3845 ( .A(n2063), .B(net331131), .ZN(n2065) );
  INV_X16 U3846 ( .A(n4325), .ZN(n2036) );
  INV_X8 U3847 ( .A(n2442), .ZN(n2282) );
  NAND2_X4 U3848 ( .A1(n1174), .A2(n1209), .ZN(n2080) );
  NAND2_X4 U3849 ( .A1(n3361), .A2(n3362), .ZN(n3363) );
  NAND2_X4 U3850 ( .A1(n3262), .A2(n3263), .ZN(n3361) );
  NOR2_X4 U3851 ( .A1(net328253), .A2(net331939), .ZN(n4253) );
  OR2_X2 U3852 ( .A1(n2405), .A2(n2404), .ZN(n2013) );
  NAND2_X4 U3853 ( .A1(n2403), .A2(n2013), .ZN(n2507) );
  INV_X4 U3854 ( .A(n2252), .ZN(n2250) );
  NAND2_X4 U3855 ( .A1(a[2]), .A2(net331307), .ZN(n2404) );
  INV_X4 U3856 ( .A(n2507), .ZN(n2511) );
  NAND2_X1 U3857 ( .A1(net328790), .A2(n1384), .ZN(n3860) );
  NOR2_X2 U3858 ( .A1(n3210), .A2(n1122), .ZN(n3215) );
  INV_X2 U3859 ( .A(n3510), .ZN(n2014) );
  NAND2_X4 U3860 ( .A1(n2872), .A2(n3038), .ZN(n2922) );
  NAND2_X4 U3861 ( .A1(n3197), .A2(n2025), .ZN(n3198) );
  INV_X4 U3862 ( .A(n2632), .ZN(n2634) );
  NOR2_X4 U3863 ( .A1(n3685), .A2(n3684), .ZN(n3692) );
  NAND2_X2 U3864 ( .A1(n1668), .A2(n3005), .ZN(n2811) );
  INV_X1 U3866 ( .A(n2623), .ZN(n2015) );
  NAND3_X2 U3867 ( .A1(net329455), .A2(net329456), .A3(net329824), .ZN(
        net329737) );
  NAND2_X2 U3868 ( .A1(n3657), .A2(n3656), .ZN(n2016) );
  INV_X2 U3869 ( .A(net331895), .ZN(net331896) );
  INV_X4 U3870 ( .A(n2339), .ZN(n2516) );
  NAND2_X4 U3871 ( .A1(n2567), .A2(n2378), .ZN(n2564) );
  NAND2_X4 U3872 ( .A1(n2031), .A2(net331480), .ZN(n4089) );
  INV_X2 U3873 ( .A(net328406), .ZN(net328403) );
  INV_X2 U3874 ( .A(n3203), .ZN(n2018) );
  NAND3_X2 U3875 ( .A1(n1661), .A2(n3039), .A3(n2921), .ZN(n2926) );
  NAND2_X4 U3876 ( .A1(net329753), .A2(net333577), .ZN(n3107) );
  NAND2_X4 U3877 ( .A1(n3401), .A2(n3502), .ZN(n3938) );
  NAND2_X2 U3878 ( .A1(n1496), .A2(net328122), .ZN(net328110) );
  NOR2_X2 U3879 ( .A1(n3837), .A2(n1644), .ZN(n3838) );
  NAND2_X2 U3882 ( .A1(n2253), .A2(n2252), .ZN(n2414) );
  NAND3_X2 U3883 ( .A1(a[1]), .A2(n2192), .A3(net331323), .ZN(n2243) );
  INV_X16 U3884 ( .A(net331357), .ZN(net331353) );
  NAND2_X1 U3885 ( .A1(a[17]), .A2(n2125), .ZN(n3048) );
  NOR2_X4 U3886 ( .A1(n2675), .A2(n2674), .ZN(n2680) );
  NAND2_X1 U3887 ( .A1(n4256), .A2(n1422), .ZN(n4359) );
  OAI21_X4 U3888 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(net328855) );
  XNOR2_X1 U3889 ( .A(n1984), .B(n2730), .ZN(product_out[13]) );
  XNOR2_X1 U3890 ( .A(n1710), .B(n1185), .ZN(product_out[11]) );
  NOR3_X2 U3891 ( .A1(n4020), .A2(n4019), .A3(net331295), .ZN(n3299) );
  OAI211_X2 U3892 ( .C1(n4372), .C2(n4373), .A(n4371), .B(net331506), .ZN(
        n4374) );
  NOR3_X4 U3893 ( .A1(n1415), .A2(n4394), .A3(net330737), .ZN(n2369) );
  NOR2_X4 U3894 ( .A1(n2020), .A2(n2219), .ZN(n2101) );
  INV_X4 U3895 ( .A(n3062), .ZN(n3063) );
  NAND2_X1 U3896 ( .A1(n2667), .A2(n2766), .ZN(n2670) );
  NAND2_X4 U3897 ( .A1(n2987), .A2(n2969), .ZN(n2972) );
  NAND2_X4 U3898 ( .A1(n2894), .A2(n2893), .ZN(n2969) );
  NAND2_X4 U3899 ( .A1(n2807), .A2(n2808), .ZN(n2964) );
  INV_X8 U3900 ( .A(n4094), .ZN(n4298) );
  NOR2_X2 U3901 ( .A1(n2850), .A2(n2851), .ZN(n2774) );
  XNOR2_X1 U3902 ( .A(n2015), .B(n2624), .ZN(product_out[12]) );
  INV_X1 U3903 ( .A(net329592), .ZN(net331798) );
  OAI21_X2 U3904 ( .B1(n3530), .B2(n3529), .A(net329112), .ZN(n3552) );
  NAND2_X4 U3905 ( .A1(n3782), .A2(n3783), .ZN(n3863) );
  NAND2_X4 U3906 ( .A1(n4288), .A2(n4331), .ZN(n4343) );
  NAND2_X4 U3907 ( .A1(n1346), .A2(n3120), .ZN(n3255) );
  NAND2_X1 U3908 ( .A1(a[25]), .A2(n1164), .ZN(n3866) );
  INV_X4 U3910 ( .A(n2537), .ZN(n2538) );
  OAI21_X4 U3911 ( .B1(net330379), .B2(n2655), .A(n1643), .ZN(n2692) );
  INV_X4 U3913 ( .A(n2022), .ZN(n2023) );
  INV_X8 U3914 ( .A(n3129), .ZN(n2931) );
  NAND2_X4 U3915 ( .A1(n2609), .A2(n2608), .ZN(n2610) );
  INV_X4 U3916 ( .A(n2268), .ZN(n2270) );
  INV_X8 U3917 ( .A(n2351), .ZN(n2353) );
  NAND2_X4 U3918 ( .A1(n2828), .A2(n2628), .ZN(n2607) );
  NAND2_X4 U3919 ( .A1(n3421), .A2(n1777), .ZN(n3516) );
  NOR2_X4 U3920 ( .A1(n3508), .A2(n1684), .ZN(n3513) );
  OAI21_X2 U3921 ( .B1(n2660), .B2(n1156), .A(net333079), .ZN(n2661) );
  NAND2_X4 U3922 ( .A1(a[16]), .A2(net331349), .ZN(n3047) );
  NAND2_X4 U3924 ( .A1(n3062), .A2(n3061), .ZN(net329345) );
  NAND2_X4 U3925 ( .A1(n3832), .A2(n3833), .ZN(n4237) );
  NAND2_X4 U3926 ( .A1(n2291), .A2(n1936), .ZN(n2442) );
  NAND2_X4 U3927 ( .A1(n2291), .A2(n1936), .ZN(n2663) );
  NAND2_X4 U3928 ( .A1(n3112), .A2(n1211), .ZN(n3239) );
  NAND2_X4 U3929 ( .A1(n3112), .A2(n1211), .ZN(n3347) );
  NAND3_X2 U3930 ( .A1(n1325), .A2(b[10]), .A3(control[1]), .ZN(n2041) );
  NAND2_X4 U3931 ( .A1(n1294), .A2(control[1]), .ZN(net328030) );
  NAND4_X4 U3932 ( .A1(n1310), .A2(b[8]), .A3(control[1]), .A4(a[3]), .ZN(
        n2054) );
  NAND4_X4 U3933 ( .A1(a[3]), .A2(b[0]), .A3(control[0]), .A4(control[1]), 
        .ZN(n2055) );
  AOI21_X1 U3934 ( .B1(n3963), .B2(n4457), .A(n3960), .ZN(n3824) );
  AOI21_X4 U3935 ( .B1(n4125), .B2(n4124), .A(n4123), .ZN(n4134) );
  NAND3_X2 U3936 ( .A1(n2426), .A2(n2266), .A3(n1626), .ZN(n2267) );
  INV_X8 U3937 ( .A(n3447), .ZN(n3352) );
  NAND3_X2 U3938 ( .A1(net333079), .A2(net330024), .A3(net333315), .ZN(n3042)
         );
  NAND3_X2 U3939 ( .A1(a[7]), .A2(n2814), .A3(net331305), .ZN(n2982) );
  NAND2_X4 U3940 ( .A1(n1729), .A2(n4449), .ZN(n3765) );
  NAND2_X4 U3941 ( .A1(n1136), .A2(net331295), .ZN(n4251) );
  NAND2_X4 U3942 ( .A1(net329457), .A2(n3340), .ZN(net329399) );
  NOR2_X2 U3943 ( .A1(net333044), .A2(net328450), .ZN(n4102) );
  OAI21_X4 U3944 ( .B1(n3338), .B2(n3382), .A(n1776), .ZN(n3683) );
  XNOR2_X1 U3948 ( .A(n3797), .B(n3796), .ZN(n3798) );
  INV_X1 U3949 ( .A(n2909), .ZN(n2836) );
  NAND2_X4 U3950 ( .A1(n2918), .A2(n2780), .ZN(n2476) );
  OAI22_X1 U3951 ( .A1(n2846), .A2(n1283), .B1(n2844), .B2(n2843), .ZN(
        net330130) );
  OAI21_X4 U3952 ( .B1(n2538), .B2(n2539), .A(n2541), .ZN(n2646) );
  NAND2_X4 U3953 ( .A1(n2089), .A2(n2088), .ZN(n2141) );
  NAND2_X4 U3954 ( .A1(n3286), .A2(n3287), .ZN(n3413) );
  NAND3_X4 U3955 ( .A1(n1310), .A2(control[1]), .A3(b[8]), .ZN(n2044) );
  NAND2_X4 U3956 ( .A1(n1828), .A2(n2176), .ZN(n2177) );
  AOI22_X4 U3957 ( .A1(n4044), .A2(n4152), .B1(n4151), .B2(n4152), .ZN(n4060)
         );
  NAND2_X4 U3958 ( .A1(n1705), .A2(n3186), .ZN(n4212) );
  OAI211_X4 U3959 ( .C1(n2991), .C2(n2990), .A(n2989), .B(net329918), .ZN(
        n2992) );
  NAND2_X4 U3960 ( .A1(n2466), .A2(n2465), .ZN(net330742) );
  NAND2_X4 U3961 ( .A1(n2240), .A2(n2239), .ZN(n2421) );
  NAND2_X4 U3962 ( .A1(net330918), .A2(n2365), .ZN(net330855) );
  NAND2_X4 U3963 ( .A1(n2235), .A2(n2234), .ZN(n2540) );
  AOI21_X4 U3964 ( .B1(n3946), .B2(n1639), .A(n3945), .ZN(n4030) );
  NAND2_X4 U3965 ( .A1(n2309), .A2(n2310), .ZN(n2541) );
  NAND2_X4 U3966 ( .A1(n2173), .A2(n1717), .ZN(n2229) );
  AOI21_X2 U3967 ( .B1(n3526), .B2(n3525), .A(n3524), .ZN(n3530) );
  NAND2_X4 U3968 ( .A1(n1726), .A2(n2308), .ZN(n2536) );
  NAND2_X4 U3969 ( .A1(n2190), .A2(n2189), .ZN(n2349) );
  NAND2_X4 U3970 ( .A1(n2992), .A2(n2993), .ZN(n3083) );
  NAND2_X4 U3971 ( .A1(n3028), .A2(n2951), .ZN(net329859) );
  OAI21_X4 U3972 ( .B1(n3215), .B2(n3214), .A(n1826), .ZN(n3329) );
  NAND3_X2 U3973 ( .A1(net332668), .A2(net330131), .A3(net329992), .ZN(n2760)
         );
  NAND2_X4 U3975 ( .A1(n3719), .A2(n3967), .ZN(n3738) );
  NAND2_X4 U3976 ( .A1(n3717), .A2(n3718), .ZN(n3967) );
  OAI22_X4 U3977 ( .A1(n2761), .A2(n2760), .B1(net330234), .B2(n2759), .ZN(
        n2793) );
  INV_X4 U3978 ( .A(n3039), .ZN(n3043) );
  INV_X8 U3979 ( .A(n3777), .ZN(n3878) );
  OAI21_X2 U3980 ( .B1(n2278), .B2(n2279), .A(n2277), .ZN(n2287) );
  NOR2_X2 U3981 ( .A1(n1741), .A2(n2096), .ZN(n2103) );
  NAND2_X4 U3982 ( .A1(n2162), .A2(n2161), .ZN(n2573) );
  NAND2_X4 U3983 ( .A1(n4117), .A2(n1332), .ZN(net328259) );
  NAND2_X4 U3984 ( .A1(n3350), .A2(n3057), .ZN(n3116) );
  INV_X1 U3985 ( .A(n3331), .ZN(n3105) );
  NOR2_X4 U3986 ( .A1(n4213), .A2(n4214), .ZN(n4218) );
  OAI22_X4 U3987 ( .A1(n3185), .A2(n3184), .B1(n3183), .B2(n3182), .ZN(n4213)
         );
  OAI221_X4 U3988 ( .B1(n3254), .B2(n3255), .C1(n3253), .C2(n1743), .A(n3252), 
        .ZN(n3257) );
  INV_X1 U3989 ( .A(n3307), .ZN(n3306) );
  NAND2_X4 U3990 ( .A1(n3249), .A2(n3248), .ZN(n3254) );
  INV_X1 U3991 ( .A(n3217), .ZN(n3218) );
  NAND4_X2 U3992 ( .A1(n3241), .A2(n3345), .A3(net329456), .A4(n3431), .ZN(
        n3243) );
  NAND2_X4 U3993 ( .A1(n3257), .A2(n3256), .ZN(n3262) );
  NAND2_X4 U3994 ( .A1(n3679), .A2(n1759), .ZN(n3564) );
  NAND3_X2 U3995 ( .A1(n3344), .A2(n3431), .A3(n3345), .ZN(n3242) );
  INV_X32 U3996 ( .A(control[0]), .ZN(net331583) );
  NAND2_X4 U3997 ( .A1(n3443), .A2(n3117), .ZN(n3058) );
  NAND2_X4 U3998 ( .A1(n2897), .A2(n2898), .ZN(n3178) );
  NAND2_X4 U4000 ( .A1(n3117), .A2(n3118), .ZN(n3447) );
  NAND2_X4 U4001 ( .A1(n2040), .A2(n2039), .ZN(n2125) );
  NAND2_X4 U4002 ( .A1(n4063), .A2(n4064), .ZN(n4177) );
  NAND2_X4 U4003 ( .A1(n3985), .A2(n3986), .ZN(n4047) );
  INV_X8 U4004 ( .A(n2206), .ZN(n2039) );
  INV_X8 U4005 ( .A(n3594), .ZN(n3510) );
  NAND3_X2 U4006 ( .A1(n2873), .A2(net330098), .A3(n1146), .ZN(n2874) );
  NAND2_X4 U4007 ( .A1(n3063), .A2(n3064), .ZN(net329464) );
  XNOR2_X2 U4008 ( .A(net328603), .B(net328604), .ZN(n3768) );
  NAND2_X4 U4009 ( .A1(n3767), .A2(n1131), .ZN(net328603) );
  NAND3_X1 U4010 ( .A1(net328937), .A2(n3755), .A3(net328936), .ZN(n3714) );
  NAND2_X1 U4011 ( .A1(net328937), .A2(net328936), .ZN(n3853) );
  NAND2_X4 U4012 ( .A1(net329289), .A2(n3470), .ZN(n3605) );
  NAND2_X4 U4013 ( .A1(n2902), .A2(n2903), .ZN(n3175) );
  NAND2_X4 U4014 ( .A1(n2488), .A2(n2489), .ZN(n2490) );
  NAND2_X4 U4015 ( .A1(n2734), .A2(n2735), .ZN(n2737) );
  NAND2_X4 U4016 ( .A1(n3285), .A2(n3284), .ZN(n3591) );
  NAND2_X4 U4017 ( .A1(n2030), .A2(n3622), .ZN(n3624) );
  INV_X4 U4018 ( .A(n2029), .ZN(n2030) );
  NAND3_X2 U4019 ( .A1(n2487), .A2(n2387), .A3(n2541), .ZN(n2488) );
  NAND2_X2 U4020 ( .A1(n4237), .A2(n4243), .ZN(n4249) );
  NAND2_X4 U4021 ( .A1(n3379), .A2(net329404), .ZN(n3686) );
  NAND3_X4 U4022 ( .A1(n2138), .A2(net333879), .A3(net331068), .ZN(net330652)
         );
  OAI21_X4 U4023 ( .B1(n2659), .B2(n2658), .A(n1629), .ZN(n2457) );
  NOR2_X2 U4024 ( .A1(n2655), .A2(n2640), .ZN(n2641) );
  NAND2_X4 U4025 ( .A1(n3742), .A2(n3741), .ZN(n3932) );
  NOR2_X2 U4026 ( .A1(net330130), .A2(net330134), .ZN(net330126) );
  NAND2_X4 U4027 ( .A1(n1632), .A2(n3290), .ZN(n3505) );
  NAND2_X4 U4028 ( .A1(n3733), .A2(n3848), .ZN(n3739) );
  NAND2_X4 U4029 ( .A1(n3962), .A2(n3961), .ZN(n3752) );
  NAND2_X4 U4030 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  AOI21_X2 U4031 ( .B1(n4091), .B2(n4099), .A(net328160), .ZN(n4097) );
  NAND2_X4 U4032 ( .A1(n2094), .A2(n2112), .ZN(net331113) );
  NAND2_X4 U4033 ( .A1(n2092), .A2(n2093), .ZN(n2112) );
  NAND2_X4 U4034 ( .A1(n2047), .A2(n2046), .ZN(n2104) );
  NAND3_X4 U4035 ( .A1(n3843), .A2(n4228), .A3(n4230), .ZN(n4124) );
  NAND2_X4 U4036 ( .A1(n3391), .A2(n3390), .ZN(n3506) );
  INV_X1 U4037 ( .A(net332747), .ZN(net331506) );
  NAND2_X1 U4038 ( .A1(a[15]), .A2(n2125), .ZN(n2863) );
  NAND3_X4 U4039 ( .A1(n1314), .A2(n1761), .A3(n2556), .ZN(n2473) );
  NAND3_X2 U4040 ( .A1(n2909), .A2(n2911), .A3(n2910), .ZN(n2912) );
  OAI21_X4 U4041 ( .B1(net330612), .B2(n2204), .A(net330752), .ZN(n2231) );
  NAND2_X4 U4042 ( .A1(n2026), .A2(n2218), .ZN(n2178) );
  NAND2_X4 U4043 ( .A1(n3071), .A2(n3406), .ZN(n3195) );
  NAND2_X4 U4044 ( .A1(n2502), .A2(n2420), .ZN(n2627) );
  NAND2_X4 U4045 ( .A1(n2544), .A2(n2545), .ZN(n2633) );
  INV_X8 U4046 ( .A(net328105), .ZN(net331359) );
  INV_X16 U4047 ( .A(net331359), .ZN(net331357) );
  OAI22_X4 U4048 ( .A1(n2823), .A2(n2822), .B1(n2821), .B2(n2820), .ZN(n2902)
         );
  NAND3_X1 U4050 ( .A1(n1107), .A2(n1334), .A3(n3483), .ZN(n2727) );
  XOR2_X1 U4051 ( .A(n2399), .B(n2001), .Z(n2405) );
  NOR2_X4 U4052 ( .A1(n3510), .A2(n4455), .ZN(n3417) );
  NAND3_X2 U4053 ( .A1(n4076), .A2(net328388), .A3(n1397), .ZN(n4145) );
  NAND2_X4 U4054 ( .A1(n1958), .A2(n3473), .ZN(n3600) );
  NAND2_X4 U4055 ( .A1(n3378), .A2(net329397), .ZN(n3518) );
  NAND2_X4 U4056 ( .A1(n2652), .A2(n2653), .ZN(n2462) );
  NAND3_X2 U4057 ( .A1(n3006), .A2(n1707), .A3(n3007), .ZN(n3197) );
  NAND2_X4 U4058 ( .A1(n4027), .A2(n4028), .ZN(net328268) );
  NAND2_X4 U4059 ( .A1(net328013), .A2(n4295), .ZN(n4302) );
  NAND2_X1 U4060 ( .A1(n2467), .A2(net330510), .ZN(n2384) );
  NAND2_X4 U4061 ( .A1(n2069), .A2(n1348), .ZN(n4325) );
  NAND3_X2 U4062 ( .A1(n3490), .A2(n3489), .A3(n3488), .ZN(n4217) );
  NAND2_X4 U4063 ( .A1(n3505), .A2(n3325), .ZN(n4020) );
  NAND3_X2 U4064 ( .A1(n1729), .A2(n4449), .A3(n4086), .ZN(n4141) );
  NAND2_X4 U4065 ( .A1(n3336), .A2(n1859), .ZN(n3382) );
  NAND3_X4 U4067 ( .A1(n2663), .A2(n2561), .A3(n2665), .ZN(n2370) );
  NAND2_X4 U4068 ( .A1(n1614), .A2(n2313), .ZN(n2346) );
  OAI21_X2 U4069 ( .B1(n3404), .B2(n3504), .A(n3403), .ZN(n3482) );
  NAND2_X1 U4070 ( .A1(n3004), .A2(n3005), .ZN(n2977) );
  NAND2_X4 U4071 ( .A1(n2306), .A2(n2307), .ZN(n2465) );
  NAND2_X4 U4072 ( .A1(n2662), .A2(n2661), .ZN(net330331) );
  NAND2_X4 U4073 ( .A1(n1123), .A2(n4010), .ZN(net328573) );
  OAI21_X4 U4074 ( .B1(n2375), .B2(n2374), .A(n2568), .ZN(n2379) );
  NAND2_X4 U4075 ( .A1(n2553), .A2(n2554), .ZN(n2781) );
  NAND2_X4 U4076 ( .A1(n3388), .A2(n3389), .ZN(n3578) );
  NAND2_X4 U4078 ( .A1(n1657), .A2(n4209), .ZN(n3570) );
  OAI21_X1 U4079 ( .B1(n3827), .B2(n3960), .A(n3753), .ZN(n3823) );
  NAND3_X2 U4080 ( .A1(n1465), .A2(n3096), .A3(n3297), .ZN(n3163) );
  NAND2_X4 U4081 ( .A1(net330987), .A2(net330986), .ZN(net330863) );
  NAND2_X4 U4082 ( .A1(n2264), .A2(n2265), .ZN(n2426) );
  AOI22_X4 U4083 ( .A1(n2624), .A2(n2623), .B1(n2622), .B2(n2621), .ZN(n2821)
         );
  NOR2_X4 U4084 ( .A1(n3175), .A2(n3176), .ZN(n3185) );
  OAI22_X4 U4085 ( .A1(n2518), .A2(n2517), .B1(n2516), .B2(n2515), .ZN(n2519)
         );
  OAI22_X4 U4086 ( .A1(n2517), .A2(n2409), .B1(n2514), .B2(n2408), .ZN(n2515)
         );
  AOI221_X4 U4087 ( .B1(n2945), .B2(net329992), .C1(net330406), .C2(n2639), 
        .A(n2640), .ZN(n2642) );
  NAND2_X4 U4088 ( .A1(n1720), .A2(n2460), .ZN(n2652) );
  NAND2_X4 U4089 ( .A1(n4088), .A2(n4142), .ZN(net328177) );
  NAND2_X4 U4090 ( .A1(n4081), .A2(n4080), .ZN(n4136) );
  NAND2_X4 U4092 ( .A1(n2714), .A2(n2715), .ZN(n2958) );
  NAND2_X4 U4093 ( .A1(n2497), .A2(n2498), .ZN(n2828) );
  NAND2_X1 U4094 ( .A1(n2064), .A2(n1703), .ZN(n2068) );
  NAND2_X4 U4095 ( .A1(n2953), .A2(n2954), .ZN(n3103) );
  AOI21_X1 U4096 ( .B1(net328035), .B2(n4024), .A(n4023), .ZN(n4025) );
  OAI21_X1 U4097 ( .B1(n2422), .B2(n2423), .A(n2421), .ZN(n2424) );
  NAND2_X4 U4098 ( .A1(n2689), .A2(n2690), .ZN(net330338) );
  NAND2_X4 U4099 ( .A1(n3352), .A2(n3351), .ZN(n3150) );
  NAND2_X4 U4100 ( .A1(n4069), .A2(n4070), .ZN(n4147) );
  NAND2_X4 U4101 ( .A1(n2778), .A2(n2779), .ZN(net330024) );
  NAND2_X4 U4102 ( .A1(n1918), .A2(n4176), .ZN(n4066) );
  NAND3_X2 U4103 ( .A1(n3211), .A2(n3092), .A3(n3007), .ZN(n3209) );
  AOI21_X4 U4104 ( .B1(n3018), .B2(n3022), .A(n3017), .ZN(n3025) );
  NAND2_X4 U4105 ( .A1(n2276), .A2(n1354), .ZN(n2676) );
  NAND2_X4 U4106 ( .A1(n2212), .A2(n2280), .ZN(n2275) );
  OAI22_X4 U4107 ( .A1(n2126), .A2(n2211), .B1(net331090), .B2(net330173), 
        .ZN(n2212) );
  NAND2_X4 U4108 ( .A1(n3415), .A2(n3416), .ZN(n3594) );
  NAND2_X4 U4109 ( .A1(n3119), .A2(n1939), .ZN(n3351) );
  NAND2_X4 U4110 ( .A1(n2861), .A2(n1487), .ZN(n2866) );
  NAND2_X4 U4112 ( .A1(n1784), .A2(n3125), .ZN(n2868) );
  XNOR2_X1 U4113 ( .A(n1693), .B(n1362), .ZN(product_out[14]) );
  XNOR2_X1 U4114 ( .A(n3938), .B(n1361), .ZN(product_out[21]) );
  NAND3_X2 U4116 ( .A1(n2627), .A2(n2629), .A3(n1905), .ZN(n2609) );
  NAND2_X4 U4117 ( .A1(n2343), .A2(n2342), .ZN(n2266) );
  NAND2_X1 U4118 ( .A1(n4098), .A2(net332287), .ZN(n4106) );
  INV_X8 U4119 ( .A(n3765), .ZN(n4014) );
  NAND2_X4 U4120 ( .A1(net331025), .A2(n2157), .ZN(n2290) );
  NAND2_X4 U4121 ( .A1(n3024), .A2(n3025), .ZN(n3334) );
  OAI21_X4 U4122 ( .B1(n4259), .B2(net328393), .A(n4143), .ZN(net328331) );
  NAND2_X4 U4123 ( .A1(net330383), .A2(net330382), .ZN(net329994) );
  NAND2_X4 U4124 ( .A1(n3565), .A2(n3566), .ZN(n3580) );
  NAND3_X2 U4125 ( .A1(n4391), .A2(n4088), .A3(n4142), .ZN(n4143) );
  INV_X8 U4126 ( .A(n3040), .ZN(n3041) );
  NAND2_X4 U4127 ( .A1(n2864), .A2(n2865), .ZN(n2867) );
  NOR2_X1 U4128 ( .A1(net331293), .A2(n1999), .ZN(n3302) );
  INV_X2 U4129 ( .A(n1999), .ZN(n4019) );
  OAI211_X4 U4130 ( .C1(n2998), .C2(n3318), .A(n3321), .B(n3317), .ZN(n3324)
         );
  NAND2_X1 U4131 ( .A1(n3746), .A2(n3745), .ZN(n3927) );
  NAND3_X2 U4132 ( .A1(n1124), .A2(n1689), .A3(n2973), .ZN(n3671) );
  NAND2_X4 U4133 ( .A1(n2361), .A2(n2362), .ZN(n2436) );
  NAND2_X4 U4134 ( .A1(n3413), .A2(n1656), .ZN(n3507) );
  NAND2_X4 U4135 ( .A1(net328911), .A2(net328585), .ZN(net328790) );
  OAI211_X4 U4136 ( .C1(net334211), .C2(n2758), .A(n2002), .B(n2757), .ZN(
        n2847) );
  NAND2_X4 U4137 ( .A1(net328564), .A2(n4011), .ZN(net328235) );
  NAND2_X4 U4138 ( .A1(n3200), .A2(n3194), .ZN(n3316) );
  NAND2_X4 U4139 ( .A1(n3073), .A2(n3196), .ZN(n3200) );
  NAND2_X4 U4140 ( .A1(n2976), .A2(n3207), .ZN(n3004) );
  NAND2_X2 U4141 ( .A1(n2554), .A2(n2553), .ZN(n2786) );
  NAND3_X2 U4142 ( .A1(n1427), .A2(n3320), .A3(n3319), .ZN(n3322) );
  NAND2_X4 U4143 ( .A1(n2484), .A2(n2485), .ZN(n2546) );
  NAND2_X4 U4144 ( .A1(n1419), .A2(n2956), .ZN(n3211) );
  NAND2_X4 U4145 ( .A1(n2967), .A2(n2881), .ZN(n3212) );
  NAND2_X4 U4146 ( .A1(n2106), .A2(n2107), .ZN(n2216) );
  NAND2_X4 U4147 ( .A1(n2436), .A2(n2437), .ZN(n2784) );
  NAND2_X4 U4148 ( .A1(net328737), .A2(net328616), .ZN(net328751) );
  OAI211_X4 U4149 ( .C1(n1267), .C2(n3705), .A(n3707), .B(n3704), .ZN(n3712)
         );
  NAND2_X4 U4150 ( .A1(n3522), .A2(n3523), .ZN(net329019) );
  NAND3_X4 U4151 ( .A1(n3438), .A2(n3437), .A3(n3436), .ZN(n3467) );
  NAND2_X4 U4152 ( .A1(n4305), .A2(n4304), .ZN(n4361) );
  NAND3_X2 U4153 ( .A1(n4141), .A2(n4140), .A3(n4139), .ZN(n4088) );
  NAND2_X4 U4154 ( .A1(n2481), .A2(n2480), .ZN(n2637) );
  OAI211_X4 U4155 ( .C1(n2438), .C2(n2439), .A(n2555), .B(n2556), .ZN(n2459)
         );
  NAND2_X4 U4156 ( .A1(n3280), .A2(n3281), .ZN(n3426) );
  NAND2_X4 U4157 ( .A1(n2158), .A2(n2168), .ZN(n2679) );
  NAND2_X4 U4158 ( .A1(n1979), .A2(n3658), .ZN(n3754) );
  NAND2_X4 U4159 ( .A1(n3916), .A2(n3917), .ZN(n4094) );
  OAI22_X4 U4160 ( .A1(n3522), .A2(n3523), .B1(n1727), .B2(n3468), .ZN(
        net329018) );
  NAND3_X2 U4161 ( .A1(n3349), .A2(n3348), .A3(net329441), .ZN(n3432) );
  NAND3_X2 U4162 ( .A1(n4237), .A2(n3834), .A3(n4238), .ZN(n3836) );
  NAND2_X1 U4164 ( .A1(n2651), .A2(n4464), .ZN(n2458) );
  NAND3_X2 U4165 ( .A1(n2663), .A2(n2561), .A3(n2665), .ZN(n2572) );
  NAND2_X4 U4167 ( .A1(n3020), .A2(n1935), .ZN(n2889) );
  OAI22_X4 U4168 ( .A1(n1244), .A2(n2750), .B1(n1472), .B2(n2749), .ZN(n2751)
         );
  OAI211_X4 U4169 ( .C1(n3204), .C2(n1659), .A(n3203), .B(n1191), .ZN(n3298)
         );
  NAND2_X4 U4170 ( .A1(n3307), .A2(n3494), .ZN(n3488) );
  NAND2_X4 U4171 ( .A1(n2318), .A2(n2319), .ZN(n2417) );
  NAND2_X4 U4172 ( .A1(n2988), .A2(n2987), .ZN(n3318) );
  NAND2_X4 U4173 ( .A1(n2103), .A2(n2102), .ZN(net331070) );
  NAND2_X4 U4174 ( .A1(n2422), .A2(n2423), .ZN(n2746) );
  NAND2_X4 U4175 ( .A1(n3016), .A2(n3015), .ZN(n3102) );
  NAND2_X1 U4176 ( .A1(a[6]), .A2(n2125), .ZN(n2127) );
  NAND2_X4 U4177 ( .A1(n2810), .A2(n1737), .ZN(n3005) );
  NAND2_X4 U4178 ( .A1(n3119), .A2(n1939), .ZN(n3443) );
  NAND2_X4 U4179 ( .A1(n3889), .A2(n3885), .ZN(n3972) );
  NAND2_X4 U4180 ( .A1(n4071), .A2(n4147), .ZN(n4148) );
  NAND2_X4 U4182 ( .A1(n2683), .A2(n2684), .ZN(n2766) );
  NAND2_X4 U4184 ( .A1(n2757), .A2(n2002), .ZN(n2945) );
  NAND2_X4 U4185 ( .A1(n2880), .A2(n2879), .ZN(n2910) );
  NAND2_X4 U4186 ( .A1(n1405), .A2(n3727), .ZN(n3963) );
  NAND2_X4 U4187 ( .A1(n3526), .A2(n3525), .ZN(n3622) );
  NAND2_X4 U4188 ( .A1(n3432), .A2(n1193), .ZN(n3525) );
  NAND2_X4 U4189 ( .A1(n3654), .A2(n3655), .ZN(net328738) );
  NAND2_X4 U4190 ( .A1(n3651), .A2(n3652), .ZN(net328872) );
  NAND2_X4 U4191 ( .A1(n2358), .A2(n2359), .ZN(net330509) );
  NAND2_X4 U4192 ( .A1(n2434), .A2(n2435), .ZN(net330595) );
  NAND2_X4 U4194 ( .A1(n3480), .A2(n3481), .ZN(n3726) );
  NAND2_X4 U4195 ( .A1(n1741), .A2(n2216), .ZN(n2674) );
  NAND3_X2 U4197 ( .A1(n2963), .A2(n2831), .A3(n1286), .ZN(n2832) );
  NAND2_X4 U4198 ( .A1(n3737), .A2(n3736), .ZN(n4226) );
  NAND2_X4 U4199 ( .A1(n2613), .A2(n2614), .ZN(n2731) );
  OAI211_X4 U4200 ( .C1(n2738), .C2(n1916), .A(n2737), .B(n2736), .ZN(n2740)
         );
  NAND3_X2 U4201 ( .A1(net332364), .A2(net333621), .A3(n2548), .ZN(n2638) );
  NAND2_X4 U4202 ( .A1(n2606), .A2(n2605), .ZN(n2962) );
  OAI211_X4 U4204 ( .C1(n2984), .C2(n2983), .A(n2981), .B(n1687), .ZN(n3315)
         );
  NAND2_X4 U4205 ( .A1(n1671), .A2(n1124), .ZN(n2981) );
  NAND2_X1 U4206 ( .A1(n4470), .A2(net328158), .ZN(n4370) );
  NAND2_X4 U4207 ( .A1(n2873), .A2(net330098), .ZN(n2845) );
  NAND3_X2 U4208 ( .A1(n2552), .A2(n2790), .A3(n2789), .ZN(n2920) );
  NOR2_X1 U4209 ( .A1(n1173), .A2(net331896), .ZN(n4098) );
  NAND3_X2 U4210 ( .A1(n3597), .A2(n3596), .A3(n3680), .ZN(n3598) );
  NAND2_X1 U4211 ( .A1(a[4]), .A2(n1640), .ZN(n2160) );
  OAI21_X4 U4212 ( .B1(n2470), .B2(net330596), .A(net330598), .ZN(n2482) );
  OAI211_X4 U4213 ( .C1(n2675), .C2(n2674), .A(n1724), .B(n2573), .ZN(n2169)
         );
  NAND2_X4 U4214 ( .A1(n3089), .A2(n3090), .ZN(n3408) );
  OAI211_X4 U4215 ( .C1(n1971), .C2(n3968), .A(n3966), .B(n1666), .ZN(n4099)
         );
  NAND2_X4 U4216 ( .A1(n2649), .A2(n2648), .ZN(net330037) );
  NAND2_X4 U4217 ( .A1(n3013), .A2(n3014), .ZN(n3022) );
  NAND2_X4 U4218 ( .A1(n2588), .A2(n2589), .ZN(net330028) );
  NAND2_X4 U4219 ( .A1(n1947), .A2(n4256), .ZN(net328142) );
  NAND2_X4 U4220 ( .A1(n2946), .A2(net329986), .ZN(net329454) );
  NAND2_X4 U4222 ( .A1(n2040), .A2(n2039), .ZN(n2032) );
  NAND2_X4 U4223 ( .A1(n2947), .A2(n2948), .ZN(net329456) );
  INV_X32 U4224 ( .A(net331353), .ZN(net331349) );
  NAND3_X4 U4225 ( .A1(n4425), .A2(control[0]), .A3(b[16]), .ZN(n2043) );
  NAND3_X4 U4226 ( .A1(control[0]), .A2(control[1]), .A3(b[0]), .ZN(n2045) );
  INV_X4 U4227 ( .A(net329043), .ZN(net331287) );
  MUX2_X2 U4228 ( .A(product_in[0]), .B(net331287), .S(net331299), .Z(
        product_out[0]) );
  NAND2_X2 U4229 ( .A1(n1376), .A2(a[0]), .ZN(n2048) );
  NAND2_X2 U4230 ( .A1(a[1]), .A2(n2125), .ZN(net331271) );
  INV_X4 U4231 ( .A(n3816), .ZN(n2038) );
  MUX2_X2 U4232 ( .A(product_in[1]), .B(n2038), .S(net331299), .Z(
        product_out[1]) );
  NAND2_X2 U4233 ( .A1(net331262), .A2(net331131), .ZN(n3173) );
  INV_X4 U4234 ( .A(n3173), .ZN(n3920) );
  MUX2_X2 U4235 ( .A(product_in[2]), .B(n3920), .S(net331299), .Z(
        product_out[2]) );
  XNOR2_X2 U4236 ( .A(n2050), .B(n2049), .ZN(n2097) );
  OAI21_X4 U4237 ( .B1(n2052), .B2(net331247), .A(n2051), .ZN(net331227) );
  NAND3_X2 U4238 ( .A1(n2062), .A2(n2061), .A3(n1679), .ZN(net331130) );
  NAND2_X2 U4239 ( .A1(b[11]), .A2(net331362), .ZN(net331221) );
  NAND2_X2 U4240 ( .A1(a[0]), .A2(net331343), .ZN(n2064) );
  INV_X4 U4242 ( .A(n4022), .ZN(n3300) );
  MUX2_X2 U4243 ( .A(product_in[3]), .B(n3300), .S(net331299), .Z(
        product_out[3]) );
  NAND2_X2 U4244 ( .A1(a[2]), .A2(net331228), .ZN(net330998) );
  INV_X4 U4245 ( .A(net330998), .ZN(net331124) );
  INV_X4 U4246 ( .A(a[1]), .ZN(net331213) );
  INV_X4 U4247 ( .A(net331202), .ZN(net331196) );
  NOR2_X4 U4248 ( .A1(n4427), .A2(net331201), .ZN(n2075) );
  INV_X4 U4249 ( .A(net331199), .ZN(net331198) );
  INV_X4 U4250 ( .A(a[4]), .ZN(net331189) );
  AOI21_X4 U4251 ( .B1(n2079), .B2(n2078), .A(net331189), .ZN(n2105) );
  INV_X4 U4252 ( .A(net330990), .ZN(net331182) );
  NAND2_X2 U4253 ( .A1(a[1]), .A2(net331341), .ZN(n2083) );
  INV_X4 U4254 ( .A(n2083), .ZN(n2093) );
  NAND2_X2 U4255 ( .A1(n2110), .A2(n2112), .ZN(n2085) );
  XNOR2_X2 U4256 ( .A(n2085), .B(n2091), .ZN(n2087) );
  NAND2_X2 U4257 ( .A1(b[12]), .A2(net331362), .ZN(net331169) );
  NAND2_X2 U4258 ( .A1(a[0]), .A2(net331329), .ZN(n2086) );
  INV_X4 U4259 ( .A(n2086), .ZN(n2089) );
  INV_X4 U4260 ( .A(n2087), .ZN(n2088) );
  NAND2_X2 U4261 ( .A1(n2090), .A2(n4453), .ZN(n4108) );
  INV_X4 U4262 ( .A(n4108), .ZN(n2526) );
  MUX2_X2 U4263 ( .A(product_in[4]), .B(n2526), .S(net331299), .Z(
        product_out[4]) );
  OAI21_X4 U4264 ( .B1(n2093), .B2(n2092), .A(n4429), .ZN(n2094) );
  INV_X4 U4265 ( .A(a[4]), .ZN(net331138) );
  XNOR2_X2 U4266 ( .A(n2134), .B(n2095), .ZN(n2215) );
  NAND3_X2 U4267 ( .A1(n2099), .A2(n2098), .A3(n1207), .ZN(n2100) );
  NOR2_X4 U4268 ( .A1(a[4]), .A2(a[3]), .ZN(n2109) );
  NAND2_X2 U4269 ( .A1(a[2]), .A2(net331341), .ZN(net331098) );
  NAND2_X2 U4270 ( .A1(a[1]), .A2(net331329), .ZN(n2115) );
  OAI21_X4 U4271 ( .B1(net331115), .B2(n2114), .A(n2115), .ZN(n2142) );
  INV_X4 U4272 ( .A(n2115), .ZN(n2116) );
  NAND2_X2 U4273 ( .A1(n2142), .A2(n4438), .ZN(n2118) );
  XNOR2_X2 U4274 ( .A(n2118), .B(n4453), .ZN(n2120) );
  NAND2_X2 U4275 ( .A1(a[0]), .A2(net331323), .ZN(n2119) );
  NAND2_X2 U4276 ( .A1(n4439), .A2(n2119), .ZN(n2123) );
  INV_X4 U4277 ( .A(n2119), .ZN(n2122) );
  INV_X4 U4278 ( .A(n2120), .ZN(n2121) );
  NAND2_X2 U4279 ( .A1(n2123), .A2(n2244), .ZN(n2124) );
  INV_X4 U4280 ( .A(n2124), .ZN(n4195) );
  MUX2_X2 U4281 ( .A(product_in[5]), .B(n4195), .S(net331299), .Z(
        product_out[5]) );
  NAND2_X2 U4282 ( .A1(a[1]), .A2(net331323), .ZN(n2193) );
  INV_X4 U4283 ( .A(a[5]), .ZN(net331091) );
  OAI21_X4 U4284 ( .B1(n2128), .B2(n2127), .A(net330834), .ZN(n2166) );
  NAND3_X2 U4285 ( .A1(n2132), .A2(n2133), .A3(n2216), .ZN(n2136) );
  NAND2_X2 U4286 ( .A1(a[4]), .A2(n2034), .ZN(net331073) );
  NAND2_X2 U4287 ( .A1(a[2]), .A2(net331329), .ZN(n2139) );
  INV_X4 U4288 ( .A(n2139), .ZN(n2140) );
  NAND2_X2 U4289 ( .A1(n2189), .A2(n2348), .ZN(n2145) );
  INV_X4 U4290 ( .A(n2141), .ZN(n2143) );
  NAND2_X2 U4291 ( .A1(n2242), .A2(n2243), .ZN(n2147) );
  XNOR2_X2 U4292 ( .A(n2147), .B(n2244), .ZN(n2152) );
  NAND2_X2 U4293 ( .A1(b[14]), .A2(net331362), .ZN(n2150) );
  NAND2_X2 U4294 ( .A1(b[6]), .A2(net331299), .ZN(n2149) );
  AOI22_X2 U4295 ( .A1(b[30]), .A2(net331613), .B1(b[22]), .B2(net328035), 
        .ZN(n2148) );
  NAND2_X2 U4296 ( .A1(a[0]), .A2(n2037), .ZN(n2151) );
  INV_X4 U4298 ( .A(n2151), .ZN(n2154) );
  INV_X4 U4299 ( .A(n2152), .ZN(n2153) );
  INV_X4 U4302 ( .A(net328250), .ZN(net331037) );
  MUX2_X2 U4303 ( .A(product_in[6]), .B(net331037), .S(net331299), .Z(
        product_out[6]) );
  NAND2_X2 U4304 ( .A1(a[1]), .A2(n2037), .ZN(n2196) );
  NAND2_X2 U4305 ( .A1(a[3]), .A2(net331329), .ZN(n2350) );
  INV_X4 U4306 ( .A(n2350), .ZN(n2354) );
  NAND2_X2 U4307 ( .A1(n2162), .A2(n2161), .ZN(n2158) );
  INV_X4 U4308 ( .A(n2163), .ZN(n2677) );
  OAI21_X4 U4309 ( .B1(n2680), .B2(n1110), .A(n2165), .ZN(n2205) );
  AOI21_X4 U4310 ( .B1(n1147), .B2(n2178), .A(n2166), .ZN(n2170) );
  NAND2_X2 U4311 ( .A1(a[5]), .A2(n2034), .ZN(n2228) );
  NOR2_X4 U4313 ( .A1(net330999), .A2(net331000), .ZN(n2181) );
  NAND2_X2 U4314 ( .A1(a[4]), .A2(net331341), .ZN(net330751) );
  INV_X4 U4315 ( .A(net330751), .ZN(net330986) );
  XNOR2_X2 U4316 ( .A(n2183), .B(n2184), .ZN(n2351) );
  NAND2_X2 U4317 ( .A1(n2354), .A2(net330983), .ZN(n2186) );
  OAI21_X4 U4318 ( .B1(n2353), .B2(n2354), .A(n1694), .ZN(n2246) );
  XNOR2_X2 U4319 ( .A(n2269), .B(n1339), .ZN(n2191) );
  XNOR2_X2 U4320 ( .A(n2199), .B(n2254), .ZN(net330965) );
  INV_X4 U4321 ( .A(net330965), .ZN(net330876) );
  NAND2_X2 U4322 ( .A1(b[15]), .A2(net331362), .ZN(n2202) );
  NAND2_X2 U4323 ( .A1(b[7]), .A2(net331299), .ZN(n2201) );
  AOI22_X2 U4324 ( .A1(b[31]), .A2(net331613), .B1(b[23]), .B2(net328035), 
        .ZN(n2200) );
  NAND2_X2 U4325 ( .A1(product_in[8]), .A2(net331295), .ZN(n2332) );
  AOI22_X2 U4326 ( .A1(n2203), .A2(n2268), .B1(n2268), .B2(n2246), .ZN(n2238)
         );
  NAND2_X2 U4327 ( .A1(a[4]), .A2(net331329), .ZN(n2234) );
  INV_X4 U4328 ( .A(n2234), .ZN(n2233) );
  NAND2_X2 U4329 ( .A1(net332690), .A2(n1902), .ZN(n2222) );
  INV_X4 U4330 ( .A(a[8]), .ZN(n2211) );
  INV_X4 U4331 ( .A(a[7]), .ZN(net330173) );
  NAND3_X2 U4332 ( .A1(n2221), .A2(n2220), .A3(net333816), .ZN(n2223) );
  OAI21_X4 U4333 ( .B1(n2282), .B2(n2225), .A(n2224), .ZN(n2226) );
  NAND2_X2 U4334 ( .A1(a[5]), .A2(net331341), .ZN(net330912) );
  XNOR2_X2 U4335 ( .A(net330917), .B(net330916), .ZN(net330911) );
  INV_X4 U4336 ( .A(net330855), .ZN(net330915) );
  AOI21_X4 U4337 ( .B1(n2230), .B2(n1618), .A(net330915), .ZN(net330913) );
  XNOR2_X2 U4338 ( .A(n2231), .B(net330910), .ZN(n2235) );
  INV_X4 U4339 ( .A(n1886), .ZN(n2232) );
  NAND2_X2 U4340 ( .A1(a[3]), .A2(net331323), .ZN(n2239) );
  INV_X4 U4341 ( .A(n2239), .ZN(n2265) );
  INV_X4 U4342 ( .A(n2242), .ZN(n2245) );
  OAI21_X4 U4343 ( .B1(n2245), .B2(n2244), .A(n2243), .ZN(n2342) );
  XNOR2_X2 U4344 ( .A(n2249), .B(n2425), .ZN(n2252) );
  NAND2_X2 U4345 ( .A1(a[2]), .A2(n2037), .ZN(n2251) );
  INV_X4 U4346 ( .A(n2251), .ZN(n2253) );
  NAND2_X2 U4347 ( .A1(n2414), .A2(n2012), .ZN(n2258) );
  INV_X4 U4349 ( .A(n2261), .ZN(n2259) );
  NAND2_X2 U4350 ( .A1(a[1]), .A2(net331305), .ZN(n2260) );
  INV_X4 U4351 ( .A(n2260), .ZN(n2262) );
  NAND2_X2 U4352 ( .A1(n2262), .A2(n2261), .ZN(n2325) );
  XNOR2_X2 U4353 ( .A(n2263), .B(net330786), .ZN(n2907) );
  OAI22_X2 U4354 ( .A1(net331363), .A2(net329043), .B1(n2907), .B2(net331293), 
        .ZN(n2333) );
  XNOR2_X2 U4355 ( .A(n2332), .B(n2333), .ZN(product_out[8]) );
  INV_X4 U4356 ( .A(net330861), .ZN(net330860) );
  INV_X4 U4357 ( .A(n1163), .ZN(n2361) );
  NAND2_X2 U4358 ( .A1(n2362), .A2(n2361), .ZN(n2300) );
  INV_X4 U4359 ( .A(n2300), .ZN(n2273) );
  NAND2_X2 U4360 ( .A1(a[6]), .A2(net331341), .ZN(n2307) );
  NOR2_X4 U4361 ( .A1(a[4]), .A2(a[3]), .ZN(n2277) );
  OAI21_X4 U4362 ( .B1(n2164), .B2(n1161), .A(n2280), .ZN(n2849) );
  NAND2_X2 U4363 ( .A1(a[8]), .A2(net331357), .ZN(n2283) );
  OAI21_X4 U4364 ( .B1(n2286), .B2(n2285), .A(n1704), .ZN(n2295) );
  NOR2_X4 U4365 ( .A1(n1721), .A2(n2288), .ZN(n2289) );
  INV_X4 U4366 ( .A(n2440), .ZN(n2293) );
  NAND2_X2 U4367 ( .A1(n2360), .A2(n2437), .ZN(n2304) );
  INV_X4 U4368 ( .A(n2307), .ZN(n2359) );
  NAND2_X2 U4369 ( .A1(n2304), .A2(n2359), .ZN(n2296) );
  XNOR2_X2 U4370 ( .A(n2297), .B(n2296), .ZN(n2466) );
  NAND2_X2 U4371 ( .A1(net330650), .A2(net330649), .ZN(n2298) );
  INV_X4 U4372 ( .A(n2298), .ZN(n2363) );
  NAND3_X2 U4373 ( .A1(n2299), .A2(n2471), .A3(net330595), .ZN(n2302) );
  NAND3_X2 U4374 ( .A1(net330738), .A2(net330595), .A3(n1617), .ZN(n2301) );
  XNOR2_X2 U4375 ( .A(net330808), .B(n2469), .ZN(n2309) );
  NAND2_X2 U4376 ( .A1(a[5]), .A2(net331329), .ZN(n2308) );
  INV_X4 U4377 ( .A(n2308), .ZN(n2310) );
  XNOR2_X2 U4378 ( .A(n2312), .B(n2311), .ZN(n2422) );
  NAND2_X2 U4379 ( .A1(a[4]), .A2(net331323), .ZN(n2313) );
  INV_X4 U4380 ( .A(n2313), .ZN(n2423) );
  NAND2_X2 U4381 ( .A1(a[3]), .A2(n2037), .ZN(n2316) );
  INV_X4 U4382 ( .A(n2316), .ZN(n2319) );
  XNOR2_X2 U4383 ( .A(n2400), .B(n2404), .ZN(n2323) );
  NAND2_X2 U4384 ( .A1(n2321), .A2(n2320), .ZN(n2322) );
  XNOR2_X2 U4385 ( .A(n2323), .B(n1676), .ZN(n2401) );
  INV_X4 U4386 ( .A(n2324), .ZN(n2326) );
  OAI21_X4 U4387 ( .B1(n2326), .B2(net330786), .A(n2325), .ZN(n2402) );
  XNOR2_X2 U4388 ( .A(n2401), .B(n2402), .ZN(n3815) );
  NAND2_X2 U4389 ( .A1(product_in[9]), .A2(net331295), .ZN(n2328) );
  INV_X4 U4390 ( .A(n2328), .ZN(n2330) );
  INV_X4 U4391 ( .A(n2332), .ZN(n2334) );
  NAND2_X2 U4392 ( .A1(n2334), .A2(n2333), .ZN(n2338) );
  XNOR2_X2 U4393 ( .A(n2335), .B(n2338), .ZN(product_out[9]) );
  NAND2_X2 U4394 ( .A1(product_in[10]), .A2(net331295), .ZN(n2517) );
  NAND2_X2 U4395 ( .A1(n3920), .A2(net331362), .ZN(n2409) );
  INV_X4 U4396 ( .A(n2517), .ZN(n2408) );
  INV_X4 U4397 ( .A(n2399), .ZN(n2340) );
  NAND3_X4 U4398 ( .A1(n2346), .A2(n2347), .A3(n2421), .ZN(n2745) );
  INV_X4 U4399 ( .A(n2352), .ZN(n2357) );
  OAI21_X4 U4400 ( .B1(n2357), .B2(n2356), .A(n2355), .ZN(n2537) );
  NAND2_X2 U4401 ( .A1(n2541), .A2(n2487), .ZN(n2388) );
  INV_X4 U4402 ( .A(a[10]), .ZN(n2376) );
  NAND2_X2 U4404 ( .A1(a[8]), .A2(n2034), .ZN(n2381) );
  INV_X4 U4405 ( .A(n2381), .ZN(n2554) );
  NAND2_X2 U4406 ( .A1(a[7]), .A2(net331341), .ZN(net330513) );
  NAND2_X2 U4407 ( .A1(a[6]), .A2(net331329), .ZN(n2385) );
  INV_X4 U4408 ( .A(n2385), .ZN(n2485) );
  INV_X4 U4409 ( .A(n2529), .ZN(n2429) );
  NAND2_X2 U4410 ( .A1(a[5]), .A2(net331323), .ZN(n2428) );
  INV_X4 U4411 ( .A(n2428), .ZN(n2530) );
  XNOR2_X2 U4412 ( .A(n2389), .B(n2390), .ZN(n2411) );
  NAND2_X2 U4413 ( .A1(a[4]), .A2(n2037), .ZN(n2391) );
  INV_X4 U4414 ( .A(n2391), .ZN(n2412) );
  NAND2_X2 U4415 ( .A1(a[3]), .A2(net331307), .ZN(n2396) );
  INV_X4 U4416 ( .A(n2396), .ZN(n2398) );
  XNOR2_X2 U4417 ( .A(n2406), .B(n2507), .ZN(n2407) );
  OAI21_X4 U4418 ( .B1(n3923), .B2(net331295), .A(n2409), .ZN(n2514) );
  XNOR2_X2 U4419 ( .A(n1880), .B(n2410), .ZN(product_out[10]) );
  NAND2_X2 U4420 ( .A1(n3300), .A2(net331362), .ZN(n2523) );
  INV_X4 U4421 ( .A(n2415), .ZN(n2419) );
  OAI21_X4 U4422 ( .B1(n2419), .B2(n2418), .A(n1983), .ZN(n2502) );
  NAND3_X2 U4423 ( .A1(n2427), .A2(n2426), .A3(n2746), .ZN(n2431) );
  NAND3_X2 U4424 ( .A1(n2432), .A2(n2431), .A3(n2430), .ZN(n2433) );
  NAND2_X2 U4425 ( .A1(a[6]), .A2(net331323), .ZN(n2493) );
  INV_X4 U4426 ( .A(n2493), .ZN(n2492) );
  NAND2_X2 U4427 ( .A1(a[8]), .A2(net331343), .ZN(n2477) );
  NAND2_X2 U4428 ( .A1(net330595), .A2(net330204), .ZN(n2439) );
  NAND3_X2 U4429 ( .A1(n2442), .A2(n2561), .A3(n2665), .ZN(n2446) );
  NAND3_X2 U4430 ( .A1(n2446), .A2(n2445), .A3(n2444), .ZN(n2449) );
  NAND2_X2 U4431 ( .A1(a[9]), .A2(n2034), .ZN(n2453) );
  OAI21_X4 U4432 ( .B1(n2452), .B2(n2451), .A(n2453), .ZN(n2918) );
  INV_X4 U4433 ( .A(n2453), .ZN(n2456) );
  INV_X4 U4434 ( .A(n2477), .ZN(n2651) );
  INV_X4 U4435 ( .A(n2458), .ZN(n2653) );
  NAND2_X2 U4436 ( .A1(n2651), .A2(n2476), .ZN(n2461) );
  XNOR2_X2 U4437 ( .A(n2462), .B(n2461), .ZN(n2481) );
  NAND2_X2 U4438 ( .A1(a[7]), .A2(net331329), .ZN(n2483) );
  INV_X4 U4439 ( .A(n2483), .ZN(n2545) );
  NAND3_X4 U4440 ( .A1(n2785), .A2(net333501), .A3(net333869), .ZN(n2552) );
  NAND2_X2 U4442 ( .A1(a[5]), .A2(n2037), .ZN(n2498) );
  INV_X4 U4443 ( .A(n2498), .ZN(n2500) );
  XNOR2_X2 U4444 ( .A(n2501), .B(n2607), .ZN(n2528) );
  XNOR2_X2 U4445 ( .A(n2505), .B(n2504), .ZN(n2506) );
  INV_X4 U4446 ( .A(n2508), .ZN(n2510) );
  NAND2_X2 U4448 ( .A1(product_in[11]), .A2(net331295), .ZN(n2522) );
  INV_X4 U4449 ( .A(n2522), .ZN(n2512) );
  XNOR2_X2 U4450 ( .A(n2513), .B(n2512), .ZN(n2521) );
  NOR2_X4 U4451 ( .A1(n2520), .A2(n2521), .ZN(n2525) );
  NOR2_X4 U4452 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  NOR2_X4 U4453 ( .A1(n2525), .A2(n2524), .ZN(n2620) );
  NAND2_X2 U4454 ( .A1(product_in[12]), .A2(net331295), .ZN(n2618) );
  NAND2_X2 U4455 ( .A1(n2526), .A2(net331362), .ZN(n2617) );
  INV_X4 U4456 ( .A(n2618), .ZN(n2622) );
  INV_X4 U4457 ( .A(n2724), .ZN(n2733) );
  OAI22_X2 U4458 ( .A1(n2723), .A2(n2733), .B1(n2722), .B2(n2733), .ZN(n2616)
         );
  NAND2_X2 U4459 ( .A1(a[7]), .A2(net331323), .ZN(n2599) );
  INV_X4 U4460 ( .A(n2599), .ZN(n2750) );
  NAND2_X2 U4461 ( .A1(n2542), .A2(n2541), .ZN(n2645) );
  NAND2_X2 U4462 ( .A1(a[8]), .A2(net331329), .ZN(n2640) );
  INV_X4 U4463 ( .A(n2640), .ZN(n2594) );
  NAND3_X4 U4464 ( .A1(n2566), .A2(n2565), .A3(n1862), .ZN(n2686) );
  OAI21_X4 U4465 ( .B1(n2577), .B2(n2576), .A(n2575), .ZN(n2664) );
  NOR2_X4 U4466 ( .A1(n2581), .A2(n2580), .ZN(n2585) );
  INV_X4 U4467 ( .A(a[11]), .ZN(n2583) );
  NAND3_X4 U4468 ( .A1(n2584), .A2(a[11]), .A3(net331349), .ZN(n2855) );
  NAND2_X2 U4469 ( .A1(a[10]), .A2(n2034), .ZN(n2586) );
  INV_X4 U4470 ( .A(n2586), .ZN(n2589) );
  INV_X4 U4471 ( .A(n2596), .ZN(n2597) );
  NAND2_X2 U4472 ( .A1(n2750), .A2(n2749), .ZN(n2711) );
  NAND2_X2 U4473 ( .A1(n2711), .A2(n3019), .ZN(n2601) );
  NAND2_X2 U4474 ( .A1(a[6]), .A2(n2037), .ZN(n2603) );
  INV_X4 U4475 ( .A(n2603), .ZN(n2606) );
  NAND2_X2 U4476 ( .A1(n2607), .A2(n1905), .ZN(n2608) );
  NAND2_X2 U4477 ( .A1(a[5]), .A2(net331307), .ZN(n2611) );
  INV_X4 U4478 ( .A(n2611), .ZN(n2614) );
  XNOR2_X2 U4479 ( .A(n2616), .B(n1917), .ZN(n4107) );
  OAI21_X4 U4480 ( .B1(n4107), .B2(net331295), .A(n2617), .ZN(n2621) );
  NAND2_X2 U4482 ( .A1(product_in[13]), .A2(net331293), .ZN(n2822) );
  NAND2_X2 U4483 ( .A1(n4195), .A2(net331362), .ZN(n2823) );
  INV_X4 U4484 ( .A(n2823), .ZN(n2625) );
  AOI21_X4 U4485 ( .B1(n2822), .B2(net331293), .A(n2625), .ZN(n2729) );
  INV_X4 U4486 ( .A(n2822), .ZN(n2626) );
  INV_X4 U4487 ( .A(n2631), .ZN(n2635) );
  NAND2_X2 U4488 ( .A1(a[8]), .A2(net331323), .ZN(n3010) );
  INV_X4 U4489 ( .A(n3010), .ZN(n2755) );
  NAND2_X2 U4490 ( .A1(n2651), .A2(n2650), .ZN(n2654) );
  XNOR2_X2 U4491 ( .A(n2654), .B(n1416), .ZN(net330382) );
  NAND2_X2 U4492 ( .A1(a[10]), .A2(net331343), .ZN(net330330) );
  AND2_X2 U4493 ( .A1(n2855), .A2(n2769), .ZN(n2667) );
  NOR2_X4 U4494 ( .A1(n2673), .A2(n2672), .ZN(n2690) );
  OAI21_X4 U4495 ( .B1(n2680), .B2(n1110), .A(n2678), .ZN(n2852) );
  INV_X4 U4496 ( .A(n2769), .ZN(n2681) );
  NAND3_X4 U4497 ( .A1(n2686), .A2(n2769), .A3(n2685), .ZN(n2932) );
  NAND2_X2 U4498 ( .A1(a[11]), .A2(n2034), .ZN(net330334) );
  INV_X4 U4499 ( .A(net330334), .ZN(net330336) );
  NAND3_X4 U4500 ( .A1(net330337), .A2(net330338), .A3(net330336), .ZN(
        net330025) );
  NAND2_X2 U4501 ( .A1(a[9]), .A2(net331329), .ZN(n2839) );
  INV_X4 U4502 ( .A(n2839), .ZN(n2695) );
  XNOR2_X2 U4503 ( .A(n2697), .B(n2696), .ZN(n2705) );
  XNOR2_X2 U4504 ( .A(n2704), .B(n1406), .ZN(n2753) );
  XNOR2_X2 U4506 ( .A(n2712), .B(n2713), .ZN(n2826) );
  NAND2_X2 U4507 ( .A1(a[7]), .A2(n2037), .ZN(n2715) );
  INV_X4 U4508 ( .A(n2715), .ZN(n2827) );
  XNOR2_X2 U4509 ( .A(n2717), .B(n2716), .ZN(n2720) );
  NAND2_X2 U4510 ( .A1(a[6]), .A2(net331307), .ZN(n2719) );
  INV_X4 U4511 ( .A(n2719), .ZN(n2721) );
  NAND3_X4 U4513 ( .A1(n3484), .A2(n1334), .A3(n2725), .ZN(n2726) );
  NOR2_X4 U4514 ( .A1(n2738), .A2(n2733), .ZN(n2735) );
  NOR2_X4 U4515 ( .A1(n2742), .A2(n2741), .ZN(n2744) );
  INV_X4 U4516 ( .A(n2886), .ZN(n2756) );
  NAND2_X2 U4517 ( .A1(a[10]), .A2(net331329), .ZN(n2796) );
  INV_X4 U4519 ( .A(n2762), .ZN(n2765) );
  INV_X4 U4520 ( .A(a[13]), .ZN(n2763) );
  OAI21_X4 U4521 ( .B1(n2765), .B2(n2764), .A(n3131), .ZN(n3121) );
  NAND3_X2 U4522 ( .A1(n2856), .A2(n2769), .A3(n2855), .ZN(n2851) );
  INV_X4 U4523 ( .A(n2856), .ZN(n2771) );
  XNOR2_X2 U4524 ( .A(n2775), .B(n2929), .ZN(n2777) );
  NAND2_X2 U4525 ( .A1(a[12]), .A2(n2034), .ZN(n2776) );
  INV_X4 U4526 ( .A(n2841), .ZN(n2842) );
  NAND4_X2 U4528 ( .A1(n2920), .A2(net330197), .A3(n2919), .A4(n1116), .ZN(
        n2873) );
  NAND2_X2 U4529 ( .A1(a[11]), .A2(net331343), .ZN(n3031) );
  INV_X4 U4530 ( .A(n3031), .ZN(n2848) );
  OAI21_X4 U4531 ( .B1(n3030), .B2(n2848), .A(n2792), .ZN(n2946) );
  XNOR2_X2 U4532 ( .A(n2801), .B(n2802), .ZN(n2804) );
  NAND2_X2 U4533 ( .A1(a[9]), .A2(net331323), .ZN(n2803) );
  NAND2_X2 U4534 ( .A1(n1407), .A2(n2803), .ZN(n2887) );
  INV_X4 U4535 ( .A(n2803), .ZN(n3014) );
  NAND2_X2 U4536 ( .A1(n3022), .A2(n2887), .ZN(n2805) );
  XNOR2_X2 U4537 ( .A(n2806), .B(n2805), .ZN(n2809) );
  INV_X4 U4538 ( .A(n2809), .ZN(n2807) );
  NAND2_X2 U4539 ( .A1(a[8]), .A2(n2037), .ZN(n2808) );
  INV_X4 U4540 ( .A(n2808), .ZN(n2810) );
  OAI21_X4 U4541 ( .B1(net331311), .B2(net330173), .A(n2813), .ZN(n2980) );
  NAND2_X2 U4542 ( .A1(product_in[14]), .A2(net331293), .ZN(n2816) );
  INV_X4 U4543 ( .A(n2816), .ZN(n2818) );
  NAND2_X2 U4544 ( .A1(n2827), .A2(n1732), .ZN(n2963) );
  NAND2_X2 U4545 ( .A1(a[9]), .A2(n2037), .ZN(n3002) );
  NAND2_X2 U4546 ( .A1(a[10]), .A2(net331323), .ZN(n2880) );
  INV_X4 U4547 ( .A(n2880), .ZN(n3015) );
  AND2_X2 U4548 ( .A1(net330043), .A2(net330042), .ZN(net330142) );
  NAND2_X2 U4549 ( .A1(n2842), .A2(n3031), .ZN(n2843) );
  NAND2_X2 U4550 ( .A1(a[12]), .A2(net331343), .ZN(n2876) );
  INV_X4 U4551 ( .A(n2876), .ZN(n2948) );
  NOR2_X4 U4552 ( .A1(n2850), .A2(n1736), .ZN(n2854) );
  INV_X4 U4553 ( .A(n2851), .ZN(n2853) );
  NAND3_X4 U4554 ( .A1(n2852), .A2(n2854), .A3(n2853), .ZN(n3129) );
  NAND2_X2 U4555 ( .A1(n1346), .A2(n2858), .ZN(n2859) );
  INV_X4 U4556 ( .A(n2863), .ZN(n2935) );
  XNOR2_X2 U4557 ( .A(n2936), .B(n2935), .ZN(n2865) );
  INV_X4 U4558 ( .A(n2867), .ZN(n2871) );
  NAND2_X2 U4559 ( .A1(a[13]), .A2(n2034), .ZN(n2869) );
  OAI21_X4 U4560 ( .B1(n2871), .B2(n2870), .A(n2869), .ZN(n2872) );
  XNOR2_X2 U4561 ( .A(n2875), .B(n1785), .ZN(n2877) );
  INV_X4 U4562 ( .A(n2877), .ZN(n2947) );
  NAND2_X2 U4563 ( .A1(a[11]), .A2(net331329), .ZN(net330089) );
  INV_X4 U4564 ( .A(net330089), .ZN(net330044) );
  INV_X4 U4565 ( .A(n3002), .ZN(n2881) );
  XNOR2_X2 U4566 ( .A(n2885), .B(n2884), .ZN(n3092) );
  NAND2_X2 U4567 ( .A1(a[8]), .A2(net331307), .ZN(n2983) );
  INV_X4 U4568 ( .A(n2983), .ZN(n2894) );
  XNOR2_X2 U4569 ( .A(n2895), .B(n2972), .ZN(n4365) );
  OAI21_X4 U4570 ( .B1(n2896), .B2(net331293), .A(net330067), .ZN(n2899) );
  INV_X4 U4571 ( .A(n2899), .ZN(n2897) );
  NAND2_X2 U4572 ( .A1(product_in[15]), .A2(net331293), .ZN(n2898) );
  INV_X4 U4573 ( .A(n2898), .ZN(n2900) );
  INV_X4 U4574 ( .A(n2906), .ZN(n3084) );
  INV_X4 U4575 ( .A(n2907), .ZN(n3675) );
  NAND2_X2 U4576 ( .A1(net331362), .A2(n3675), .ZN(n2993) );
  NAND2_X2 U4577 ( .A1(a[9]), .A2(net331307), .ZN(n2985) );
  INV_X4 U4578 ( .A(n2985), .ZN(n2997) );
  INV_X4 U4579 ( .A(n2888), .ZN(n2911) );
  NAND2_X2 U4580 ( .A1(net330040), .A2(net330088), .ZN(n2916) );
  NAND2_X2 U4581 ( .A1(a[12]), .A2(net331329), .ZN(net329972) );
  NAND2_X2 U4582 ( .A1(a[13]), .A2(net331343), .ZN(n2943) );
  INV_X4 U4583 ( .A(n2943), .ZN(n2950) );
  NAND4_X2 U4584 ( .A1(n1652), .A2(net330029), .A3(n2919), .A4(n1116), .ZN(
        n3039) );
  INV_X4 U4585 ( .A(n3042), .ZN(n2921) );
  NAND3_X4 U4586 ( .A1(n2923), .A2(net330021), .A3(n2924), .ZN(n3040) );
  NAND2_X2 U4587 ( .A1(n1661), .A2(n3040), .ZN(n2925) );
  NAND2_X2 U4588 ( .A1(a[14]), .A2(n2034), .ZN(n2939) );
  INV_X4 U4589 ( .A(a[15]), .ZN(n2927) );
  NAND3_X4 U4590 ( .A1(a[15]), .A2(n1340), .A3(net331349), .ZN(n3136) );
  OAI21_X4 U4591 ( .B1(n1340), .B2(n2928), .A(n3136), .ZN(n3122) );
  NAND3_X2 U4592 ( .A1(n2929), .A2(n3124), .A3(n3125), .ZN(n2930) );
  NAND2_X2 U4593 ( .A1(n2936), .A2(n2935), .ZN(n3132) );
  XNOR2_X2 U4594 ( .A(n2942), .B(n3045), .ZN(n2944) );
  INV_X4 U4595 ( .A(n2944), .ZN(n2949) );
  NAND2_X2 U4597 ( .A1(a[11]), .A2(net331323), .ZN(n3229) );
  INV_X4 U4598 ( .A(n3229), .ZN(n2954) );
  XNOR2_X2 U4599 ( .A(net329753), .B(n2952), .ZN(n2953) );
  NAND3_X2 U4600 ( .A1(n1646), .A2(a[10]), .A3(n2037), .ZN(n3410) );
  NAND2_X2 U4601 ( .A1(a[10]), .A2(n2037), .ZN(n2956) );
  INV_X4 U4602 ( .A(n2957), .ZN(n2961) );
  OAI21_X4 U4603 ( .B1(n2960), .B2(n2961), .A(n2959), .ZN(n3207) );
  OAI21_X4 U4604 ( .B1(n2966), .B2(n3205), .A(n3005), .ZN(n3093) );
  XNOR2_X2 U4605 ( .A(n2968), .B(n2995), .ZN(n2970) );
  INV_X4 U4606 ( .A(n2971), .ZN(n3669) );
  NAND2_X2 U4608 ( .A1(control[1]), .A2(n3670), .ZN(n2990) );
  XNOR2_X2 U4609 ( .A(n2978), .B(n2977), .ZN(n2984) );
  XNOR2_X2 U4610 ( .A(n2994), .B(n2985), .ZN(n2986) );
  XNOR2_X2 U4611 ( .A(n2986), .B(n2995), .ZN(n2988) );
  XNOR2_X2 U4612 ( .A(n3084), .B(n3082), .ZN(product_out[16]) );
  NAND3_X2 U4614 ( .A1(n3021), .A2(n3022), .A3(n3023), .ZN(n3024) );
  NAND2_X2 U4615 ( .A1(n3034), .A2(net329873), .ZN(n3037) );
  INV_X4 U4617 ( .A(net332761), .ZN(net329866) );
  AOI21_X4 U4618 ( .B1(n3033), .B2(n3032), .A(net329866), .ZN(n3035) );
  NAND3_X2 U4619 ( .A1(n3036), .A2(net329857), .A3(n3037), .ZN(n3060) );
  OAI21_X4 U4620 ( .B1(n3043), .B2(n3042), .A(n3041), .ZN(n3119) );
  OAI21_X4 U4621 ( .B1(n3046), .B2(n3122), .A(n3136), .ZN(n3051) );
  INV_X4 U4622 ( .A(n3048), .ZN(n3139) );
  XNOR2_X2 U4623 ( .A(n3140), .B(n3139), .ZN(n3050) );
  INV_X4 U4624 ( .A(n3056), .ZN(n3054) );
  NAND2_X2 U4625 ( .A1(n3133), .A2(n3051), .ZN(n3055) );
  NAND2_X2 U4626 ( .A1(a[15]), .A2(n2034), .ZN(n3052) );
  OAI21_X4 U4627 ( .B1(n3054), .B2(n3053), .A(n3052), .ZN(n3057) );
  XNOR2_X2 U4628 ( .A(n3060), .B(n1291), .ZN(n3062) );
  NAND2_X2 U4629 ( .A1(a[13]), .A2(net331329), .ZN(n3061) );
  INV_X4 U4630 ( .A(n3061), .ZN(n3064) );
  XNOR2_X2 U4631 ( .A(n3068), .B(n3217), .ZN(n3070) );
  NAND2_X2 U4632 ( .A1(a[11]), .A2(n2037), .ZN(n3069) );
  INV_X4 U4633 ( .A(n3069), .ZN(n3090) );
  INV_X4 U4634 ( .A(n3070), .ZN(n3089) );
  NAND2_X2 U4636 ( .A1(a[10]), .A2(net331307), .ZN(n3072) );
  INV_X4 U4637 ( .A(n3072), .ZN(n3196) );
  INV_X4 U4639 ( .A(n3182), .ZN(n3077) );
  OAI21_X4 U4640 ( .B1(n4417), .B2(net331293), .A(n3077), .ZN(n3080) );
  NAND2_X2 U4641 ( .A1(product_in[17]), .A2(net331293), .ZN(n3079) );
  NAND2_X2 U4642 ( .A1(n3078), .A2(n3079), .ZN(n3081) );
  INV_X4 U4643 ( .A(n3079), .ZN(n3183) );
  NAND2_X2 U4644 ( .A1(a[11]), .A2(net331307), .ZN(n3170) );
  INV_X4 U4645 ( .A(n3170), .ZN(n3297) );
  INV_X4 U4646 ( .A(n3209), .ZN(n3094) );
  INV_X4 U4647 ( .A(n3097), .ZN(n3100) );
  NAND3_X2 U4648 ( .A1(n3219), .A2(n3220), .A3(n3106), .ZN(n3158) );
  NAND2_X2 U4649 ( .A1(net329467), .A2(n4485), .ZN(n3275) );
  NAND3_X2 U4650 ( .A1(n3276), .A2(n1277), .A3(n3275), .ZN(n3108) );
  INV_X4 U4651 ( .A(n3239), .ZN(n3114) );
  AOI211_X4 U4652 ( .C1(n3115), .C2(net329737), .A(n3114), .B(n3113), .ZN(
        net329690) );
  NAND2_X2 U4653 ( .A1(a[15]), .A2(net331343), .ZN(n3152) );
  INV_X4 U4654 ( .A(n3152), .ZN(n3236) );
  NAND2_X2 U4655 ( .A1(a[16]), .A2(n2034), .ZN(n3146) );
  INV_X4 U4656 ( .A(n3123), .ZN(n3128) );
  INV_X4 U4657 ( .A(n3124), .ZN(n3127) );
  NAND2_X2 U4658 ( .A1(n3125), .A2(n3133), .ZN(n3126) );
  NOR3_X4 U4659 ( .A1(n3126), .A2(n3127), .A3(n3128), .ZN(n3130) );
  NAND2_X2 U4660 ( .A1(n3140), .A2(n3139), .ZN(n3248) );
  INV_X4 U4661 ( .A(a[17]), .ZN(n3142) );
  XNOR2_X2 U4662 ( .A(n3144), .B(n3251), .ZN(n3147) );
  NAND2_X2 U4663 ( .A1(n3146), .A2(n3145), .ZN(n3148) );
  NAND3_X2 U4664 ( .A1(n3147), .A2(a[16]), .A3(n2034), .ZN(n3354) );
  XNOR2_X2 U4665 ( .A(n3151), .B(n1447), .ZN(n3149) );
  XNOR2_X2 U4666 ( .A(n3151), .B(n1447), .ZN(n3235) );
  XNOR2_X2 U4667 ( .A(n3154), .B(n1390), .ZN(n3225) );
  NAND2_X2 U4668 ( .A1(a[13]), .A2(net331323), .ZN(n3156) );
  INV_X4 U4669 ( .A(n3156), .ZN(n3226) );
  NAND2_X2 U4670 ( .A1(a[12]), .A2(n2037), .ZN(n3222) );
  INV_X4 U4671 ( .A(n3222), .ZN(n3160) );
  INV_X4 U4672 ( .A(n3168), .ZN(n3161) );
  XNOR2_X2 U4673 ( .A(n3163), .B(n3162), .ZN(n3319) );
  NOR3_X4 U4674 ( .A1(n1662), .A2(n3164), .A3(n2024), .ZN(n3165) );
  XNOR2_X2 U4675 ( .A(n3169), .B(n3168), .ZN(n3295) );
  NAND2_X2 U4676 ( .A1(n3320), .A2(n3319), .ZN(n3202) );
  NAND2_X2 U4677 ( .A1(product_in[18]), .A2(net331293), .ZN(n3188) );
  INV_X4 U4678 ( .A(n3174), .ZN(n3496) );
  INV_X4 U4679 ( .A(n3191), .ZN(n3309) );
  INV_X4 U4680 ( .A(n3188), .ZN(n3190) );
  NAND2_X2 U4681 ( .A1(n3190), .A2(n3189), .ZN(n3489) );
  INV_X4 U4682 ( .A(n3489), .ZN(n3495) );
  XNOR2_X2 U4683 ( .A(n3199), .B(n1675), .ZN(n3201) );
  INV_X4 U4684 ( .A(n3202), .ZN(n3203) );
  NAND2_X2 U4685 ( .A1(a[12]), .A2(net331307), .ZN(n3291) );
  INV_X4 U4686 ( .A(n3291), .ZN(n3290) );
  INV_X4 U4687 ( .A(n3329), .ZN(n3224) );
  OAI211_X2 U4688 ( .C1(n3232), .C2(n3231), .A(n1141), .B(n1482), .ZN(n3233)
         );
  NAND2_X2 U4689 ( .A1(a[16]), .A2(net331343), .ZN(n3272) );
  INV_X4 U4690 ( .A(n3272), .ZN(n3269) );
  NAND2_X2 U4691 ( .A1(a[17]), .A2(n2034), .ZN(n3265) );
  INV_X4 U4692 ( .A(n3251), .ZN(n3252) );
  NAND2_X2 U4693 ( .A1(a[18]), .A2(net331349), .ZN(n3258) );
  INV_X4 U4694 ( .A(n3258), .ZN(n3360) );
  INV_X4 U4695 ( .A(n3259), .ZN(n3359) );
  XNOR2_X2 U4696 ( .A(n3360), .B(n3359), .ZN(n3261) );
  NAND2_X2 U4697 ( .A1(n3260), .A2(n3261), .ZN(n3264) );
  INV_X4 U4698 ( .A(n3261), .ZN(n3263) );
  NAND3_X4 U4699 ( .A1(n3267), .A2(a[17]), .A3(n2034), .ZN(n3445) );
  NAND2_X2 U4700 ( .A1(n3440), .A2(n3445), .ZN(n3353) );
  XNOR2_X2 U4701 ( .A(n3268), .B(n3353), .ZN(n3270) );
  NAND2_X2 U4703 ( .A1(a[15]), .A2(net331329), .ZN(net329340) );
  XNOR2_X2 U4704 ( .A(n3424), .B(net329352), .ZN(n3274) );
  NAND2_X2 U4705 ( .A1(a[14]), .A2(net331323), .ZN(n3423) );
  INV_X4 U4706 ( .A(n3423), .ZN(n3281) );
  XNOR2_X2 U4707 ( .A(n3279), .B(net329545), .ZN(n3280) );
  XNOR2_X2 U4708 ( .A(n3283), .B(n3282), .ZN(n3285) );
  NAND2_X2 U4709 ( .A1(a[13]), .A2(n2037), .ZN(n3284) );
  INV_X4 U4710 ( .A(n3284), .ZN(n3287) );
  INV_X4 U4711 ( .A(n1653), .ZN(n3286) );
  XNOR2_X2 U4712 ( .A(n4467), .B(n3288), .ZN(n3292) );
  NOR2_X4 U4713 ( .A1(n3293), .A2(net331295), .ZN(n3294) );
  NAND2_X2 U4714 ( .A1(n4018), .A2(n3294), .ZN(n3305) );
  NAND2_X2 U4715 ( .A1(n3300), .A2(net328035), .ZN(n3301) );
  NAND3_X2 U4716 ( .A1(n3305), .A2(n3304), .A3(n3303), .ZN(n3307) );
  NAND2_X2 U4717 ( .A1(product_in[19]), .A2(net331293), .ZN(n3493) );
  NAND2_X2 U4718 ( .A1(n3306), .A2(n3493), .ZN(n3310) );
  INV_X4 U4719 ( .A(n3493), .ZN(n3494) );
  NAND2_X2 U4721 ( .A1(n3309), .A2(n3489), .ZN(n3311) );
  INV_X4 U4722 ( .A(n3316), .ZN(n3317) );
  NAND3_X4 U4723 ( .A1(n3323), .A2(n3325), .A3(n3324), .ZN(n3504) );
  NAND2_X2 U4724 ( .A1(a[14]), .A2(n2037), .ZN(n3589) );
  INV_X4 U4725 ( .A(n3589), .ZN(n3416) );
  NAND3_X2 U4726 ( .A1(n1849), .A2(n3334), .A3(n3333), .ZN(n3336) );
  NAND2_X2 U4727 ( .A1(n3345), .A2(net329456), .ZN(n3343) );
  OAI21_X4 U4728 ( .B1(n3342), .B2(n3343), .A(n3341), .ZN(n3434) );
  INV_X4 U4729 ( .A(n3434), .ZN(n3526) );
  INV_X4 U4730 ( .A(n3353), .ZN(n3356) );
  NAND2_X2 U4731 ( .A1(n3355), .A2(n3354), .ZN(n3439) );
  NAND2_X2 U4732 ( .A1(a[18]), .A2(n2034), .ZN(n3369) );
  NAND2_X2 U4733 ( .A1(n3360), .A2(n3359), .ZN(n3362) );
  INV_X4 U4734 ( .A(n3365), .ZN(n3366) );
  INV_X4 U4735 ( .A(n3370), .ZN(n3368) );
  XNOR2_X2 U4736 ( .A(n3372), .B(n3441), .ZN(n3375) );
  NAND2_X2 U4737 ( .A1(a[17]), .A2(net331343), .ZN(n3374) );
  NAND2_X2 U4738 ( .A1(n3373), .A2(n3374), .ZN(n3618) );
  INV_X4 U4739 ( .A(n3374), .ZN(n3376) );
  XNOR2_X2 U4740 ( .A(n3377), .B(n3430), .ZN(net329410) );
  NAND2_X2 U4741 ( .A1(a[15]), .A2(net331323), .ZN(net329397) );
  INV_X4 U4742 ( .A(net329397), .ZN(net329404) );
  XNOR2_X2 U4743 ( .A(net329395), .B(n3384), .ZN(n3517) );
  XNOR2_X2 U4744 ( .A(n4443), .B(n3385), .ZN(n3590) );
  NAND2_X2 U4745 ( .A1(a[13]), .A2(net331307), .ZN(n3389) );
  INV_X4 U4746 ( .A(n3389), .ZN(n3391) );
  INV_X4 U4747 ( .A(n3500), .ZN(n3394) );
  OAI21_X4 U4748 ( .B1(n1364), .B2(net331295), .A(n3394), .ZN(n4211) );
  XNOR2_X2 U4750 ( .A(n3395), .B(n1337), .ZN(n3400) );
  NAND3_X2 U4751 ( .A1(n3398), .A2(n3400), .A3(n3399), .ZN(n3401) );
  NAND2_X2 U4752 ( .A1(n1337), .A2(n4211), .ZN(n3502) );
  NAND2_X2 U4753 ( .A1(a[15]), .A2(n2037), .ZN(n3474) );
  INV_X4 U4754 ( .A(n3474), .ZN(n3473) );
  XNOR2_X2 U4755 ( .A(n3425), .B(n3424), .ZN(n3427) );
  NAND3_X2 U4756 ( .A1(n3519), .A2(n1138), .A3(n3517), .ZN(n3684) );
  NAND2_X2 U4757 ( .A1(a[16]), .A2(net331323), .ZN(n3470) );
  INV_X4 U4758 ( .A(n3470), .ZN(n3521) );
  NAND2_X2 U4759 ( .A1(a[17]), .A2(net331329), .ZN(n3468) );
  INV_X4 U4760 ( .A(n3468), .ZN(n3523) );
  NAND2_X2 U4761 ( .A1(n3430), .A2(n1649), .ZN(n3438) );
  NAND3_X2 U4762 ( .A1(n3623), .A2(n1788), .A3(n1193), .ZN(n3437) );
  NAND2_X2 U4763 ( .A1(a[18]), .A2(net331343), .ZN(n3466) );
  NAND2_X2 U4764 ( .A1(n3440), .A2(n3439), .ZN(n3442) );
  AOI21_X4 U4765 ( .B1(n3445), .B2(n3442), .A(n3441), .ZN(n3452) );
  INV_X4 U4766 ( .A(n3444), .ZN(n3446) );
  AOI21_X4 U4767 ( .B1(n3452), .B2(n3451), .A(n3450), .ZN(n3533) );
  NAND2_X2 U4768 ( .A1(a[19]), .A2(n2035), .ZN(n3461) );
  OAI21_X4 U4769 ( .B1(n3455), .B2(n3454), .A(n3453), .ZN(n3637) );
  NAND2_X2 U4770 ( .A1(a[20]), .A2(net331349), .ZN(n3456) );
  INV_X4 U4771 ( .A(n3456), .ZN(n3536) );
  INV_X4 U4772 ( .A(n3457), .ZN(n3535) );
  XNOR2_X2 U4773 ( .A(n3536), .B(n3535), .ZN(n3459) );
  NAND2_X2 U4774 ( .A1(n3458), .A2(n3459), .ZN(n3460) );
  INV_X4 U4775 ( .A(n3459), .ZN(n3638) );
  NAND2_X2 U4776 ( .A1(n3460), .A2(n3537), .ZN(n3462) );
  NAND2_X2 U4777 ( .A1(n3461), .A2(n3462), .ZN(n3464) );
  INV_X4 U4778 ( .A(n3462), .ZN(n3463) );
  NAND3_X4 U4779 ( .A1(n3463), .A2(a[19]), .A3(n2035), .ZN(n3531) );
  INV_X4 U4780 ( .A(n3532), .ZN(n3465) );
  XNOR2_X2 U4781 ( .A(n3533), .B(n3465), .ZN(net329295) );
  XNOR2_X2 U4782 ( .A(n3477), .B(n3476), .ZN(n3479) );
  NAND2_X2 U4783 ( .A1(a[14]), .A2(net331305), .ZN(n3478) );
  INV_X4 U4784 ( .A(n3478), .ZN(n3481) );
  INV_X4 U4785 ( .A(n4194), .ZN(n3486) );
  NAND2_X2 U4786 ( .A1(n4195), .A2(net328035), .ZN(n3485) );
  OAI21_X4 U4787 ( .B1(n3486), .B2(net331363), .A(n3485), .ZN(n3487) );
  AOI21_X4 U4788 ( .B1(product_in[21]), .B2(net331293), .A(n3487), .ZN(n4222)
         );
  NAND2_X2 U4789 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  OAI211_X2 U4790 ( .C1(n1337), .C2(n3500), .A(n3499), .B(n3498), .ZN(n4215)
         );
  NAND3_X4 U4791 ( .A1(n3504), .A2(n1879), .A3(n1907), .ZN(n3730) );
  NOR2_X4 U4792 ( .A1(n3510), .A2(n3763), .ZN(n3511) );
  OAI21_X4 U4793 ( .B1(n3513), .B2(n3512), .A(n3511), .ZN(n3679) );
  NAND3_X2 U4794 ( .A1(n3519), .A2(n3518), .A3(n3517), .ZN(n3520) );
  INV_X4 U4795 ( .A(n3554), .ZN(n3560) );
  OAI21_X4 U4796 ( .B1(net329225), .B2(net333991), .A(net328741), .ZN(n3553)
         );
  INV_X4 U4797 ( .A(n3527), .ZN(n3528) );
  NAND2_X2 U4798 ( .A1(n3528), .A2(n3618), .ZN(n3529) );
  NAND2_X2 U4799 ( .A1(a[19]), .A2(net331343), .ZN(n3549) );
  OAI21_X4 U4800 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3534) );
  NAND2_X2 U4801 ( .A1(a[20]), .A2(n2034), .ZN(n3544) );
  NAND2_X2 U4802 ( .A1(n3536), .A2(n3535), .ZN(n3632) );
  NAND2_X2 U4803 ( .A1(n3537), .A2(n3632), .ZN(n3542) );
  INV_X4 U4804 ( .A(n3539), .ZN(n3540) );
  NAND2_X2 U4805 ( .A1(n3541), .A2(n3631), .ZN(n3635) );
  XNOR2_X2 U4806 ( .A(n3542), .B(n3635), .ZN(n3545) );
  NAND2_X2 U4807 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  NAND3_X2 U4808 ( .A1(a[20]), .A2(n3545), .A3(n2034), .ZN(n3627) );
  NAND2_X2 U4809 ( .A1(n3625), .A2(n3708), .ZN(n3551) );
  NAND2_X2 U4810 ( .A1(a[18]), .A2(net331329), .ZN(net329194) );
  NAND2_X2 U4811 ( .A1(n3606), .A2(n3687), .ZN(n3610) );
  NAND2_X2 U4813 ( .A1(a[15]), .A2(net331305), .ZN(n3727) );
  INV_X4 U4814 ( .A(n3727), .ZN(n3566) );
  NAND2_X2 U4815 ( .A1(product_in[22]), .A2(net331295), .ZN(n3571) );
  XNOR2_X2 U4816 ( .A(n3572), .B(n3571), .ZN(n3568) );
  INV_X4 U4817 ( .A(n3568), .ZN(n4221) );
  NAND2_X2 U4818 ( .A1(n1360), .A2(n3840), .ZN(n3937) );
  INV_X4 U4819 ( .A(n3571), .ZN(n3573) );
  NAND2_X2 U4820 ( .A1(n3573), .A2(n3572), .ZN(n4230) );
  OAI21_X4 U4821 ( .B1(n3574), .B2(n4209), .A(n4230), .ZN(n3940) );
  OAI21_X4 U4822 ( .B1(n3576), .B2(n3937), .A(n3575), .ZN(n3577) );
  NAND3_X2 U4823 ( .A1(n3592), .A2(n3591), .A3(n3593), .ZN(n3595) );
  NAND2_X2 U4824 ( .A1(n1735), .A2(n1771), .ZN(n3603) );
  NAND2_X2 U4825 ( .A1(a[17]), .A2(n2037), .ZN(n3658) );
  INV_X4 U4826 ( .A(n3658), .ZN(n3657) );
  NOR2_X4 U4827 ( .A1(n3607), .A2(n3611), .ZN(n3608) );
  NAND2_X2 U4828 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  NAND2_X2 U4829 ( .A1(a[19]), .A2(net331329), .ZN(n3655) );
  INV_X4 U4830 ( .A(n3655), .ZN(n3652) );
  INV_X4 U4831 ( .A(n3619), .ZN(n3620) );
  AOI21_X4 U4832 ( .B1(net329112), .B2(n3621), .A(n3620), .ZN(n3626) );
  NAND3_X4 U4833 ( .A1(n3624), .A2(n3626), .A3(n3625), .ZN(n3706) );
  NAND2_X2 U4834 ( .A1(a[20]), .A2(net331343), .ZN(n3649) );
  INV_X4 U4835 ( .A(n3649), .ZN(n3646) );
  OAI21_X4 U4836 ( .B1(n1298), .B2(n3628), .A(n1144), .ZN(n3694) );
  INV_X4 U4837 ( .A(n3630), .ZN(n3695) );
  XNOR2_X2 U4838 ( .A(n1213), .B(n3695), .ZN(n3643) );
  INV_X4 U4839 ( .A(n3643), .ZN(n3641) );
  INV_X4 U4840 ( .A(n3632), .ZN(n3633) );
  NOR2_X4 U4841 ( .A1(n3634), .A2(n3633), .ZN(n3640) );
  INV_X4 U4842 ( .A(n3635), .ZN(n3636) );
  NAND3_X2 U4843 ( .A1(n3637), .A2(n3638), .A3(n3636), .ZN(n3639) );
  NAND2_X2 U4844 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  NAND3_X4 U4845 ( .A1(n1218), .A2(a[21]), .A3(n2034), .ZN(n3775) );
  XNOR2_X2 U4846 ( .A(n1658), .B(n3769), .ZN(n3647) );
  NAND2_X2 U4847 ( .A1(n3646), .A2(n3647), .ZN(n3707) );
  INV_X4 U4848 ( .A(n3647), .ZN(n3648) );
  XNOR2_X2 U4849 ( .A(n3650), .B(n3705), .ZN(n3651) );
  NAND2_X2 U4850 ( .A1(a[16]), .A2(net331305), .ZN(n3661) );
  INV_X4 U4851 ( .A(n3661), .ZN(n3721) );
  NAND2_X2 U4852 ( .A1(product_in[23]), .A2(net331295), .ZN(n3666) );
  INV_X4 U4853 ( .A(n4229), .ZN(n3664) );
  OAI21_X4 U4854 ( .B1(n1121), .B2(net331295), .A(n3664), .ZN(n4225) );
  INV_X4 U4855 ( .A(net329055), .ZN(net329052) );
  INV_X4 U4856 ( .A(n3666), .ZN(n3667) );
  OAI21_X4 U4857 ( .B1(n3668), .B2(net329052), .A(n3667), .ZN(n4228) );
  NAND2_X2 U4858 ( .A1(net328035), .A2(n3675), .ZN(n3676) );
  OAI21_X4 U4859 ( .B1(n3677), .B2(control[0]), .A(n3676), .ZN(n3745) );
  NAND2_X2 U4860 ( .A1(product_in[24]), .A2(net331295), .ZN(n4232) );
  INV_X4 U4861 ( .A(n4232), .ZN(n3746) );
  XNOR2_X2 U4862 ( .A(n4233), .B(n3746), .ZN(n3724) );
  NAND2_X2 U4863 ( .A1(a[17]), .A2(net331305), .ZN(n3718) );
  INV_X4 U4864 ( .A(n3718), .ZN(n3813) );
  INV_X4 U4865 ( .A(net328980), .ZN(net328982) );
  INV_X4 U4866 ( .A(n3683), .ZN(n3685) );
  NAND2_X2 U4867 ( .A1(n1688), .A2(n3471), .ZN(n3691) );
  INV_X4 U4868 ( .A(n3687), .ZN(n3689) );
  NOR2_X4 U4869 ( .A1(n3688), .A2(n3689), .ZN(n3690) );
  OAI21_X4 U4870 ( .B1(net329017), .B2(n1392), .A(n1388), .ZN(n3693) );
  NAND3_X4 U4871 ( .A1(net329015), .A2(n3693), .A3(net329014), .ZN(n3767) );
  INV_X4 U4872 ( .A(a[22]), .ZN(net329000) );
  NAND2_X2 U4873 ( .A1(n1213), .A2(n3695), .ZN(n3697) );
  INV_X4 U4874 ( .A(a[23]), .ZN(net329006) );
  OAI21_X4 U4875 ( .B1(n1342), .B2(n3699), .A(n3779), .ZN(n3780) );
  INV_X4 U4876 ( .A(n3780), .ZN(n3700) );
  OAI21_X4 U4877 ( .B1(n1172), .B2(net329000), .A(n3701), .ZN(n3770) );
  NAND2_X2 U4878 ( .A1(a[21]), .A2(net331343), .ZN(n3795) );
  XNOR2_X2 U4879 ( .A(n3796), .B(n3795), .ZN(n3703) );
  XNOR2_X2 U4880 ( .A(n3797), .B(n3703), .ZN(n3710) );
  NAND3_X4 U4881 ( .A1(n3706), .A2(n3707), .A3(n1237), .ZN(n3709) );
  NAND3_X4 U4882 ( .A1(n3709), .A2(n3710), .A3(n1296), .ZN(n3889) );
  NAND2_X2 U4883 ( .A1(a[20]), .A2(net331329), .ZN(n3803) );
  INV_X4 U4884 ( .A(n3803), .ZN(n3713) );
  NAND3_X4 U4885 ( .A1(n3712), .A2(n1414), .A3(n3713), .ZN(net328616) );
  NAND2_X2 U4886 ( .A1(a[18]), .A2(n2037), .ZN(n3852) );
  INV_X4 U4887 ( .A(n3852), .ZN(n3755) );
  XNOR2_X2 U4888 ( .A(n3716), .B(n3715), .ZN(n3812) );
  INV_X4 U4889 ( .A(n3812), .ZN(n3717) );
  NAND2_X2 U4890 ( .A1(n3960), .A2(net331299), .ZN(n3722) );
  NOR2_X4 U4891 ( .A1(n3753), .A2(n3722), .ZN(n3723) );
  NOR2_X4 U4892 ( .A1(n3724), .A2(n3723), .ZN(n3737) );
  NOR2_X4 U4893 ( .A1(n3752), .A2(n3725), .ZN(n3733) );
  OAI21_X4 U4895 ( .B1(n3751), .B2(n3743), .A(n4228), .ZN(n3744) );
  XNOR2_X2 U4896 ( .A(n3744), .B(n1644), .ZN(product_out[24]) );
  NAND2_X2 U4898 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  OAI21_X4 U4899 ( .B1(n3751), .B2(n3750), .A(n3749), .ZN(n3835) );
  NAND3_X2 U4900 ( .A1(net328936), .A2(net328937), .A3(n3755), .ZN(n3757) );
  NOR3_X4 U4901 ( .A1(n3761), .A2(n1955), .A3(n3760), .ZN(n3762) );
  INV_X4 U4902 ( .A(n3766), .ZN(n3947) );
  NAND2_X2 U4903 ( .A1(net328737), .A2(net328616), .ZN(net328604) );
  NAND2_X2 U4905 ( .A1(a[21]), .A2(net331329), .ZN(n3904) );
  INV_X4 U4906 ( .A(n3904), .ZN(n3800) );
  NAND2_X2 U4907 ( .A1(a[22]), .A2(net331343), .ZN(n3793) );
  INV_X4 U4908 ( .A(n3769), .ZN(n3771) );
  INV_X4 U4909 ( .A(n3778), .ZN(n3862) );
  XNOR2_X2 U4910 ( .A(n1214), .B(n3862), .ZN(n3784) );
  INV_X4 U4911 ( .A(n3784), .ZN(n3782) );
  OAI21_X4 U4912 ( .B1(n3781), .B2(n3780), .A(n3779), .ZN(n3783) );
  NAND2_X2 U4913 ( .A1(n3785), .A2(n3784), .ZN(n3789) );
  INV_X4 U4914 ( .A(n3789), .ZN(n3787) );
  NAND2_X2 U4915 ( .A1(a[23]), .A2(n2034), .ZN(n3786) );
  OAI21_X4 U4916 ( .B1(n3788), .B2(n3787), .A(n3786), .ZN(n3790) );
  NAND2_X2 U4917 ( .A1(n3790), .A2(n3876), .ZN(n3877) );
  INV_X4 U4918 ( .A(n3877), .ZN(n3791) );
  XNOR2_X2 U4919 ( .A(n3878), .B(n3791), .ZN(n3794) );
  NAND2_X2 U4920 ( .A1(n3793), .A2(n3792), .ZN(n3887) );
  NAND3_X2 U4921 ( .A1(n3794), .A2(a[22]), .A3(net331341), .ZN(n3884) );
  NAND2_X2 U4922 ( .A1(n3887), .A2(n3884), .ZN(n3976) );
  INV_X4 U4923 ( .A(n3795), .ZN(n3799) );
  NAND2_X2 U4924 ( .A1(n3799), .A2(n3798), .ZN(n3885) );
  XNOR2_X2 U4926 ( .A(n3807), .B(n3806), .ZN(n3809) );
  INV_X4 U4927 ( .A(net328790), .ZN(net328853) );
  NAND2_X2 U4928 ( .A1(n3813), .A2(n1366), .ZN(n4090) );
  OAI21_X4 U4930 ( .B1(n4417), .B2(net331363), .A(n3819), .ZN(n3928) );
  INV_X4 U4931 ( .A(n3928), .ZN(n3821) );
  NAND2_X2 U4932 ( .A1(product_in[25]), .A2(net331295), .ZN(n3825) );
  NAND2_X2 U4933 ( .A1(n3821), .A2(n3825), .ZN(n4241) );
  INV_X4 U4934 ( .A(n4241), .ZN(n3833) );
  OAI211_X2 U4935 ( .C1(n3824), .C2(n3823), .A(n3822), .B(n3833), .ZN(n3834)
         );
  INV_X4 U4936 ( .A(n3825), .ZN(n3930) );
  NAND2_X2 U4937 ( .A1(n3930), .A2(n3928), .ZN(n4238) );
  INV_X4 U4938 ( .A(n3828), .ZN(n3849) );
  NAND2_X2 U4939 ( .A1(n4090), .A2(n1630), .ZN(n3847) );
  NAND2_X2 U4940 ( .A1(n3829), .A2(n3847), .ZN(n3830) );
  NAND3_X2 U4941 ( .A1(n3831), .A2(n3830), .A3(net331299), .ZN(n3832) );
  NAND2_X2 U4942 ( .A1(n3838), .A2(n3933), .ZN(n3839) );
  INV_X4 U4943 ( .A(n3839), .ZN(n4125) );
  OAI21_X4 U4944 ( .B1(n1125), .B2(n3841), .A(n1725), .ZN(n3843) );
  NAND2_X2 U4945 ( .A1(n3930), .A2(n3928), .ZN(n3929) );
  XNOR2_X2 U4946 ( .A(n3845), .B(n3950), .ZN(n3846) );
  INV_X4 U4947 ( .A(n3855), .ZN(n4013) );
  NAND2_X2 U4948 ( .A1(net328791), .A2(n3859), .ZN(n3861) );
  NAND3_X2 U4949 ( .A1(n3861), .A2(net328588), .A3(n3860), .ZN(n3909) );
  NAND2_X2 U4950 ( .A1(n1214), .A2(n3862), .ZN(n3864) );
  NAND2_X2 U4951 ( .A1(n3866), .A2(n3867), .ZN(n3869) );
  INV_X4 U4952 ( .A(n3867), .ZN(n3868) );
  NAND2_X2 U4953 ( .A1(n3869), .A2(n3982), .ZN(n3983) );
  INV_X4 U4954 ( .A(n3983), .ZN(n3870) );
  XNOR2_X2 U4955 ( .A(n3984), .B(n3870), .ZN(n3873) );
  INV_X4 U4956 ( .A(n3873), .ZN(n3871) );
  NAND2_X2 U4957 ( .A1(a[24]), .A2(n2034), .ZN(n3872) );
  INV_X4 U4958 ( .A(n3872), .ZN(n3874) );
  XNOR2_X2 U4959 ( .A(n1175), .B(n3996), .ZN(n3881) );
  NAND2_X2 U4960 ( .A1(a[23]), .A2(net331343), .ZN(n3880) );
  INV_X4 U4961 ( .A(n3880), .ZN(n3882) );
  INV_X4 U4962 ( .A(n3884), .ZN(n3974) );
  INV_X4 U4963 ( .A(n3885), .ZN(n3886) );
  INV_X4 U4964 ( .A(n3887), .ZN(n3888) );
  AOI21_X4 U4965 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n3891) );
  NAND2_X2 U4966 ( .A1(a[22]), .A2(net331329), .ZN(n3892) );
  INV_X4 U4967 ( .A(n3892), .ZN(n4006) );
  NAND2_X2 U4968 ( .A1(a[21]), .A2(net331323), .ZN(n4009) );
  NAND3_X2 U4969 ( .A1(a[21]), .A2(net328607), .A3(net331323), .ZN(n3895) );
  XNOR2_X2 U4970 ( .A(n3909), .B(n3908), .ZN(n3912) );
  NAND2_X2 U4971 ( .A1(a[20]), .A2(n2037), .ZN(n3911) );
  INV_X4 U4972 ( .A(n3911), .ZN(n3913) );
  NAND2_X2 U4973 ( .A1(n3913), .A2(n3912), .ZN(n4082) );
  NAND2_X2 U4974 ( .A1(a[19]), .A2(net331305), .ZN(n3954) );
  INV_X4 U4975 ( .A(n3954), .ZN(n3917) );
  INV_X4 U4976 ( .A(n3955), .ZN(n3916) );
  NAND2_X2 U4977 ( .A1(product_in[26]), .A2(net331295), .ZN(n3943) );
  NAND2_X2 U4978 ( .A1(n3920), .A2(net331613), .ZN(n3921) );
  XNOR2_X2 U4979 ( .A(n1647), .B(n3943), .ZN(n4243) );
  INV_X4 U4980 ( .A(n3927), .ZN(n4239) );
  INV_X4 U4981 ( .A(n3929), .ZN(n4032) );
  NAND2_X2 U4982 ( .A1(n4239), .A2(n3930), .ZN(n3931) );
  INV_X4 U4983 ( .A(n3931), .ZN(n4031) );
  NOR3_X4 U4984 ( .A1(n1341), .A2(n4032), .A3(n4031), .ZN(n3935) );
  AOI21_X4 U4985 ( .B1(n3935), .B2(n4034), .A(n3934), .ZN(n3946) );
  INV_X4 U4986 ( .A(n3937), .ZN(n3939) );
  NAND3_X4 U4987 ( .A1(n3938), .A2(n3939), .A3(n1404), .ZN(n3942) );
  INV_X4 U4988 ( .A(n3943), .ZN(n3944) );
  XNOR2_X2 U4989 ( .A(n3949), .B(n3948), .ZN(n3951) );
  XNOR2_X2 U4990 ( .A(n3951), .B(n3950), .ZN(n3952) );
  INV_X4 U4991 ( .A(n3958), .ZN(n3968) );
  NAND2_X2 U4992 ( .A1(a[21]), .A2(n2037), .ZN(net328404) );
  OAI21_X4 U4993 ( .B1(n3977), .B2(n4389), .A(n3975), .ZN(n4041) );
  NAND2_X2 U4994 ( .A1(n3979), .A2(n3978), .ZN(n4042) );
  NAND2_X2 U4995 ( .A1(n4041), .A2(n4042), .ZN(n4002) );
  INV_X4 U4996 ( .A(n3980), .ZN(n4046) );
  INV_X4 U4997 ( .A(n3981), .ZN(n4045) );
  XNOR2_X2 U4998 ( .A(n4046), .B(n4045), .ZN(n3987) );
  INV_X4 U4999 ( .A(n3987), .ZN(n3985) );
  OAI21_X4 U5000 ( .B1(n3984), .B2(n3983), .A(n3982), .ZN(n3986) );
  NAND2_X2 U5001 ( .A1(a[25]), .A2(n2035), .ZN(n3989) );
  OAI21_X4 U5002 ( .B1(n3991), .B2(n3990), .A(n3989), .ZN(n3993) );
  INV_X4 U5003 ( .A(n1175), .ZN(n3997) );
  OAI21_X4 U5004 ( .B1(n3997), .B2(n1198), .A(n3995), .ZN(n4154) );
  NAND2_X2 U5005 ( .A1(a[24]), .A2(net331343), .ZN(n3998) );
  NAND2_X2 U5006 ( .A1(n3998), .A2(n1391), .ZN(n4043) );
  INV_X4 U5007 ( .A(n3998), .ZN(n4000) );
  XNOR2_X2 U5009 ( .A(n4002), .B(n4001), .ZN(n4004) );
  NAND2_X2 U5010 ( .A1(a[23]), .A2(net331329), .ZN(n4003) );
  NOR2_X4 U5011 ( .A1(net328605), .A2(net328606), .ZN(n4008) );
  INV_X4 U5012 ( .A(net328604), .ZN(net328602) );
  NAND3_X4 U5013 ( .A1(net328603), .A2(net328602), .A3(net328601), .ZN(n4007)
         );
  NAND3_X4 U5014 ( .A1(n4008), .A2(n4007), .A3(net328599), .ZN(n4072) );
  INV_X4 U5015 ( .A(n4009), .ZN(n4010) );
  NAND2_X2 U5016 ( .A1(a[20]), .A2(net331305), .ZN(net328528) );
  NOR2_X4 U5017 ( .A1(n4014), .A2(n1642), .ZN(n4016) );
  OAI21_X4 U5018 ( .B1(n4016), .B2(n4015), .A(n4422), .ZN(net328527) );
  XNOR2_X2 U5019 ( .A(n4017), .B(n4454), .ZN(n4029) );
  NOR2_X4 U5020 ( .A1(n4019), .A2(n4018), .ZN(n4021) );
  XNOR2_X2 U5021 ( .A(n4021), .B(n1245), .ZN(n4026) );
  NAND2_X2 U5022 ( .A1(product_in[27]), .A2(net331295), .ZN(n4118) );
  INV_X4 U5023 ( .A(n4118), .ZN(n4028) );
  XNOR2_X2 U5024 ( .A(n4030), .B(n1742), .ZN(product_out[27]) );
  NOR3_X4 U5025 ( .A1(n1341), .A2(n4032), .A3(n4031), .ZN(n4035) );
  AOI21_X4 U5026 ( .B1(n4035), .B2(n4034), .A(n4033), .ZN(n4040) );
  INV_X4 U5027 ( .A(net328533), .ZN(net328272) );
  AOI21_X4 U5028 ( .B1(n4037), .B2(net333918), .A(net328272), .ZN(n4038) );
  AOI21_X4 U5029 ( .B1(n4040), .B2(n4039), .A(n4038), .ZN(n4116) );
  NAND2_X2 U5030 ( .A1(a[22]), .A2(n2037), .ZN(n4080) );
  INV_X4 U5031 ( .A(n4080), .ZN(n4256) );
  INV_X4 U5032 ( .A(net328392), .ZN(net328389) );
  INV_X4 U5033 ( .A(n4154), .ZN(n4044) );
  NAND2_X2 U5034 ( .A1(n4046), .A2(n4045), .ZN(n4048) );
  INV_X4 U5035 ( .A(n4049), .ZN(n4162) );
  INV_X4 U5036 ( .A(n4051), .ZN(n4052) );
  NAND2_X2 U5037 ( .A1(n4053), .A2(n4160), .ZN(n4161) );
  NAND2_X2 U5038 ( .A1(a[26]), .A2(n2034), .ZN(n4055) );
  NAND2_X2 U5039 ( .A1(n4054), .A2(n4055), .ZN(n4058) );
  INV_X4 U5040 ( .A(n4055), .ZN(n4057) );
  NAND2_X2 U5041 ( .A1(a[25]), .A2(net331343), .ZN(n4061) );
  INV_X4 U5042 ( .A(n4061), .ZN(n4064) );
  NAND2_X2 U5043 ( .A1(a[24]), .A2(net331329), .ZN(n4068) );
  INV_X4 U5044 ( .A(n4068), .ZN(n4070) );
  XNOR2_X2 U5045 ( .A(n4074), .B(n4073), .ZN(n4077) );
  XNOR2_X2 U5046 ( .A(n4079), .B(n4452), .ZN(n4255) );
  XNOR2_X2 U5047 ( .A(net331520), .B(n4089), .ZN(net328158) );
  NAND2_X2 U5048 ( .A1(n4093), .A2(n4092), .ZN(n4297) );
  INV_X4 U5049 ( .A(n4296), .ZN(n4095) );
  OAI21_X4 U5050 ( .B1(n4096), .B2(n4095), .A(n1795), .ZN(n4105) );
  NOR3_X4 U5051 ( .A1(n4101), .A2(n4298), .A3(n4472), .ZN(net328168) );
  INV_X4 U5052 ( .A(net328160), .ZN(net328450) );
  OAI21_X4 U5053 ( .B1(n1364), .B2(net331363), .A(n4111), .ZN(n4117) );
  XNOR2_X2 U5054 ( .A(n4112), .B(n1332), .ZN(n4252) );
  NAND2_X2 U5055 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  INV_X4 U5056 ( .A(n4126), .ZN(n4129) );
  NOR2_X4 U5057 ( .A1(n4129), .A2(n4128), .ZN(n4131) );
  NOR3_X4 U5058 ( .A1(n4134), .A2(n4133), .A3(n4132), .ZN(n4205) );
  NAND2_X2 U5059 ( .A1(a[25]), .A2(net331329), .ZN(n4185) );
  INV_X4 U5060 ( .A(n4185), .ZN(n4182) );
  OAI21_X4 U5061 ( .B1(n4158), .B2(n4157), .A(n4156), .ZN(n4274) );
  INV_X4 U5062 ( .A(n4159), .ZN(n4278) );
  XNOR2_X2 U5063 ( .A(n1215), .B(n4278), .ZN(n4165) );
  INV_X4 U5064 ( .A(n4165), .ZN(n4163) );
  OAI21_X4 U5065 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n4164) );
  NAND2_X2 U5066 ( .A1(n4279), .A2(n4167), .ZN(n4169) );
  INV_X4 U5067 ( .A(n4169), .ZN(n4168) );
  NAND3_X4 U5068 ( .A1(n4168), .A2(a[27]), .A3(n2034), .ZN(n4275) );
  NAND2_X2 U5069 ( .A1(a[27]), .A2(n2035), .ZN(n4170) );
  NAND2_X2 U5070 ( .A1(n4170), .A2(n4169), .ZN(n4171) );
  XNOR2_X2 U5071 ( .A(n4274), .B(n4276), .ZN(n4173) );
  NAND2_X2 U5072 ( .A1(a[26]), .A2(net331343), .ZN(n4172) );
  NAND2_X2 U5073 ( .A1(n1165), .A2(n4172), .ZN(n4175) );
  INV_X4 U5074 ( .A(n4172), .ZN(n4174) );
  XNOR2_X2 U5075 ( .A(n4285), .B(n4181), .ZN(n4183) );
  NAND2_X2 U5076 ( .A1(n4182), .A2(n4183), .ZN(n4271) );
  INV_X4 U5077 ( .A(n4183), .ZN(n4184) );
  XNOR2_X2 U5078 ( .A(n4187), .B(n4186), .ZN(n4188) );
  NAND2_X2 U5079 ( .A1(a[23]), .A2(n2037), .ZN(n4304) );
  INV_X4 U5080 ( .A(n4304), .ZN(n4190) );
  XNOR2_X2 U5081 ( .A(net328331), .B(n4303), .ZN(n4191) );
  XNOR2_X2 U5082 ( .A(n4193), .B(n4192), .ZN(n4203) );
  NAND2_X2 U5083 ( .A1(product_in[29]), .A2(net331295), .ZN(net328118) );
  NAND2_X2 U5084 ( .A1(n4195), .A2(net331613), .ZN(n4206) );
  XNOR2_X2 U5085 ( .A(n4205), .B(n4204), .ZN(product_out[29]) );
  NOR2_X4 U5086 ( .A1(net328118), .A2(net328309), .ZN(n4254) );
  INV_X4 U5087 ( .A(n4209), .ZN(n4210) );
  INV_X4 U5088 ( .A(n4212), .ZN(n4214) );
  INV_X4 U5089 ( .A(n4215), .ZN(n4216) );
  NOR2_X4 U5090 ( .A1(n4222), .A2(n4221), .ZN(n4223) );
  NAND4_X2 U5091 ( .A1(n4224), .A2(n4225), .A3(n1421), .A4(n4223), .ZN(n4227)
         );
  INV_X4 U5092 ( .A(n4227), .ZN(n4236) );
  NOR2_X4 U5093 ( .A1(n2017), .A2(n4228), .ZN(n4235) );
  NAND2_X2 U5094 ( .A1(n4229), .A2(n4228), .ZN(n4231) );
  NOR3_X4 U5095 ( .A1(n4236), .A2(n4235), .A3(n4234), .ZN(n4250) );
  INV_X4 U5096 ( .A(n4238), .ZN(n4240) );
  NAND3_X2 U5098 ( .A1(net328264), .A2(n4247), .A3(n4246), .ZN(n4248) );
  OAI21_X4 U5099 ( .B1(n4250), .B2(n4249), .A(n4248), .ZN(net328113) );
  INV_X4 U5100 ( .A(net328113), .ZN(net328253) );
  NOR2_X4 U5101 ( .A1(n4253), .A2(n4254), .ZN(n4308) );
  INV_X4 U5102 ( .A(n4263), .ZN(n4266) );
  AOI21_X4 U5104 ( .B1(n4264), .B2(n4263), .A(n1860), .ZN(n4265) );
  OAI21_X4 U5105 ( .B1(net328222), .B2(n4266), .A(n4265), .ZN(n4292) );
  INV_X4 U5106 ( .A(net328051), .ZN(net328192) );
  NAND2_X2 U5107 ( .A1(a[26]), .A2(net331329), .ZN(n4342) );
  INV_X4 U5108 ( .A(n4342), .ZN(n4289) );
  OAI21_X4 U5109 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n4322) );
  NAND2_X2 U5110 ( .A1(n1215), .A2(n4278), .ZN(n4280) );
  INV_X4 U5111 ( .A(n4281), .ZN(n4282) );
  NAND2_X2 U5112 ( .A1(n1216), .A2(n4282), .ZN(n4339) );
  OAI21_X4 U5113 ( .B1(n1216), .B2(n4282), .A(n4339), .ZN(n4314) );
  XNOR2_X2 U5114 ( .A(n4316), .B(n4314), .ZN(n4309) );
  NAND2_X2 U5115 ( .A1(a[28]), .A2(n2035), .ZN(n4311) );
  XNOR2_X2 U5116 ( .A(n4322), .B(n4321), .ZN(n4333) );
  NAND2_X2 U5117 ( .A1(a[27]), .A2(net331341), .ZN(n4332) );
  NAND2_X2 U5118 ( .A1(n4287), .A2(n1368), .ZN(n4288) );
  NAND2_X2 U5119 ( .A1(a[24]), .A2(n2037), .ZN(net328083) );
  NAND2_X2 U5120 ( .A1(a[23]), .A2(net331305), .ZN(net328020) );
  INV_X4 U5121 ( .A(n4370), .ZN(n4301) );
  NOR3_X4 U5122 ( .A1(n4302), .A2(n4373), .A3(n4301), .ZN(net328128) );
  XNOR2_X2 U5123 ( .A(n4360), .B(n4303), .ZN(net328026) );
  AOI22_X2 U5124 ( .A1(n4305), .A2(n4359), .B1(n4304), .B2(n4391), .ZN(n4306)
         );
  OAI21_X4 U5125 ( .B1(n4307), .B2(n4306), .A(n1135), .ZN(net328025) );
  NAND2_X2 U5126 ( .A1(product_in[30]), .A2(net331295), .ZN(net328123) );
  XNOR2_X2 U5127 ( .A(n4313), .B(n4312), .ZN(n4320) );
  INV_X4 U5128 ( .A(n4314), .ZN(n4315) );
  XNOR2_X2 U5129 ( .A(n4318), .B(n4317), .ZN(n4319) );
  XNOR2_X2 U5130 ( .A(n4320), .B(n4319), .ZN(n4329) );
  NAND2_X2 U5131 ( .A1(net331341), .A2(a[28]), .ZN(n4323) );
  XNOR2_X2 U5132 ( .A(n4324), .B(n4323), .ZN(n4327) );
  NAND2_X2 U5133 ( .A1(a[29]), .A2(n2035), .ZN(n4326) );
  XNOR2_X2 U5134 ( .A(n4327), .B(n4326), .ZN(n4328) );
  XNOR2_X2 U5135 ( .A(n4329), .B(n4328), .ZN(n4351) );
  INV_X4 U5137 ( .A(n4334), .ZN(n4338) );
  NAND2_X2 U5138 ( .A1(a[26]), .A2(net331323), .ZN(n4336) );
  NAND2_X2 U5139 ( .A1(n2037), .A2(a[25]), .ZN(n4335) );
  XNOR2_X2 U5140 ( .A(n4336), .B(n4335), .ZN(n4337) );
  FA_X1 U5141 ( .A(n4338), .B(n1350), .CI(n4337), .S(n4348) );
  INV_X4 U5142 ( .A(n4339), .ZN(n4341) );
  NAND2_X2 U5143 ( .A1(a[24]), .A2(net331307), .ZN(n4340) );
  XNOR2_X2 U5144 ( .A(n4341), .B(n4340), .ZN(n4346) );
  OAI22_X2 U5145 ( .A1(n4344), .A2(n4352), .B1(n1770), .B2(n4342), .ZN(n4345)
         );
  XNOR2_X2 U5146 ( .A(n4345), .B(n4346), .ZN(n4347) );
  XNOR2_X2 U5147 ( .A(n4347), .B(n4348), .ZN(n4349) );
  FA_X1 U5148 ( .A(n4349), .B(n4351), .CI(n4350), .S(n4358) );
  INV_X4 U5149 ( .A(net328019), .ZN(net328039) );
  NAND2_X2 U5150 ( .A1(n4362), .A2(n1134), .ZN(n4364) );
  INV_X4 U5151 ( .A(net327997), .ZN(net328028) );
  NAND2_X2 U5152 ( .A1(product_in[31]), .A2(net331295), .ZN(net328003) );
  NOR2_X4 U5153 ( .A1(net328028), .A2(net327998), .ZN(net327999) );
  XNOR2_X2 U5154 ( .A(net328023), .B(n1112), .ZN(n4366) );
  NAND2_X2 U5155 ( .A1(net328021), .A2(n4366), .ZN(n4369) );
  INV_X4 U5156 ( .A(net328020), .ZN(net328016) );
  NAND2_X2 U5158 ( .A1(n4369), .A2(n4371), .ZN(n4375) );
  NAND2_X2 U1136 ( .A1(n3285), .A2(n3284), .ZN(n4455) );
  NAND2_X2 U1141 ( .A1(n2295), .A2(n2294), .ZN(n2441) );
  INV_X8 U1153 ( .A(net333677), .ZN(net333678) );
  INV_X4 U1158 ( .A(n1895), .ZN(n4386) );
  INV_X4 U1164 ( .A(n3227), .ZN(n1895) );
  INV_X2 U1165 ( .A(n3728), .ZN(n4387) );
  INV_X8 U1177 ( .A(n3728), .ZN(n3565) );
  NAND2_X4 U1181 ( .A1(n4406), .A2(n4420), .ZN(n3728) );
  OAI22_X4 U1182 ( .A1(net330942), .A2(n2377), .B1(n2371), .B2(n2376), .ZN(
        n2378) );
  INV_X8 U1190 ( .A(net330244), .ZN(n4388) );
  INV_X8 U1193 ( .A(net330244), .ZN(net334211) );
  CLKBUF_X3 U1196 ( .A(n4139), .Z(n4422) );
  NAND2_X4 U1218 ( .A1(n2195), .A2(n2343), .ZN(n2194) );
  OAI21_X4 U1221 ( .B1(n2195), .B2(n2343), .A(n2194), .ZN(n2197) );
  OAI221_X4 U1226 ( .B1(n2244), .B2(n2193), .C1(n2146), .C2(n2244), .A(n2243), 
        .ZN(n2195) );
  INV_X1 U1236 ( .A(n2706), .ZN(n2532) );
  INV_X4 U1242 ( .A(net331025), .ZN(net333770) );
  INV_X4 U1245 ( .A(n3763), .ZN(n1771) );
  INV_X2 U1253 ( .A(n3514), .ZN(n1776) );
  BUF_X8 U1271 ( .A(n2026), .Z(n1147) );
  INV_X4 U1282 ( .A(n3801), .ZN(n4389) );
  INV_X8 U1292 ( .A(n3976), .ZN(n3801) );
  AND2_X2 U1296 ( .A1(net330043), .A2(net330042), .ZN(n4390) );
  BUF_X4 U1303 ( .A(net329965), .Z(n4445) );
  INV_X8 U1309 ( .A(n2283), .ZN(n2372) );
  NAND2_X4 U1319 ( .A1(n1947), .A2(n4256), .ZN(n4391) );
  NAND2_X4 U1334 ( .A1(n4410), .A2(n4411), .ZN(n1947) );
  NAND2_X2 U1335 ( .A1(net332894), .A2(net332895), .ZN(n4392) );
  NAND2_X4 U1342 ( .A1(n3771), .A2(n3770), .ZN(n3773) );
  INV_X4 U1343 ( .A(net328585), .ZN(n1544) );
  NAND2_X4 U1344 ( .A1(net328912), .A2(n3768), .ZN(net328585) );
  NAND2_X2 U1358 ( .A1(n3564), .A2(n3563), .ZN(n4406) );
  INV_X8 U1360 ( .A(n1206), .ZN(n1207) );
  INV_X4 U1362 ( .A(net329990), .ZN(net329452) );
  NAND2_X4 U1370 ( .A1(n3094), .A2(n3093), .ZN(n1794) );
  XNOR2_X2 U1371 ( .A(n3979), .B(n3891), .ZN(n4393) );
  NAND2_X2 U1373 ( .A1(n1991), .A2(n2169), .ZN(n2173) );
  INV_X8 U1385 ( .A(net331476), .ZN(net331477) );
  AND2_X2 U1387 ( .A1(n2434), .A2(n2435), .ZN(n4394) );
  INV_X8 U1397 ( .A(net328229), .ZN(n1397) );
  NAND2_X4 U1410 ( .A1(net329451), .A2(n3431), .ZN(n3342) );
  INV_X2 U1415 ( .A(net328607), .ZN(net328606) );
  NAND2_X2 U1416 ( .A1(net328385), .A2(net328485), .ZN(n4395) );
  NAND2_X4 U1420 ( .A1(n3112), .A2(n1211), .ZN(n4396) );
  INV_X8 U1421 ( .A(n3562), .ZN(n1992) );
  NOR2_X4 U1423 ( .A1(net328389), .A2(n4269), .ZN(n4073) );
  INV_X8 U1442 ( .A(n4012), .ZN(n1956) );
  NAND2_X1 U1449 ( .A1(net328864), .A2(net328865), .ZN(n4399) );
  NAND2_X2 U1455 ( .A1(n4397), .A2(n4398), .ZN(n4400) );
  NAND2_X2 U1476 ( .A1(n4399), .A2(n4400), .ZN(n1518) );
  INV_X1 U1479 ( .A(net328864), .ZN(n4397) );
  INV_X2 U1485 ( .A(net328865), .ZN(n4398) );
  NAND2_X2 U1510 ( .A1(net328616), .A2(n3894), .ZN(n4401) );
  NAND2_X4 U1514 ( .A1(n4402), .A2(net328752), .ZN(n3896) );
  INV_X4 U1520 ( .A(n4401), .ZN(n4402) );
  INV_X2 U1524 ( .A(n3515), .ZN(n1688) );
  INV_X8 U1571 ( .A(n4392), .ZN(net328583) );
  AND2_X4 U1574 ( .A1(net332558), .A2(net328167), .ZN(net328148) );
  INV_X4 U1593 ( .A(n1979), .ZN(n3656) );
  INV_X2 U1607 ( .A(n1700), .ZN(n4144) );
  INV_X8 U1616 ( .A(n3415), .ZN(n1925) );
  NAND2_X4 U1690 ( .A1(n4163), .A2(n4164), .ZN(n4279) );
  BUF_X4 U1694 ( .A(n4343), .Z(n1770) );
  XNOR2_X2 U1697 ( .A(n4343), .B(n4342), .ZN(n4352) );
  INV_X8 U1698 ( .A(net328573), .ZN(n1546) );
  INV_X8 U1706 ( .A(n1970), .ZN(n4444) );
  INV_X4 U1724 ( .A(n3412), .ZN(n3508) );
  INV_X2 U1728 ( .A(net328593), .ZN(n4403) );
  INV_X8 U1740 ( .A(net328794), .ZN(net328593) );
  NAND2_X4 U1744 ( .A1(n4404), .A2(n4405), .ZN(n4407) );
  NAND2_X4 U1746 ( .A1(n4406), .A2(n4407), .ZN(n1405) );
  INV_X2 U1747 ( .A(n3564), .ZN(n4404) );
  INV_X1 U1748 ( .A(n3563), .ZN(n4405) );
  NAND2_X1 U1779 ( .A1(n4079), .A2(n4078), .ZN(n4410) );
  NAND2_X2 U1815 ( .A1(n4408), .A2(n4409), .ZN(n4411) );
  INV_X2 U1817 ( .A(n4079), .ZN(n4408) );
  INV_X4 U1825 ( .A(n4078), .ZN(n4409) );
  INV_X8 U1831 ( .A(net329598), .ZN(n4477) );
  NAND2_X1 U1858 ( .A1(n3198), .A2(n3195), .ZN(n4414) );
  NAND2_X4 U1861 ( .A1(n4412), .A2(n4413), .ZN(n4415) );
  NAND2_X4 U1869 ( .A1(n4414), .A2(n4415), .ZN(n3073) );
  INV_X4 U1870 ( .A(n3198), .ZN(n4412) );
  INV_X2 U1902 ( .A(n3195), .ZN(n4413) );
  INV_X4 U1920 ( .A(n3477), .ZN(n1488) );
  CLKBUF_X3 U1924 ( .A(n3899), .Z(n1507) );
  NOR2_X4 U1938 ( .A1(n4258), .A2(n4257), .ZN(n4261) );
  INV_X2 U1946 ( .A(n1655), .ZN(n3246) );
  INV_X8 U1948 ( .A(n4148), .ZN(n4270) );
  NAND2_X2 U1950 ( .A1(n1933), .A2(n1934), .ZN(n4416) );
  XNOR2_X2 U1955 ( .A(n3088), .B(n3087), .ZN(n4417) );
  NAND2_X2 U1986 ( .A1(n4418), .A2(n4419), .ZN(n4420) );
  INV_X4 U2065 ( .A(n3564), .ZN(n4418) );
  INV_X1 U2066 ( .A(n3563), .ZN(n4419) );
  OAI221_X4 U2067 ( .B1(n3514), .B2(n3420), .C1(n3421), .C2(n1836), .A(n3383), 
        .ZN(n4443) );
  INV_X8 U2081 ( .A(n3758), .ZN(n1734) );
  INV_X2 U2095 ( .A(n1955), .ZN(n4421) );
  INV_X8 U2099 ( .A(n1963), .ZN(n3678) );
  OAI21_X2 U2110 ( .B1(n3030), .B2(n2848), .A(n2792), .ZN(n1128) );
  NAND2_X2 U2114 ( .A1(n3030), .A2(n2848), .ZN(net329986) );
  INV_X2 U2122 ( .A(n3030), .ZN(n1201) );
  BUF_X16 U2138 ( .A(net328593), .Z(net332214) );
  INV_X8 U2141 ( .A(net329985), .ZN(net334441) );
  INV_X4 U2167 ( .A(n3315), .ZN(n4423) );
  INV_X4 U2177 ( .A(n3315), .ZN(n2998) );
  INV_X2 U2217 ( .A(n1187), .ZN(n2503) );
  INV_X2 U2228 ( .A(n2911), .ZN(n4424) );
  INV_X32 U2232 ( .A(control[1]), .ZN(n4425) );
  INV_X32 U2234 ( .A(control[1]), .ZN(n4426) );
  INV_X16 U2241 ( .A(control[1]), .ZN(n4427) );
  INV_X32 U2242 ( .A(control[1]), .ZN(n4428) );
  NOR2_X4 U2245 ( .A1(n2064), .A2(n2065), .ZN(n4429) );
  INV_X4 U2255 ( .A(n4429), .ZN(n2091) );
  INV_X2 U2258 ( .A(n2065), .ZN(n2066) );
  BUF_X32 U2272 ( .A(n3923), .Z(n4430) );
  INV_X4 U2282 ( .A(n2407), .ZN(n3923) );
  NAND2_X4 U2285 ( .A1(n2974), .A2(n2973), .ZN(n3670) );
  NAND3_X2 U2292 ( .A1(n1124), .A2(n1689), .A3(n2973), .ZN(n4431) );
  INV_X2 U2308 ( .A(n2825), .ZN(n1689) );
  NAND2_X4 U2318 ( .A1(n1622), .A2(n1115), .ZN(n2994) );
  INV_X8 U2336 ( .A(n3393), .ZN(n1364) );
  XNOR2_X2 U2366 ( .A(n3577), .B(n3743), .ZN(product_out[23]) );
  INV_X4 U2374 ( .A(n3577), .ZN(n3751) );
  NAND2_X2 U2385 ( .A1(n2694), .A2(n2695), .ZN(n4432) );
  NAND2_X4 U2410 ( .A1(n2694), .A2(n2695), .ZN(n4433) );
  NAND2_X2 U2433 ( .A1(n2694), .A2(n2695), .ZN(n2838) );
  NAND2_X4 U2436 ( .A1(n1316), .A2(n1317), .ZN(n2694) );
  NAND2_X2 U2449 ( .A1(n1787), .A2(n3829), .ZN(n3831) );
  NAND2_X2 U2465 ( .A1(n3481), .A2(n3480), .ZN(n4434) );
  NAND2_X2 U2473 ( .A1(n3481), .A2(n3480), .ZN(n1619) );
  INV_X4 U2479 ( .A(n3390), .ZN(n3388) );
  INV_X4 U2491 ( .A(n3600), .ZN(n3763) );
  OAI21_X2 U2523 ( .B1(n4014), .B2(n3947), .A(n1280), .ZN(n1962) );
  INV_X4 U2525 ( .A(n3850), .ZN(n3829) );
  NAND2_X4 U2563 ( .A1(net332668), .A2(n3031), .ZN(n3032) );
  CLKBUF_X2 U2573 ( .A(n3726), .Z(n4435) );
  INV_X4 U2574 ( .A(n1786), .ZN(n1787) );
  XNOR2_X1 U2576 ( .A(n2186), .B(n2185), .ZN(n4436) );
  OAI21_X4 U2578 ( .B1(n1738), .B2(net331295), .A(n4221), .ZN(n3840) );
  INV_X8 U2582 ( .A(n3840), .ZN(n3574) );
  INV_X4 U2589 ( .A(n2187), .ZN(n4437) );
  INV_X4 U2616 ( .A(n4437), .ZN(n4438) );
  XNOR2_X1 U2640 ( .A(n2118), .B(n4453), .ZN(n4439) );
  NAND2_X2 U2664 ( .A1(n2089), .A2(n2088), .ZN(n4453) );
  XNOR2_X2 U2683 ( .A(n2269), .B(n4440), .ZN(n1624) );
  INV_X32 U2696 ( .A(n1339), .ZN(n4440) );
  XNOR2_X2 U2744 ( .A(n2955), .B(n3026), .ZN(n1299) );
  INV_X2 U2745 ( .A(n3332), .ZN(n4441) );
  INV_X4 U2779 ( .A(n4441), .ZN(n4442) );
  INV_X8 U2781 ( .A(n4211), .ZN(n3395) );
  NAND2_X2 U2818 ( .A1(n4087), .A2(n4085), .ZN(n3845) );
  INV_X2 U2834 ( .A(n2966), .ZN(n1677) );
  AND2_X4 U2836 ( .A1(n3963), .A2(n3580), .ZN(n1970) );
  INV_X4 U2838 ( .A(net328562), .ZN(net332946) );
  INV_X8 U2851 ( .A(n3759), .ZN(n4449) );
  INV_X4 U2856 ( .A(n2177), .ZN(n2471) );
  NAND3_X2 U2871 ( .A1(n3349), .A2(n3348), .A3(net329441), .ZN(n1788) );
  XNOR2_X1 U2890 ( .A(net333311), .B(n4446), .ZN(n1574) );
  XOR2_X2 U2893 ( .A(net328047), .B(net328020), .Z(n4446) );
  INV_X2 U2894 ( .A(net333311), .ZN(net328046) );
  NAND2_X2 U2912 ( .A1(n1898), .A2(n1899), .ZN(n4447) );
  INV_X4 U2914 ( .A(n1171), .ZN(n1899) );
  INV_X8 U2925 ( .A(n2482), .ZN(n1921) );
  INV_X2 U2929 ( .A(n4076), .ZN(n4264) );
  XOR2_X2 U2941 ( .A(n1647), .B(n3943), .Z(n4469) );
  NAND4_X2 U2946 ( .A1(n2073), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2074)
         );
  NAND2_X4 U2948 ( .A1(n2082), .A2(n2178), .ZN(n1808) );
  NAND2_X4 U2980 ( .A1(n3063), .A2(n3064), .ZN(n4448) );
  INV_X8 U2985 ( .A(n1344), .ZN(n1406) );
  NOR2_X4 U2994 ( .A1(n4298), .A2(n4100), .ZN(n4091) );
  INV_X2 U3019 ( .A(n3759), .ZN(n4085) );
  NAND2_X2 U3021 ( .A1(net332856), .A2(net332855), .ZN(n4450) );
  NAND2_X4 U3022 ( .A1(n1875), .A2(n1876), .ZN(net332856) );
  NAND2_X2 U3030 ( .A1(n2230), .A2(n1618), .ZN(net330854) );
  INV_X2 U3040 ( .A(n2757), .ZN(n2021) );
  INV_X4 U3042 ( .A(n2382), .ZN(n1745) );
  INV_X2 U3044 ( .A(net333621), .ZN(net330596) );
  NAND2_X1 U3050 ( .A1(net330918), .A2(n2365), .ZN(n4451) );
  NAND2_X4 U3078 ( .A1(n2360), .A2(n2557), .ZN(n2658) );
  NAND2_X4 U3085 ( .A1(net328472), .A2(n1506), .ZN(net328176) );
  NAND2_X2 U3112 ( .A1(net328473), .A2(net328474), .ZN(n1506) );
  INV_X4 U3113 ( .A(net333078), .ZN(net332292) );
  INV_X2 U3115 ( .A(net330029), .ZN(net333078) );
  INV_X2 U3118 ( .A(net328584), .ZN(net328917) );
  NAND2_X4 U3132 ( .A1(net331084), .A2(net331083), .ZN(n2130) );
  NAND2_X2 U3139 ( .A1(n1127), .A2(n2139), .ZN(n2189) );
  INV_X4 U3146 ( .A(n2591), .ZN(n1964) );
  NAND2_X4 U3147 ( .A1(n4077), .A2(n4076), .ZN(n4452) );
  NAND2_X2 U3166 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  AOI21_X2 U3169 ( .B1(n1641), .B2(n1291), .A(n3238), .ZN(n3244) );
  NAND2_X4 U3188 ( .A1(net328016), .A2(n4368), .ZN(n4371) );
  OAI21_X4 U3191 ( .B1(n3629), .B2(n3628), .A(n1144), .ZN(n1658) );
  INV_X2 U3196 ( .A(n2276), .ZN(n1171) );
  NAND2_X4 U3221 ( .A1(n3599), .A2(n1331), .ZN(n3758) );
  NOR2_X4 U3228 ( .A1(n2931), .A2(n2930), .ZN(n2934) );
  INV_X16 U3256 ( .A(n2443), .ZN(n2566) );
  INV_X2 U3276 ( .A(n3270), .ZN(n3271) );
  OAI221_X4 U3286 ( .B1(net329339), .B2(net329340), .C1(net333569), .C2(
        net329459), .A(n4482), .ZN(n1523) );
  INV_X4 U3312 ( .A(n3029), .ZN(n3034) );
  INV_X8 U3335 ( .A(n4354), .ZN(n4344) );
  OAI21_X4 U3347 ( .B1(n4272), .B2(n4273), .A(n1775), .ZN(n4354) );
  NAND2_X4 U3363 ( .A1(n2345), .A2(n2426), .ZN(n2347) );
  NAND2_X2 U3374 ( .A1(n2389), .A2(n1223), .ZN(n1224) );
  OAI211_X4 U3381 ( .C1(n2984), .C2(n2983), .A(n2981), .B(n1687), .ZN(n1680)
         );
  NAND2_X1 U3399 ( .A1(n2152), .A2(n2151), .ZN(n2155) );
  NAND2_X4 U3403 ( .A1(n2155), .A2(n2254), .ZN(net328250) );
  INV_X2 U3420 ( .A(n2254), .ZN(n2256) );
  NAND2_X4 U3423 ( .A1(n2154), .A2(n2153), .ZN(n2254) );
  INV_X8 U3459 ( .A(n2619), .ZN(n2624) );
  XNOR2_X1 U3462 ( .A(n3308), .B(n1220), .ZN(product_out[19]) );
  AOI21_X2 U3465 ( .B1(n3313), .B2(n3314), .A(n3312), .ZN(n3396) );
  AOI21_X4 U3472 ( .B1(n1557), .B2(n1315), .A(net329971), .ZN(net329968) );
  INV_X4 U3476 ( .A(n3065), .ZN(n1398) );
  INV_X8 U3497 ( .A(n1865), .ZN(n4460) );
  NAND2_X2 U3503 ( .A1(n2380), .A2(n2381), .ZN(n2557) );
  INV_X16 U3505 ( .A(net332666), .ZN(net332668) );
  INV_X4 U3522 ( .A(n3739), .ZN(n3735) );
  INV_X2 U3532 ( .A(n1644), .ZN(n1627) );
  NAND2_X2 U3571 ( .A1(n1644), .A2(n3927), .ZN(n3747) );
  AND2_X2 U3584 ( .A1(n3579), .A2(n1619), .ZN(n1401) );
  INV_X2 U3588 ( .A(net328450), .ZN(n4454) );
  INV_X4 U3596 ( .A(n3738), .ZN(n3753) );
  NAND2_X2 U3633 ( .A1(n3738), .A2(net331299), .ZN(n4479) );
  INV_X8 U3667 ( .A(n1906), .ZN(n1907) );
  OR2_X2 U3683 ( .A1(n4012), .A2(n4013), .ZN(n3854) );
  OAI21_X4 U3691 ( .B1(n1683), .B2(n3727), .A(n4434), .ZN(n3959) );
  INV_X8 U3701 ( .A(n3959), .ZN(n3732) );
  NAND2_X4 U3751 ( .A1(n3579), .A2(n3578), .ZN(n3729) );
  NAND2_X4 U3762 ( .A1(n3579), .A2(n3578), .ZN(n1418) );
  INV_X4 U3765 ( .A(n2117), .ZN(n2114) );
  INV_X8 U3789 ( .A(n2174), .ZN(n2221) );
  OAI21_X4 U3814 ( .B1(n3224), .B2(n3326), .A(n3327), .ZN(n4467) );
  OAI211_X2 U3841 ( .C1(n3329), .C2(n3330), .A(n3328), .B(n1113), .ZN(n3387)
         );
  AOI211_X4 U3865 ( .C1(n1192), .C2(n1774), .A(n4215), .B(n3570), .ZN(n1125)
         );
  INV_X1 U3880 ( .A(n1360), .ZN(n1361) );
  NOR2_X2 U3881 ( .A1(n3826), .A2(n3814), .ZN(n3822) );
  NAND2_X4 U3909 ( .A1(n2027), .A2(n3227), .ZN(n2028) );
  NOR3_X2 U3912 ( .A1(n2282), .A2(n1736), .A3(n1110), .ZN(n2285) );
  INV_X8 U3923 ( .A(n1150), .ZN(n3338) );
  INV_X8 U3945 ( .A(n3338), .ZN(n1777) );
  NAND2_X4 U3946 ( .A1(n3311), .A2(n3310), .ZN(n3397) );
  NAND2_X4 U3947 ( .A1(n2380), .A2(n2381), .ZN(n4456) );
  NAND2_X4 U3974 ( .A1(net331499), .A2(net330994), .ZN(net331068) );
  INV_X8 U3999 ( .A(n2218), .ZN(n2219) );
  NAND2_X2 U4049 ( .A1(n3732), .A2(n3958), .ZN(n4457) );
  NAND2_X2 U4066 ( .A1(n3732), .A2(n3958), .ZN(n3848) );
  INV_X8 U4077 ( .A(n3295), .ZN(n3296) );
  NAND2_X4 U4091 ( .A1(n2593), .A2(n2594), .ZN(n4458) );
  NAND2_X2 U4111 ( .A1(n2593), .A2(n2594), .ZN(n2837) );
  NAND2_X2 U4115 ( .A1(n2229), .A2(n2175), .ZN(n1829) );
  NAND2_X2 U4163 ( .A1(n3953), .A2(n1795), .ZN(n3971) );
  CLKBUF_X3 U4166 ( .A(net331097), .Z(net333618) );
  NAND2_X4 U4181 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  NAND3_X2 U4183 ( .A1(net328415), .A2(net333918), .A3(n1584), .ZN(net328414)
         );
  BUF_X4 U4193 ( .A(n1111), .Z(net333918) );
  INV_X1 U4196 ( .A(n3080), .ZN(n3078) );
  NAND2_X4 U4203 ( .A1(n2363), .A2(n1143), .ZN(n2299) );
  NAND2_X4 U4221 ( .A1(n3940), .A2(n1404), .ZN(n3941) );
  INV_X4 U4241 ( .A(n3207), .ZN(n2966) );
  INV_X4 U4297 ( .A(n3171), .ZN(n1913) );
  NAND2_X4 U4300 ( .A1(net332987), .A2(net332988), .ZN(n1848) );
  XNOR2_X2 U4301 ( .A(net333311), .B(n4459), .ZN(net328024) );
  INV_X32 U4312 ( .A(n1690), .ZN(n4459) );
  NAND2_X4 U4348 ( .A1(n4491), .A2(n4492), .ZN(n1865) );
  BUF_X8 U4403 ( .A(net328024), .Z(n1112) );
  INV_X4 U4441 ( .A(net327992), .ZN(n1478) );
  OAI21_X2 U4447 ( .B1(n2172), .B2(n1881), .A(n2228), .ZN(n2176) );
  NAND2_X4 U4481 ( .A1(n1611), .A2(net331073), .ZN(net334039) );
  NAND2_X1 U4505 ( .A1(n1611), .A2(net331073), .ZN(n1608) );
  INV_X8 U4512 ( .A(n3672), .ZN(n3204) );
  NAND2_X2 U4518 ( .A1(n4262), .A2(n4263), .ZN(n4461) );
  INV_X2 U4527 ( .A(n1860), .ZN(n4262) );
  NAND2_X4 U4596 ( .A1(net329558), .A2(net329557), .ZN(n4462) );
  INV_X1 U4607 ( .A(n2088), .ZN(n4463) );
  NAND2_X2 U4613 ( .A1(net328851), .A2(n3808), .ZN(n1425) );
  NOR2_X4 U4616 ( .A1(net328171), .A2(net328475), .ZN(net328170) );
  INV_X4 U4635 ( .A(net328475), .ZN(net328409) );
  NAND4_X4 U4638 ( .A1(n2556), .A2(n2555), .A3(n1460), .A4(n1667), .ZN(n2558)
         );
  OAI21_X2 U4702 ( .B1(n1606), .B2(net330039), .A(n1607), .ZN(net334227) );
  OAI211_X4 U4720 ( .C1(n2709), .C2(n2708), .A(n3019), .B(n2707), .ZN(n2710)
         );
  NAND2_X2 U4749 ( .A1(n1682), .A2(n2531), .ZN(n2708) );
  NAND2_X4 U4812 ( .A1(n4228), .A2(n1404), .ZN(n3743) );
  NAND2_X1 U4894 ( .A1(n4228), .A2(n3927), .ZN(n3748) );
  AOI211_X4 U4897 ( .C1(n4233), .C2(n4232), .A(n4231), .B(n4230), .ZN(n4234)
         );
  INV_X8 U4904 ( .A(net330843), .ZN(n1313) );
  INV_X4 U4925 ( .A(n2656), .ZN(n4464) );
  INV_X8 U4929 ( .A(n2281), .ZN(n1902) );
  CLKBUF_X3 U5008 ( .A(net330834), .Z(net333816) );
  INV_X1 U5097 ( .A(n2134), .ZN(n2135) );
  INV_X8 U5103 ( .A(n1648), .ZN(n3030) );
  OAI21_X4 U5136 ( .B1(n2511), .B2(n2510), .A(n2509), .ZN(n4465) );
  OAI21_X2 U5157 ( .B1(n2511), .B2(n2510), .A(n2509), .ZN(n2722) );
  INV_X8 U5159 ( .A(n2476), .ZN(n2560) );
  INV_X4 U5160 ( .A(n2099), .ZN(n2052) );
  INV_X8 U5161 ( .A(n4360), .ZN(n4307) );
  BUF_X32 U5162 ( .A(n3815), .Z(n1133) );
  INV_X1 U5163 ( .A(n1277), .ZN(n4466) );
  OAI21_X4 U5164 ( .B1(n1297), .B2(n3222), .A(n3408), .ZN(n3326) );
  INV_X2 U5165 ( .A(net333275), .ZN(net330612) );
  INV_X8 U5166 ( .A(net329965), .ZN(net329753) );
  NAND2_X4 U5167 ( .A1(n1540), .A2(net330330), .ZN(n4468) );
  INV_X4 U5168 ( .A(n1168), .ZN(n4112) );
  INV_X2 U5169 ( .A(n3483), .ZN(n2725) );
  XNOR2_X2 U5170 ( .A(n3484), .B(n3483), .ZN(n4194) );
  OAI21_X4 U5171 ( .B1(n1357), .B2(n1917), .A(n1238), .ZN(n3483) );
  INV_X2 U5172 ( .A(n1376), .ZN(net330942) );
  NAND2_X1 U5173 ( .A1(net331479), .A2(net328408), .ZN(n4470) );
  INV_X4 U5174 ( .A(n2182), .ZN(n1875) );
  INV_X2 U5175 ( .A(net333424), .ZN(net328247) );
  AOI21_X1 U5176 ( .B1(n3192), .B2(n3191), .A(n3495), .ZN(n3308) );
  INV_X8 U5177 ( .A(net329453), .ZN(net329824) );
  INV_X4 U5178 ( .A(n4100), .ZN(n4471) );
  INV_X4 U5179 ( .A(n4471), .ZN(n4472) );
  INV_X4 U5180 ( .A(n3250), .ZN(n3253) );
  NAND2_X4 U5181 ( .A1(n3249), .A2(n3248), .ZN(n1743) );
  NOR2_X2 U5182 ( .A1(net328254), .A2(n4241), .ZN(n4242) );
  NAND2_X4 U5183 ( .A1(n2794), .A2(n2795), .ZN(n3065) );
  INV_X1 U5184 ( .A(n2796), .ZN(n2795) );
  NAND2_X2 U5185 ( .A1(n1384), .A2(n4473), .ZN(n4474) );
  INV_X2 U5186 ( .A(net328794), .ZN(n4473) );
  INV_X4 U5187 ( .A(n4474), .ZN(net328791) );
  AOI21_X4 U5188 ( .B1(n2367), .B2(n2369), .A(n2368), .ZN(n2383) );
  NAND3_X4 U5189 ( .A1(n4294), .A2(n4355), .A3(n4475), .ZN(n4476) );
  INV_X4 U5190 ( .A(net328083), .ZN(n4475) );
  INV_X8 U5191 ( .A(n4476), .ZN(n4350) );
  NAND2_X2 U5192 ( .A1(n4176), .A2(n4043), .ZN(n4001) );
  NAND3_X4 U5193 ( .A1(n3110), .A2(n4396), .A3(n4477), .ZN(n4478) );
  INV_X8 U5194 ( .A(n4478), .ZN(n3113) );
  OAI211_X4 U5195 ( .C1(n2782), .C2(n1415), .A(n2780), .B(n2781), .ZN(n2919)
         );
  INV_X8 U5196 ( .A(n4456), .ZN(n2782) );
  AOI21_X4 U5197 ( .B1(n2435), .B2(n2434), .A(n1829), .ZN(n2783) );
  AOI21_X2 U5198 ( .B1(n1991), .B2(n2169), .A(n2221), .ZN(n2172) );
  OAI21_X2 U5199 ( .B1(n4454), .B2(n4299), .A(net328162), .ZN(n4300) );
  NOR2_X4 U5200 ( .A1(n2787), .A2(n2788), .ZN(n2789) );
  INV_X4 U5201 ( .A(n4479), .ZN(n3734) );
  INV_X16 U5202 ( .A(net328006), .ZN(net331299) );
  CLKBUF_X3 U5203 ( .A(n2166), .Z(n1650) );
  NAND3_X2 U5204 ( .A1(n2566), .A2(n2565), .A3(n1862), .ZN(n4480) );
  BUF_X16 U5205 ( .A(n4355), .Z(n4481) );
  NAND2_X2 U5206 ( .A1(n1330), .A2(net329556), .ZN(n4482) );
  NAND2_X2 U5207 ( .A1(n1330), .A2(net329556), .ZN(net329343) );
  INV_X8 U5208 ( .A(net331353), .ZN(net331351) );
  XNOR2_X2 U5209 ( .A(net331072), .B(net331061), .ZN(net331030) );
  INV_X8 U5210 ( .A(n1410), .ZN(n1411) );
  INV_X1 U5211 ( .A(net331357), .ZN(n4483) );
  INV_X4 U5212 ( .A(n3102), .ZN(n2883) );
  INV_X2 U5213 ( .A(n4257), .ZN(n4484) );
  INV_X2 U5214 ( .A(n4359), .ZN(n4257) );
  NAND3_X4 U5215 ( .A1(a[13]), .A2(n2765), .A3(net331349), .ZN(n3131) );
  NOR2_X2 U5216 ( .A1(n3121), .A2(n3122), .ZN(n3123) );
  BUF_X4 U5217 ( .A(n3131), .Z(n1487) );
  INV_X8 U5218 ( .A(n2177), .ZN(n1420) );
  INV_X4 U5219 ( .A(net329472), .ZN(n4485) );
  INV_X8 U5220 ( .A(n2643), .ZN(n4486) );
  INV_X4 U5221 ( .A(n2643), .ZN(n2702) );
  INV_X8 U5222 ( .A(n3098), .ZN(n3099) );
  INV_X4 U5223 ( .A(n1422), .ZN(n4487) );
  XNOR2_X2 U5224 ( .A(n1645), .B(n4452), .ZN(n1422) );
  INV_X4 U5225 ( .A(net328873), .ZN(net329014) );
  NAND2_X1 U5226 ( .A1(n2563), .A2(n2562), .ZN(n2565) );
  NAND2_X4 U5227 ( .A1(n2420), .A2(n2392), .ZN(n2393) );
  NAND2_X2 U5228 ( .A1(n2412), .A2(n2411), .ZN(n2392) );
  NAND2_X1 U5229 ( .A1(n2557), .A2(n2781), .ZN(n2382) );
  INV_X4 U5230 ( .A(net331353), .ZN(n4488) );
  XNOR2_X2 U5231 ( .A(n2060), .B(n2059), .ZN(n1679) );
  INV_X8 U5232 ( .A(n1387), .ZN(n1388) );
  INV_X2 U5233 ( .A(n2125), .ZN(n2371) );
  NAND2_X1 U5234 ( .A1(n2490), .A2(n2547), .ZN(n4491) );
  NAND2_X2 U5235 ( .A1(n4489), .A2(n4490), .ZN(n4492) );
  INV_X2 U5236 ( .A(n2490), .ZN(n4489) );
  INV_X1 U5237 ( .A(n2547), .ZN(n4490) );
  NAND2_X4 U5238 ( .A1(n4460), .A2(n2492), .ZN(n4493) );
endmodule

