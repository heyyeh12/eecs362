module testbench;
	reg [31:0] A;
	wire Z;

	nor32to1 nor32to1(.a(A),.z(Z));

	initial begin
		$monitor("A = %h Z = %b", A, Z);
		#0 A = 32'h00000000;
		#1 A = 32'h00000001;
		#1 A = 32'h00000002; 
		#1 A = 32'h00000004;
		#1 A = 32'h00000008;
		#1 A = 32'h00000010;
		#1 A = 32'h00000020; 
		#1 A = 32'h00000040;
		#1 A = 32'h00000080;
		#1 A = 32'h00000100;
		#1 A = 32'h00000200; 
		#1 A = 32'h00000400;
		#1 A = 32'h00000800;
		#1 A = 32'h00001000;
		#1 A = 32'h00002000; 
		#1 A = 32'h00004000;
		#1 A = 32'h00008000;
		#1 A = 32'h00010000;
		#1 A = 32'h00020000; 
		#1 A = 32'h00040000;
		#1 A = 32'h00080000;
		#1 A = 32'h00100000;
		#1 A = 32'h00200000; 
		#1 A = 32'h00400000;
		#1 A = 32'h00800000;
		
	end
endmodule

