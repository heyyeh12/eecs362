
module ex ( aluSrc, aluCtrl, setInv, zeroExt, busA, busB, imm32, aluRes, 
        isZero, fp );
  input [3:0] aluCtrl;
  input [31:0] busA;
  input [31:0] busB;
  input [31:0] imm32;
  output [31:0] aluRes;
  input aluSrc, setInv, zeroExt, fp;
  output isZero;
  wire   n184, n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n267, n299, n439, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178;

  NAND4_X2 U3 ( .A1(n196), .A2(n197), .A3(n198), .A4(n199), .ZN(n195) );
  NOR4_X2 U4 ( .A1(busA[23]), .A2(busA[22]), .A3(busA[21]), .A4(busA[20]), 
        .ZN(n199) );
  NOR4_X2 U5 ( .A1(busA[1]), .A2(busA[19]), .A3(busA[18]), .A4(busA[17]), .ZN(
        n198) );
  NOR4_X2 U6 ( .A1(busA[16]), .A2(busA[15]), .A3(busA[14]), .A4(busA[13]), 
        .ZN(n197) );
  NOR4_X2 U7 ( .A1(busA[12]), .A2(busA[11]), .A3(busA[10]), .A4(busA[0]), .ZN(
        n196) );
  NAND4_X2 U8 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(n194) );
  NOR4_X2 U9 ( .A1(busA[9]), .A2(busA[8]), .A3(busA[7]), .A4(busA[6]), .ZN(
        n203) );
  NOR4_X2 U10 ( .A1(busA[5]), .A2(busA[4]), .A3(busA[3]), .A4(busA[31]), .ZN(
        n202) );
  NOR4_X2 U11 ( .A1(busA[30]), .A2(busA[2]), .A3(busA[29]), .A4(busA[28]), 
        .ZN(n201) );
  NOR4_X2 U12 ( .A1(busA[27]), .A2(busA[26]), .A3(busA[25]), .A4(busA[24]), 
        .ZN(n200) );
  OAI22_X2 U55 ( .A1(n190), .A2(n853), .B1(fp), .B2(n267), .ZN(aluRes[3]) );
  OAI22_X2 U75 ( .A1(n191), .A2(n853), .B1(fp), .B2(n299), .ZN(aluRes[2]) );
  OAI22_X2 U179 ( .A1(n192), .A2(n853), .B1(fp), .B2(n439), .ZN(aluRes[1]) );
  INV_X4 U800 ( .A(busA[9]), .ZN(n184) );
  INV_X4 U806 ( .A(busA[3]), .ZN(n190) );
  INV_X4 U807 ( .A(busA[2]), .ZN(n191) );
  INV_X4 U808 ( .A(busA[1]), .ZN(n192) );
  NAND2_X4 U811 ( .A1(n1771), .A2(n1526), .ZN(n969) );
  NAND4_X4 U812 ( .A1(n1396), .A2(n1397), .A3(n1395), .A4(n1394), .ZN(n1453)
         );
  NOR2_X2 U813 ( .A1(n1930), .A2(n1824), .ZN(n1395) );
  INV_X8 U814 ( .A(n830), .ZN(n831) );
  OAI221_X2 U815 ( .B1(n831), .B2(n1521), .C1(n829), .C2(n2082), .A(n837), 
        .ZN(n1771) );
  INV_X1 U816 ( .A(n827), .ZN(n1415) );
  NAND2_X4 U817 ( .A1(n1829), .A2(n1093), .ZN(n1264) );
  INV_X8 U818 ( .A(n1091), .ZN(n1111) );
  XNOR2_X2 U819 ( .A(n1028), .B(n1027), .ZN(n1056) );
  XNOR2_X2 U820 ( .A(n1329), .B(n1328), .ZN(n1824) );
  INV_X4 U821 ( .A(n839), .ZN(n838) );
  INV_X8 U822 ( .A(n839), .ZN(n837) );
  INV_X8 U823 ( .A(n822), .ZN(n1591) );
  NOR2_X2 U824 ( .A1(n1792), .A2(n1791), .ZN(n1793) );
  NOR2_X2 U825 ( .A1(n1833), .A2(n798), .ZN(n1792) );
  NOR2_X2 U826 ( .A1(n1832), .A2(n784), .ZN(n1791) );
  NOR2_X2 U827 ( .A1(n1759), .A2(n1758), .ZN(n1760) );
  NOR2_X2 U828 ( .A1(n1756), .A2(n798), .ZN(n1759) );
  NOR2_X2 U829 ( .A1(n1757), .A2(n784), .ZN(n1758) );
  NOR3_X2 U830 ( .A1(n925), .A2(n924), .A3(n2067), .ZN(n926) );
  NOR3_X2 U831 ( .A1(n1984), .A2(n790), .A3(n1393), .ZN(n1394) );
  NAND3_X2 U832 ( .A1(n824), .A2(n1131), .A3(n1130), .ZN(n1421) );
  NAND2_X2 U833 ( .A1(n1129), .A2(n1128), .ZN(n1130) );
  NOR2_X2 U834 ( .A1(n1260), .A2(n1127), .ZN(n1125) );
  INV_X4 U835 ( .A(n958), .ZN(n1770) );
  NAND2_X2 U836 ( .A1(n810), .A2(n1408), .ZN(n1193) );
  NAND3_X2 U837 ( .A1(n1001), .A2(n1000), .A3(n999), .ZN(n1531) );
  AOI21_X2 U838 ( .B1(n1474), .B2(n2138), .A(n839), .ZN(n988) );
  NOR2_X2 U839 ( .A1(n1912), .A2(n1856), .ZN(n1303) );
  NOR2_X2 U840 ( .A1(n2106), .A2(n800), .ZN(n1304) );
  INV_X4 U841 ( .A(n1849), .ZN(n832) );
  INV_X4 U842 ( .A(n1973), .ZN(n1979) );
  OAI21_X2 U843 ( .B1(n1607), .B2(n1703), .A(n1606), .ZN(n1033) );
  INV_X4 U844 ( .A(n783), .ZN(n1864) );
  OAI21_X2 U845 ( .B1(n1607), .B2(n1635), .A(n1606), .ZN(n1034) );
  INV_X4 U846 ( .A(n833), .ZN(n1868) );
  AOI21_X2 U847 ( .B1(n1052), .B2(n1591), .A(n1051), .ZN(n1053) );
  AOI21_X2 U848 ( .B1(n805), .B2(n2134), .A(n1063), .ZN(n1051) );
  NOR2_X2 U849 ( .A1(n843), .A2(n1519), .ZN(n1524) );
  NOR2_X2 U850 ( .A1(n843), .A2(n1550), .ZN(n1555) );
  NOR2_X2 U851 ( .A1(n1961), .A2(n843), .ZN(n1964) );
  INV_X4 U852 ( .A(n2170), .ZN(n2124) );
  INV_X8 U853 ( .A(aluCtrl[1]), .ZN(n1092) );
  INV_X4 U854 ( .A(n1119), .ZN(n1137) );
  OAI21_X2 U855 ( .B1(n1423), .B2(n1133), .A(n1100), .ZN(n1118) );
  AOI22_X2 U856 ( .A1(n789), .A2(n1886), .B1(n786), .B2(n1875), .ZN(n978) );
  NOR2_X2 U857 ( .A1(n989), .A2(n1470), .ZN(n990) );
  INV_X8 U858 ( .A(n997), .ZN(n839) );
  INV_X4 U859 ( .A(n973), .ZN(n1474) );
  NAND3_X2 U860 ( .A1(n1149), .A2(n1288), .A3(n794), .ZN(n1292) );
  NOR2_X2 U861 ( .A1(n1221), .A2(n1218), .ZN(n1149) );
  NOR2_X2 U862 ( .A1(aluCtrl[2]), .A2(aluCtrl[3]), .ZN(n954) );
  NOR2_X2 U863 ( .A1(n1494), .A2(n1493), .ZN(n1495) );
  NOR2_X2 U864 ( .A1(n2156), .A2(n1491), .ZN(n1496) );
  NOR2_X2 U865 ( .A1(n1498), .A2(n1499), .ZN(n1504) );
  OAI21_X2 U866 ( .B1(n1284), .B2(n1283), .A(n1282), .ZN(n1286) );
  NOR3_X1 U867 ( .A1(n1281), .A2(n1280), .A3(n1279), .ZN(n1284) );
  NAND3_X2 U868 ( .A1(n1838), .A2(n1837), .A3(n1836), .ZN(n1892) );
  NOR2_X2 U869 ( .A1(n1835), .A2(n1834), .ZN(n1836) );
  AOI21_X2 U870 ( .B1(n1425), .B2(n1424), .A(n1423), .ZN(n1426) );
  AOI21_X2 U871 ( .B1(n785), .B2(n2031), .A(n846), .ZN(n2033) );
  AOI21_X2 U872 ( .B1(n785), .B2(n2048), .A(n848), .ZN(n2050) );
  NOR2_X2 U873 ( .A1(n2067), .A2(n850), .ZN(n2069) );
  OAI21_X2 U874 ( .B1(n846), .B2(n2066), .A(n2067), .ZN(n2071) );
  OAI21_X2 U875 ( .B1(n1411), .B2(n1410), .A(n1409), .ZN(n1435) );
  AOI21_X2 U876 ( .B1(n785), .B2(n2081), .A(n846), .ZN(n2083) );
  NOR2_X2 U877 ( .A1(n1063), .A2(n972), .ZN(n975) );
  AOI21_X2 U878 ( .B1(n785), .B2(n2098), .A(n848), .ZN(n2100) );
  AOI21_X2 U879 ( .B1(n1433), .B2(n1198), .A(n787), .ZN(n1199) );
  NOR2_X2 U880 ( .A1(n1219), .A2(n1218), .ZN(n1224) );
  NOR2_X2 U881 ( .A1(aluCtrl[0]), .A2(aluCtrl[2]), .ZN(n1004) );
  AOI21_X2 U882 ( .B1(n1061), .B2(n1041), .A(n1040), .ZN(n1042) );
  NOR2_X2 U883 ( .A1(n1345), .A2(n1346), .ZN(n1062) );
  OAI21_X2 U884 ( .B1(n2097), .B2(n1529), .A(n1076), .ZN(n1077) );
  INV_X8 U885 ( .A(n1520), .ZN(n1526) );
  NOR2_X2 U886 ( .A1(n1522), .A2(n1521), .ZN(n1523) );
  OAI21_X2 U887 ( .B1(n1383), .B2(n1382), .A(n1381), .ZN(n1385) );
  NOR2_X2 U888 ( .A1(n1553), .A2(n1552), .ZN(n1554) );
  NOR2_X2 U889 ( .A1(n843), .A2(n1578), .ZN(n1583) );
  NOR2_X2 U890 ( .A1(n1581), .A2(n1580), .ZN(n1582) );
  AOI21_X2 U891 ( .B1(n785), .B2(n1579), .A(n846), .ZN(n1581) );
  NOR2_X2 U892 ( .A1(n2020), .A2(n843), .ZN(n1616) );
  NOR2_X2 U893 ( .A1(n1614), .A2(n1613), .ZN(n1615) );
  AOI21_X2 U894 ( .B1(n785), .B2(n1612), .A(n846), .ZN(n1614) );
  AOI21_X2 U895 ( .B1(n1369), .B2(n1368), .A(n1367), .ZN(n1371) );
  AOI21_X2 U896 ( .B1(n1378), .B2(n1364), .A(n1362), .ZN(n1369) );
  NOR2_X2 U897 ( .A1(n2019), .A2(n843), .ZN(n1646) );
  NOR2_X2 U898 ( .A1(n1644), .A2(n1643), .ZN(n1645) );
  AOI21_X2 U899 ( .B1(n785), .B2(n1642), .A(n848), .ZN(n1644) );
  NOR2_X2 U900 ( .A1(n2000), .A2(n843), .ZN(n1680) );
  NOR2_X2 U901 ( .A1(n1678), .A2(n1677), .ZN(n1679) );
  AOI21_X2 U902 ( .B1(n785), .B2(n1676), .A(n848), .ZN(n1678) );
  NAND3_X2 U903 ( .A1(n1641), .A2(n1640), .A3(n1639), .ZN(n1683) );
  NOR2_X2 U904 ( .A1(n1684), .A2(n1788), .ZN(n1685) );
  NOR2_X2 U905 ( .A1(n184), .A2(n853), .ZN(n1686) );
  NOR2_X2 U906 ( .A1(n1981), .A2(n843), .ZN(n1715) );
  NOR2_X2 U907 ( .A1(n1713), .A2(n1712), .ZN(n1714) );
  AOI21_X2 U908 ( .B1(n785), .B2(n1711), .A(n848), .ZN(n1713) );
  INV_X4 U909 ( .A(n1744), .ZN(n1750) );
  NOR2_X2 U910 ( .A1(n1966), .A2(n843), .ZN(n1748) );
  NOR2_X2 U911 ( .A1(n1746), .A2(n1745), .ZN(n1747) );
  INV_X4 U912 ( .A(n1780), .ZN(n1786) );
  NOR2_X2 U913 ( .A1(n1937), .A2(n843), .ZN(n1784) );
  NOR2_X2 U914 ( .A1(n1782), .A2(n1781), .ZN(n1783) );
  NOR2_X2 U915 ( .A1(n1789), .A2(n1788), .ZN(n1790) );
  NOR2_X2 U916 ( .A1(n1947), .A2(n2170), .ZN(n1823) );
  NOR2_X2 U917 ( .A1(n1900), .A2(n2157), .ZN(n1822) );
  INV_X4 U918 ( .A(n1807), .ZN(n1813) );
  NOR2_X2 U919 ( .A1(n1927), .A2(n843), .ZN(n1811) );
  NOR2_X2 U920 ( .A1(n1809), .A2(n1808), .ZN(n1810) );
  AOI21_X2 U921 ( .B1(n785), .B2(n1807), .A(n848), .ZN(n1809) );
  NAND3_X2 U922 ( .A1(n1779), .A2(n1778), .A3(n1777), .ZN(n1814) );
  AOI21_X2 U923 ( .B1(n1862), .B2(n1831), .A(n1776), .ZN(n1777) );
  NOR2_X2 U924 ( .A1(n1909), .A2(n843), .ZN(n1843) );
  NAND3_X2 U925 ( .A1(n1806), .A2(n1805), .A3(n1804), .ZN(n1846) );
  AOI21_X2 U926 ( .B1(n1862), .B2(n1865), .A(n1803), .ZN(n1804) );
  OAI21_X2 U927 ( .B1(aluSrc), .B2(n889), .A(n888), .ZN(n1879) );
  NOR2_X2 U928 ( .A1(n1909), .A2(n2151), .ZN(n1877) );
  AOI21_X2 U929 ( .B1(n843), .B2(n2157), .A(n796), .ZN(n1873) );
  OAI21_X2 U930 ( .B1(n850), .B2(n1879), .A(n847), .ZN(n1874) );
  NOR2_X2 U931 ( .A1(n843), .A2(n1888), .ZN(n1889) );
  AOI21_X2 U932 ( .B1(n2151), .B2(n2170), .A(n796), .ZN(n1884) );
  OAI21_X2 U933 ( .B1(n1891), .B2(n851), .A(n847), .ZN(n1885) );
  NOR2_X2 U934 ( .A1(n1909), .A2(n2170), .ZN(n1911) );
  NOR2_X2 U935 ( .A1(n1927), .A2(n2157), .ZN(n1910) );
  AOI211_X2 U936 ( .C1(n1907), .C2(n1906), .A(n1905), .B(n1904), .ZN(n1916) );
  NOR2_X2 U937 ( .A1(n1903), .A2(n1902), .ZN(n1904) );
  NOR2_X2 U938 ( .A1(n1900), .A2(n843), .ZN(n1905) );
  NOR2_X2 U939 ( .A1(n1927), .A2(n2170), .ZN(n1929) );
  NOR2_X2 U940 ( .A1(n1937), .A2(n2157), .ZN(n1928) );
  AOI211_X2 U941 ( .C1(n1925), .C2(n1924), .A(n1923), .B(n1922), .ZN(n1934) );
  NOR2_X2 U942 ( .A1(n1921), .A2(n1920), .ZN(n1922) );
  NOR2_X2 U943 ( .A1(n1947), .A2(n843), .ZN(n1923) );
  NOR2_X2 U944 ( .A1(n1966), .A2(n2157), .ZN(n1938) );
  NOR2_X2 U945 ( .A1(n1937), .A2(n2170), .ZN(n1939) );
  NOR3_X2 U946 ( .A1(n1950), .A2(n1949), .A3(n1948), .ZN(n1951) );
  NOR2_X2 U947 ( .A1(n1947), .A2(n2151), .ZN(n1948) );
  NOR2_X2 U948 ( .A1(n1962), .A2(n843), .ZN(n1949) );
  NOR2_X2 U949 ( .A1(n1962), .A2(n2151), .ZN(n1963) );
  OAI21_X2 U950 ( .B1(n846), .B2(n1958), .A(n1957), .ZN(n1959) );
  OAI21_X2 U951 ( .B1(n846), .B2(n1955), .A(n1956), .ZN(n1960) );
  NOR2_X2 U952 ( .A1(n1956), .A2(n850), .ZN(n1958) );
  NOR2_X2 U953 ( .A1(n1726), .A2(n1725), .ZN(n1727) );
  NOR2_X2 U954 ( .A1(n1724), .A2(n833), .ZN(n1726) );
  NOR2_X2 U955 ( .A1(n2000), .A2(n2157), .ZN(n1982) );
  NOR2_X2 U956 ( .A1(n1981), .A2(n2170), .ZN(n1983) );
  NOR2_X2 U957 ( .A1(n1975), .A2(n1974), .ZN(n1976) );
  NOR2_X2 U958 ( .A1(n843), .A2(n1972), .ZN(n1977) );
  NAND3_X2 U959 ( .A1(n1695), .A2(n1694), .A3(n1693), .ZN(n1999) );
  NOR2_X2 U960 ( .A1(n2000), .A2(n2170), .ZN(n2002) );
  NOR2_X2 U961 ( .A1(n2019), .A2(n2157), .ZN(n2001) );
  AOI211_X2 U962 ( .C1(n1998), .C2(n1997), .A(n1996), .B(n1995), .ZN(n2007) );
  NOR2_X2 U963 ( .A1(n1994), .A2(n1993), .ZN(n1995) );
  NOR2_X2 U964 ( .A1(n843), .A2(n1991), .ZN(n1996) );
  NOR2_X2 U965 ( .A1(n1312), .A2(n1413), .ZN(n1313) );
  NAND3_X2 U966 ( .A1(n1661), .A2(n1660), .A3(n1659), .ZN(n2018) );
  NOR2_X2 U967 ( .A1(n1658), .A2(n1657), .ZN(n1659) );
  NOR2_X2 U968 ( .A1(n2020), .A2(n2157), .ZN(n2021) );
  NOR2_X2 U969 ( .A1(n2019), .A2(n2170), .ZN(n2022) );
  AOI211_X2 U970 ( .C1(n2017), .C2(n2016), .A(n2015), .B(n2014), .ZN(n2027) );
  NOR2_X2 U971 ( .A1(n2013), .A2(n2012), .ZN(n2014) );
  NOR2_X2 U972 ( .A1(n843), .A2(n2010), .ZN(n2015) );
  NAND3_X2 U973 ( .A1(n1627), .A2(n1626), .A3(n1625), .ZN(n2038) );
  NOR2_X2 U974 ( .A1(n1624), .A2(n1623), .ZN(n1625) );
  NAND3_X2 U975 ( .A1(n1598), .A2(n1597), .A3(n1596), .ZN(n2055) );
  NOR2_X2 U976 ( .A1(n1595), .A2(n1594), .ZN(n1596) );
  NAND3_X2 U977 ( .A1(n1549), .A2(n1548), .A3(n1547), .ZN(n2063) );
  AOI21_X2 U978 ( .B1(n1605), .B2(n1862), .A(n802), .ZN(n1547) );
  NAND3_X2 U979 ( .A1(n1075), .A2(n1074), .A3(n1073), .ZN(n2088) );
  NOR2_X2 U980 ( .A1(n1072), .A2(n1071), .ZN(n1073) );
  NAND3_X2 U981 ( .A1(n1518), .A2(n1517), .A3(n1516), .ZN(n2089) );
  AOI21_X2 U982 ( .B1(n1573), .B2(n1862), .A(n802), .ZN(n1516) );
  AOI21_X2 U983 ( .B1(n1672), .B2(n1868), .A(n801), .ZN(n1049) );
  INV_X4 U984 ( .A(n2157), .ZN(n2108) );
  OAI21_X2 U985 ( .B1(n846), .B2(n2118), .A(n2117), .ZN(n2119) );
  OAI21_X2 U986 ( .B1(n846), .B2(n2115), .A(n2116), .ZN(n2120) );
  NOR2_X2 U987 ( .A1(n2116), .A2(n850), .ZN(n2118) );
  OAI21_X2 U988 ( .B1(n2140), .B2(n2157), .A(n2125), .ZN(n2126) );
  NOR3_X2 U989 ( .A1(n2168), .A2(n2167), .A3(n2166), .ZN(n2169) );
  NOR2_X2 U990 ( .A1(n2157), .A2(n2156), .ZN(n2168) );
  NOR2_X2 U991 ( .A1(n2159), .A2(n847), .ZN(n2167) );
  NOR3_X2 U992 ( .A1(n1585), .A2(n793), .A3(n1618), .ZN(n1391) );
  NOR2_X2 U993 ( .A1(n795), .A2(n788), .ZN(n1392) );
  OAI21_X2 U994 ( .B1(n1107), .B2(n827), .A(n1321), .ZN(n1134) );
  NAND2_X2 U995 ( .A1(n930), .A2(n1092), .ZN(n994) );
  NAND2_X2 U996 ( .A1(n930), .A2(aluCtrl[1]), .ZN(n995) );
  OAI21_X2 U997 ( .B1(n1503), .B2(n835), .A(n1471), .ZN(n1166) );
  NAND2_X2 U998 ( .A1(n1351), .A2(n1353), .ZN(n1156) );
  NAND2_X2 U999 ( .A1(n1257), .A2(n1278), .ZN(n1277) );
  NOR2_X2 U1000 ( .A1(n1832), .A2(n833), .ZN(n1835) );
  NOR2_X2 U1001 ( .A1(n1833), .A2(n783), .ZN(n1834) );
  NOR2_X2 U1002 ( .A1(n1239), .A2(n1238), .ZN(n1240) );
  OAI21_X2 U1003 ( .B1(aluCtrl[1]), .B2(n1458), .A(n962), .ZN(n1376) );
  OAI21_X2 U1004 ( .B1(n1607), .B2(n1687), .A(n1606), .ZN(n1802) );
  OAI21_X2 U1005 ( .B1(n1592), .B2(n1591), .A(n1590), .ZN(n1593) );
  INV_X4 U1006 ( .A(n1180), .ZN(n1331) );
  NAND3_X2 U1007 ( .A1(n1339), .A2(n1343), .A3(n1344), .ZN(n1180) );
  OAI21_X2 U1008 ( .B1(n1607), .B2(n1720), .A(n1606), .ZN(n1775) );
  NOR2_X2 U1009 ( .A1(n1470), .A2(n971), .ZN(n976) );
  OAI21_X2 U1010 ( .B1(n2099), .B2(n973), .A(n837), .ZN(n974) );
  OAI21_X2 U1011 ( .B1(aluSrc), .B2(n893), .A(n892), .ZN(n2161) );
  NOR2_X2 U1012 ( .A1(n1481), .A2(n784), .ZN(n1482) );
  NAND3_X2 U1013 ( .A1(n1477), .A2(n1476), .A3(n1475), .ZN(n1485) );
  AOI21_X2 U1014 ( .B1(n1474), .B2(n2162), .A(n839), .ZN(n1475) );
  INV_X4 U1015 ( .A(n834), .ZN(n835) );
  OAI21_X2 U1016 ( .B1(n2133), .B2(n807), .A(n1059), .ZN(n1039) );
  NOR3_X2 U1017 ( .A1(n1346), .A2(n1382), .A3(n1345), .ZN(n1386) );
  OAI21_X2 U1018 ( .B1(n1058), .B2(n1057), .A(n1056), .ZN(n1380) );
  NAND2_X2 U1019 ( .A1(n1544), .A2(n1151), .ZN(n1364) );
  NAND3_X2 U1020 ( .A1(n1365), .A2(n1364), .A3(n1363), .ZN(n1368) );
  OAI21_X2 U1021 ( .B1(n1174), .B2(n1381), .A(n1387), .ZN(n1175) );
  NOR2_X2 U1022 ( .A1(n798), .A2(n1775), .ZN(n1776) );
  NAND3_X2 U1023 ( .A1(n1671), .A2(n1773), .A3(n1670), .ZN(n1865) );
  NOR2_X2 U1024 ( .A1(n798), .A2(n1802), .ZN(n1803) );
  OAI21_X2 U1025 ( .B1(n1268), .B2(n1267), .A(n1266), .ZN(n1269) );
  NAND3_X2 U1026 ( .A1(n1774), .A2(n1773), .A3(n1772), .ZN(n1848) );
  NAND3_X2 U1027 ( .A1(n1705), .A2(n1773), .A3(n1704), .ZN(n1847) );
  OAI22_X2 U1028 ( .A1(n1260), .A2(n1112), .B1(n1111), .B2(n1260), .ZN(n1113)
         );
  NAND3_X2 U1029 ( .A1(n1738), .A2(n1773), .A3(n1737), .ZN(n1861) );
  NAND3_X2 U1030 ( .A1(n1755), .A2(n1773), .A3(n1754), .ZN(n1863) );
  OAI21_X2 U1031 ( .B1(n846), .B2(n1940), .A(n1941), .ZN(n1945) );
  OAI21_X2 U1032 ( .B1(n846), .B2(n1943), .A(n1942), .ZN(n1944) );
  NOR2_X2 U1033 ( .A1(n1941), .A2(n850), .ZN(n1943) );
  NAND3_X2 U1034 ( .A1(n1247), .A2(n1132), .A3(n1421), .ZN(n1139) );
  NAND3_X2 U1035 ( .A1(n1656), .A2(n1655), .A3(n1654), .ZN(n1850) );
  NAND3_X2 U1036 ( .A1(n1722), .A2(n1773), .A3(n1721), .ZN(n1851) );
  NOR2_X2 U1037 ( .A1(n1795), .A2(n783), .ZN(n1725) );
  NAND3_X2 U1038 ( .A1(n1561), .A2(n1655), .A3(n1560), .ZN(n1691) );
  NAND3_X2 U1039 ( .A1(n1622), .A2(n1655), .A3(n1621), .ZN(n1817) );
  NAND3_X2 U1040 ( .A1(n1690), .A2(n1773), .A3(n1689), .ZN(n1867) );
  AOI21_X2 U1041 ( .B1(n785), .B2(n1992), .A(n846), .ZN(n1994) );
  NOR2_X2 U1042 ( .A1(n1795), .A2(n784), .ZN(n1657) );
  NOR2_X2 U1043 ( .A1(n1794), .A2(n798), .ZN(n1658) );
  NAND3_X2 U1044 ( .A1(n1535), .A2(n1655), .A3(n1534), .ZN(n1649) );
  AOI21_X2 U1045 ( .B1(n785), .B2(n2011), .A(n848), .ZN(n2013) );
  NOR2_X2 U1046 ( .A1(n1762), .A2(n784), .ZN(n1623) );
  NOR2_X2 U1047 ( .A1(n1761), .A2(n798), .ZN(n1624) );
  NOR2_X2 U1048 ( .A1(n1795), .A2(n798), .ZN(n1594) );
  NOR2_X2 U1049 ( .A1(n1724), .A2(n784), .ZN(n1595) );
  NOR2_X2 U1050 ( .A1(n1481), .A2(n833), .ZN(n1071) );
  NOR2_X2 U1051 ( .A1(n1069), .A2(n784), .ZN(n1072) );
  NAND3_X2 U1052 ( .A1(n1068), .A2(n1655), .A3(n1067), .ZN(n1692) );
  NAND3_X2 U1053 ( .A1(n1019), .A2(n1655), .A3(n1018), .ZN(n1650) );
  OAI21_X2 U1054 ( .B1(n1607), .B2(n1736), .A(n1606), .ZN(n1046) );
  AOI211_X2 U1055 ( .C1(n1017), .C2(n1591), .A(n991), .B(n990), .ZN(n992) );
  NAND3_X2 U1056 ( .A1(n936), .A2(n935), .A3(n934), .ZN(n1070) );
  INV_X4 U1057 ( .A(n798), .ZN(n1866) );
  AOI22_X2 U1058 ( .A1(n1299), .A2(n1298), .B1(n1297), .B2(n1296), .ZN(n1301)
         );
  NOR2_X2 U1059 ( .A1(n1293), .A2(n1292), .ZN(n1298) );
  AOI21_X2 U1060 ( .B1(n2162), .B2(n2161), .A(n2160), .ZN(n2164) );
  NOR2_X2 U1061 ( .A1(n1490), .A2(n1489), .ZN(n1509) );
  AOI21_X2 U1062 ( .B1(n1507), .B2(n1506), .A(n809), .ZN(n1508) );
  AOI211_X2 U1063 ( .C1(n2143), .C2(n1497), .A(n1496), .B(n1495), .ZN(n1507)
         );
  NOR3_X2 U1064 ( .A1(n1466), .A2(fp), .A3(n1465), .ZN(n1467) );
  AOI21_X2 U1065 ( .B1(n1058), .B2(n1011), .A(n1010), .ZN(n1012) );
  OAI21_X2 U1066 ( .B1(n2133), .B2(n806), .A(n1478), .ZN(n1009) );
  AOI211_X2 U1067 ( .C1(n2037), .C2(n2036), .A(n2035), .B(n2034), .ZN(n2044)
         );
  NOR2_X2 U1068 ( .A1(n2033), .A2(n2032), .ZN(n2034) );
  NOR2_X2 U1069 ( .A1(n843), .A2(n2030), .ZN(n2035) );
  AOI211_X2 U1070 ( .C1(n2054), .C2(n2053), .A(n2052), .B(n2051), .ZN(n2061)
         );
  NOR2_X2 U1071 ( .A1(n2050), .A2(n2049), .ZN(n2051) );
  NOR2_X2 U1072 ( .A1(n2065), .A2(n843), .ZN(n2052) );
  NOR2_X2 U1073 ( .A1(n2073), .A2(n2072), .ZN(n2074) );
  OAI21_X2 U1074 ( .B1(n846), .B2(n2069), .A(n2068), .ZN(n2070) );
  AOI21_X2 U1075 ( .B1(n1435), .B2(n1434), .A(n1227), .ZN(n1436) );
  AOI211_X2 U1076 ( .C1(n2087), .C2(n2086), .A(n2085), .B(n2084), .ZN(n2094)
         );
  NOR2_X2 U1077 ( .A1(n2083), .A2(n2082), .ZN(n2084) );
  NOR2_X2 U1078 ( .A1(n2080), .A2(n2151), .ZN(n2085) );
  OAI21_X2 U1079 ( .B1(n1231), .B2(n787), .A(n1230), .ZN(n1232) );
  AOI21_X2 U1080 ( .B1(n1229), .B2(n1228), .A(n1227), .ZN(n1231) );
  AOI21_X2 U1081 ( .B1(n1638), .B2(n1868), .A(n801), .ZN(n1036) );
  AOI211_X2 U1082 ( .C1(n2104), .C2(n2103), .A(n2102), .B(n2101), .ZN(n2112)
         );
  NOR2_X2 U1083 ( .A1(n2100), .A2(n2099), .ZN(n2101) );
  NOR2_X2 U1084 ( .A1(n2097), .A2(n2151), .ZN(n2102) );
  OAI21_X2 U1085 ( .B1(n2133), .B2(n2132), .A(n2136), .ZN(n2147) );
  OAI21_X2 U1086 ( .B1(n2136), .B2(n2135), .A(n2134), .ZN(n2137) );
  NOR2_X2 U1087 ( .A1(n194), .A2(n195), .ZN(isZero) );
  NOR2_X2 U1088 ( .A1(n1375), .A2(n1493), .ZN(n1078) );
  AOI211_X2 U1089 ( .C1(n1526), .C2(n1525), .A(n1524), .B(n1523), .ZN(n1543)
         );
  AOI211_X2 U1090 ( .C1(n1557), .C2(n1556), .A(n1555), .B(n1554), .ZN(n1570)
         );
  AOI211_X2 U1091 ( .C1(n925), .C2(n1584), .A(n1583), .B(n1582), .ZN(n1602) );
  AOI211_X2 U1092 ( .C1(n924), .C2(n1617), .A(n1616), .B(n1615), .ZN(n1631) );
  AOI211_X2 U1093 ( .C1(n1648), .C2(n1647), .A(n1646), .B(n1645), .ZN(n1665)
         );
  NOR2_X2 U1094 ( .A1(n1686), .A2(n1685), .ZN(n1697) );
  AOI211_X2 U1095 ( .C1(n1682), .C2(n1681), .A(n1680), .B(n1679), .ZN(n1699)
         );
  AOI211_X2 U1096 ( .C1(n1717), .C2(n1716), .A(n1715), .B(n1714), .ZN(n1732)
         );
  AOI211_X2 U1097 ( .C1(n1750), .C2(n1749), .A(n1748), .B(n1747), .ZN(n1766)
         );
  NOR2_X2 U1098 ( .A1(n812), .A2(n1790), .ZN(n1797) );
  AOI211_X2 U1099 ( .C1(n1813), .C2(n1812), .A(n1811), .B(n1810), .ZN(n1828)
         );
  NOR2_X2 U1100 ( .A1(n1823), .A2(n1822), .ZN(n1826) );
  AOI211_X2 U1101 ( .C1(n1845), .C2(n1844), .A(n1843), .B(n1842), .ZN(n1860)
         );
  AOI21_X2 U1102 ( .B1(n1875), .B2(n1874), .A(n1873), .ZN(n1883) );
  AOI21_X2 U1103 ( .B1(n1879), .B2(n1878), .A(n1877), .ZN(n1882) );
  AOI21_X2 U1104 ( .B1(n1886), .B2(n1885), .A(n1884), .ZN(n1897) );
  AOI21_X2 U1105 ( .B1(n1891), .B2(n1890), .A(n1889), .ZN(n1896) );
  NOR2_X2 U1106 ( .A1(n1911), .A2(n1910), .ZN(n1914) );
  NOR2_X2 U1107 ( .A1(n1929), .A2(n1928), .ZN(n1932) );
  NOR2_X2 U1108 ( .A1(n1939), .A2(n1938), .ZN(n1952) );
  AOI211_X2 U1109 ( .C1(n852), .C2(n790), .A(n1967), .B(n808), .ZN(n1968) );
  NOR3_X2 U1110 ( .A1(n1965), .A2(n1964), .A3(n1963), .ZN(n1969) );
  NOR2_X2 U1111 ( .A1(n1983), .A2(n1982), .ZN(n1986) );
  NOR2_X2 U1112 ( .A1(n2002), .A2(n2001), .ZN(n2005) );
  NOR2_X2 U1113 ( .A1(n2022), .A2(n2021), .ZN(n2025) );
  NOR2_X2 U1114 ( .A1(n2122), .A2(n2121), .ZN(n2129) );
  AOI21_X2 U1115 ( .B1(n852), .B2(n2173), .A(n2172), .ZN(n2178) );
  OAI21_X2 U1116 ( .B1(n2171), .B2(n2170), .A(n2169), .ZN(n2172) );
  INV_X4 U1117 ( .A(n995), .ZN(n830) );
  OAI21_X2 U1118 ( .B1(n1607), .B2(n1669), .A(n1606), .ZN(n1047) );
  NAND2_X1 U1119 ( .A1(n799), .A2(n1669), .ZN(n1670) );
  INV_X4 U1120 ( .A(n784), .ZN(n1862) );
  NAND2_X2 U1121 ( .A1(n1478), .A2(n1027), .ZN(n783) );
  NAND2_X2 U1122 ( .A1(n1002), .A2(n1059), .ZN(n784) );
  AND2_X4 U1123 ( .A1(n2131), .A2(n853), .ZN(n785) );
  AND2_X4 U1124 ( .A1(n828), .A2(n1520), .ZN(n786) );
  XOR2_X2 U1125 ( .A(n1197), .B(n2082), .Z(n787) );
  XOR2_X2 U1126 ( .A(n1342), .B(n1341), .Z(n788) );
  NAND2_X2 U1127 ( .A1(n2141), .A2(n853), .ZN(n2170) );
  INV_X4 U1128 ( .A(n785), .ZN(n850) );
  INV_X4 U1129 ( .A(n2158), .ZN(n848) );
  INV_X4 U1130 ( .A(n848), .ZN(n847) );
  INV_X1 U1131 ( .A(n1276), .ZN(n825) );
  AND2_X4 U1132 ( .A1(n830), .A2(n1520), .ZN(n789) );
  XOR2_X2 U1133 ( .A(n1340), .B(n1339), .Z(n790) );
  XOR2_X2 U1134 ( .A(n1191), .B(n2012), .Z(n791) );
  XOR2_X2 U1135 ( .A(n1388), .B(n1387), .Z(n792) );
  XOR2_X2 U1136 ( .A(n1361), .B(n1360), .Z(n793) );
  AND2_X4 U1137 ( .A1(n1405), .A2(n803), .ZN(n794) );
  XOR2_X1 U1138 ( .A(n1419), .B(n820), .Z(n795) );
  AND4_X4 U1139 ( .A1(n1872), .A2(n1871), .A3(n1870), .A4(n1869), .ZN(n796) );
  INV_X4 U1140 ( .A(zeroExt), .ZN(n955) );
  OR2_X4 U1141 ( .A1(n992), .A2(n833), .ZN(n797) );
  INV_X4 U1142 ( .A(n834), .ZN(n842) );
  INV_X8 U1143 ( .A(n842), .ZN(n840) );
  NAND2_X2 U1144 ( .A1(n1478), .A2(n1059), .ZN(n798) );
  INV_X4 U1145 ( .A(n2151), .ZN(n845) );
  AND2_X4 U1146 ( .A1(n1520), .A2(n1591), .ZN(n799) );
  XOR2_X2 U1147 ( .A(n1259), .B(n1265), .Z(n800) );
  AND2_X4 U1148 ( .A1(n2160), .A2(n1059), .ZN(n801) );
  AND2_X4 U1149 ( .A1(n1866), .A2(n2160), .ZN(n802) );
  AND2_X4 U1150 ( .A1(n1407), .A2(n1400), .ZN(n803) );
  AND2_X4 U1151 ( .A1(n954), .A2(aluCtrl[1]), .ZN(n804) );
  INV_X4 U1152 ( .A(n2113), .ZN(n844) );
  INV_X4 U1153 ( .A(n844), .ZN(n843) );
  INV_X4 U1154 ( .A(n828), .ZN(n829) );
  INV_X4 U1155 ( .A(n994), .ZN(n828) );
  OR2_X4 U1156 ( .A1(n1591), .A2(n2135), .ZN(n805) );
  INV_X4 U1157 ( .A(fp), .ZN(n853) );
  AND2_X4 U1158 ( .A1(n2131), .A2(n1008), .ZN(n806) );
  AND2_X4 U1159 ( .A1(n2131), .A2(n1038), .ZN(n807) );
  INV_X4 U1160 ( .A(n2163), .ZN(n849) );
  INV_X4 U1161 ( .A(n1376), .ZN(n834) );
  AND2_X4 U1162 ( .A1(busA[20]), .A2(fp), .ZN(n808) );
  AND2_X4 U1163 ( .A1(n1505), .A2(fp), .ZN(n809) );
  AND2_X4 U1164 ( .A1(n1407), .A2(n1409), .ZN(n810) );
  NAND2_X2 U1165 ( .A1(n1530), .A2(n853), .ZN(n2157) );
  OR2_X4 U1166 ( .A1(n1021), .A2(n784), .ZN(n811) );
  AND2_X4 U1167 ( .A1(busA[12]), .A2(fp), .ZN(n812) );
  INV_X8 U1168 ( .A(zeroExt), .ZN(n836) );
  OR3_X4 U1169 ( .A1(n1216), .A2(aluCtrl[0]), .A3(fp), .ZN(n813) );
  INV_X4 U1170 ( .A(n1788), .ZN(n852) );
  AND2_X4 U1171 ( .A1(busA[29]), .A2(fp), .ZN(n814) );
  INV_X4 U1172 ( .A(n785), .ZN(n851) );
  OR2_X4 U1173 ( .A1(n2154), .A2(n2153), .ZN(aluRes[30]) );
  INV_X4 U1174 ( .A(n832), .ZN(n833) );
  INV_X4 U1175 ( .A(n2158), .ZN(n846) );
  NAND2_X2 U1176 ( .A1(n1135), .A2(n1320), .ZN(n1322) );
  NAND2_X4 U1177 ( .A1(n1235), .A2(n1354), .ZN(n1245) );
  OAI21_X2 U1178 ( .B1(n1242), .B2(n1241), .A(n1240), .ZN(n1244) );
  AOI21_X1 U1179 ( .B1(n785), .B2(n1919), .A(n846), .ZN(n1921) );
  INV_X4 U1180 ( .A(n1919), .ZN(n1925) );
  XNOR2_X2 U1181 ( .A(n1188), .B(n834), .ZN(n816) );
  INV_X2 U1182 ( .A(n1419), .ZN(n1318) );
  OAI21_X2 U1183 ( .B1(n1607), .B2(n1753), .A(n1606), .ZN(n1546) );
  OAI221_X2 U1184 ( .B1(n831), .B2(n1552), .C1(n829), .C2(n1195), .A(n838), 
        .ZN(n1753) );
  OAI21_X2 U1185 ( .B1(n1453), .B2(n1454), .A(n1457), .ZN(n1450) );
  NOR2_X1 U1186 ( .A1(n1226), .A2(n1225), .ZN(n1229) );
  INV_X4 U1187 ( .A(n1193), .ZN(n1226) );
  INV_X4 U1188 ( .A(n1551), .ZN(n817) );
  INV_X4 U1189 ( .A(n817), .ZN(n818) );
  AOI21_X1 U1190 ( .B1(n785), .B2(n1839), .A(n848), .ZN(n1841) );
  NAND2_X1 U1191 ( .A1(n1408), .A2(n1407), .ZN(n1441) );
  NAND2_X1 U1192 ( .A1(n794), .A2(n1440), .ZN(n1442) );
  INV_X2 U1193 ( .A(n1440), .ZN(n1432) );
  INV_X2 U1194 ( .A(n1089), .ZN(n1886) );
  OAI221_X1 U1195 ( .B1(n829), .B2(n1089), .C1(n831), .C2(n1084), .A(n837), 
        .ZN(n1688) );
  NAND2_X1 U1196 ( .A1(n1311), .A2(n1310), .ZN(n1314) );
  NAND3_X2 U1197 ( .A1(n1400), .A2(n1399), .A3(n1398), .ZN(n1402) );
  OAI21_X1 U1198 ( .B1(n1307), .B2(n1413), .A(n1311), .ZN(n1309) );
  AOI211_X4 U1199 ( .C1(n1485), .C2(n1484), .A(n1483), .B(n1482), .ZN(n1487)
         );
  NAND2_X1 U1200 ( .A1(n1295), .A2(n1294), .ZN(n1296) );
  OAI211_X4 U1201 ( .C1(n1246), .C2(n1245), .A(n1244), .B(n1243), .ZN(n1342)
         );
  INV_X4 U1202 ( .A(n1418), .ZN(n819) );
  INV_X8 U1203 ( .A(n819), .ZN(n820) );
  NOR2_X2 U1204 ( .A1(n1841), .A2(n1840), .ZN(n1842) );
  OAI221_X1 U1205 ( .B1(n831), .B2(n1840), .C1(n829), .C2(n1902), .A(n837), 
        .ZN(n1719) );
  INV_X2 U1206 ( .A(n1840), .ZN(n1829) );
  INV_X1 U1207 ( .A(n2155), .ZN(n2173) );
  NAND2_X1 U1208 ( .A1(n1917), .A2(n1098), .ZN(n1132) );
  INV_X4 U1209 ( .A(n1652), .ZN(n821) );
  INV_X4 U1210 ( .A(n821), .ZN(n822) );
  OAI21_X1 U1211 ( .B1(n1280), .B2(n825), .A(n1265), .ZN(n1283) );
  XNOR2_X2 U1212 ( .A(n1813), .B(n1154), .ZN(n1101) );
  NAND2_X1 U1213 ( .A1(n1868), .A2(n1562), .ZN(n1564) );
  NAND2_X1 U1214 ( .A1(n1864), .A2(n1562), .ZN(n1075) );
  INV_X4 U1215 ( .A(n931), .ZN(n930) );
  NAND2_X2 U1216 ( .A1(n1331), .A2(n1330), .ZN(n1217) );
  INV_X4 U1217 ( .A(n1420), .ZN(n823) );
  INV_X8 U1218 ( .A(n823), .ZN(n824) );
  AOI21_X1 U1219 ( .B1(n785), .B2(n1520), .A(n846), .ZN(n1522) );
  XNOR2_X1 U1220 ( .A(n1173), .B(n1520), .ZN(n1387) );
  OAI21_X1 U1221 ( .B1(n1607), .B2(n1771), .A(n1606), .ZN(n1515) );
  NAND2_X1 U1222 ( .A1(n799), .A2(n1771), .ZN(n1772) );
  XNOR2_X2 U1223 ( .A(n1161), .B(n1632), .ZN(n826) );
  INV_X4 U1224 ( .A(n826), .ZN(n1360) );
  NAND2_X1 U1225 ( .A1(busA[8]), .A2(n836), .ZN(n1643) );
  OAI221_X1 U1226 ( .B1(n829), .B2(n1920), .C1(n831), .C2(n1808), .A(n838), 
        .ZN(n1752) );
  OAI221_X1 U1227 ( .B1(n829), .B2(n2099), .C1(n831), .C2(n1063), .A(n838), 
        .ZN(n1736) );
  XNOR2_X2 U1228 ( .A(n1097), .B(n841), .ZN(n827) );
  INV_X4 U1229 ( .A(n842), .ZN(n841) );
  OAI21_X2 U1230 ( .B1(n1260), .B2(n1251), .A(n1319), .ZN(n1106) );
  NAND3_X1 U1231 ( .A1(n1349), .A2(n1348), .A3(n1387), .ZN(n1363) );
  NAND2_X4 U1232 ( .A1(n1172), .A2(n1348), .ZN(n1359) );
  INV_X4 U1233 ( .A(n1437), .ZN(n1443) );
  AOI22_X1 U1234 ( .A1(busA[27]), .A2(fp), .B1(n852), .B2(n2090), .ZN(n2091)
         );
  NOR3_X2 U1235 ( .A1(n1446), .A2(n2090), .A3(n2057), .ZN(n1447) );
  XNOR2_X1 U1236 ( .A(n1277), .B(n1276), .ZN(n1856) );
  NOR3_X2 U1237 ( .A1(n1893), .A2(n2127), .A3(n2149), .ZN(n1302) );
  NAND2_X1 U1238 ( .A1(n852), .A2(n2149), .ZN(n2150) );
  NAND3_X2 U1239 ( .A1(n1456), .A2(n1457), .A3(n1455), .ZN(n1463) );
  NOR2_X1 U1240 ( .A1(n1459), .A2(n1458), .ZN(n1461) );
  AOI211_X1 U1241 ( .C1(n1979), .C2(n1978), .A(n1977), .B(n1976), .ZN(n1988)
         );
  AOI21_X1 U1242 ( .B1(n785), .B2(n1973), .A(n846), .ZN(n1975) );
  XNOR2_X1 U1243 ( .A(n1979), .B(n841), .ZN(n1147) );
  NAND3_X4 U1244 ( .A1(n1250), .A2(n1108), .A3(n1266), .ZN(n1091) );
  NAND2_X4 U1245 ( .A1(n1088), .A2(n1282), .ZN(n1108) );
  AOI22_X1 U1246 ( .A1(busA[13]), .A2(fp), .B1(n852), .B2(n1824), .ZN(n1825)
         );
  AOI222_X2 U1247 ( .A1(n1587), .A2(n1070), .B1(n1479), .B2(n1002), .C1(n1866), 
        .C2(n1619), .ZN(n2152) );
  OAI211_X1 U1248 ( .C1(n1359), .C2(n1358), .A(n1357), .B(n1356), .ZN(n1361)
         );
  OAI21_X1 U1249 ( .B1(n1026), .B2(n1025), .A(n1170), .ZN(n1029) );
  NAND2_X4 U1250 ( .A1(n1118), .A2(n1117), .ZN(n1119) );
  NAND3_X4 U1251 ( .A1(n979), .A2(n838), .A3(n978), .ZN(n1651) );
  NAND3_X4 U1252 ( .A1(n957), .A2(n956), .A3(n838), .ZN(n1635) );
  NAND2_X1 U1253 ( .A1(n828), .A2(n2162), .ZN(n956) );
  NAND3_X2 U1254 ( .A1(n1176), .A2(n1160), .A3(n1370), .ZN(n1357) );
  NOR2_X4 U1255 ( .A1(n1163), .A2(n1162), .ZN(n1179) );
  NAND2_X4 U1256 ( .A1(n1404), .A2(n1401), .ZN(n1408) );
  INV_X1 U1257 ( .A(n2142), .ZN(n1014) );
  AOI21_X1 U1258 ( .B1(n785), .B2(n1901), .A(n846), .ZN(n1903) );
  INV_X4 U1259 ( .A(n2142), .ZN(n1486) );
  INV_X2 U1260 ( .A(n1901), .ZN(n1907) );
  NAND3_X2 U1261 ( .A1(n1901), .A2(n1102), .A3(n1919), .ZN(n884) );
  INV_X8 U1262 ( .A(n1171), .ZN(n1382) );
  OAI21_X1 U1263 ( .B1(n1062), .B2(n1380), .A(n1171), .ZN(n1065) );
  NAND3_X2 U1264 ( .A1(n820), .A2(n1419), .A3(n1256), .ZN(n1254) );
  NAND2_X4 U1265 ( .A1(n1061), .A2(n1060), .ZN(n1171) );
  XNOR2_X1 U1266 ( .A(n1552), .B(n1154), .ZN(n1155) );
  OAI22_X4 U1267 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n1154) );
  NAND2_X4 U1268 ( .A1(n816), .A2(n1220), .ZN(n1311) );
  AOI211_X1 U1269 ( .C1(n1786), .C2(n1785), .A(n1784), .B(n1783), .ZN(n1799)
         );
  OAI21_X2 U1270 ( .B1(n1327), .B2(n827), .A(n1326), .ZN(n1329) );
  NAND2_X1 U1271 ( .A1(n1134), .A2(n1133), .ZN(n1136) );
  XNOR2_X1 U1272 ( .A(n1786), .B(n840), .ZN(n1105) );
  NAND3_X2 U1273 ( .A1(n1264), .A2(n1282), .A3(n1253), .ZN(n1110) );
  NAND3_X2 U1274 ( .A1(n1282), .A2(n1276), .A3(n1264), .ZN(n1109) );
  OAI21_X2 U1275 ( .B1(n1464), .B2(n1463), .A(n1462), .ZN(n1468) );
  NAND3_X1 U1276 ( .A1(n1271), .A2(n1328), .A3(n1270), .ZN(n1272) );
  NAND3_X1 U1277 ( .A1(n1338), .A2(n1337), .A3(n1336), .ZN(n1340) );
  INV_X8 U1278 ( .A(n1337), .ZN(n1142) );
  XNOR2_X1 U1279 ( .A(n925), .B(n1154), .ZN(n1153) );
  NAND2_X4 U1280 ( .A1(n1226), .A2(n1433), .ZN(n1200) );
  INV_X32 U1281 ( .A(aluCtrl[0]), .ZN(n1458) );
  AOI21_X1 U1282 ( .B1(n785), .B2(n1744), .A(n848), .ZN(n1746) );
  INV_X1 U1283 ( .A(n1413), .ZN(n1299) );
  NAND3_X1 U1284 ( .A1(n824), .A2(n1419), .A3(n820), .ZN(n1422) );
  INV_X2 U1285 ( .A(n820), .ZN(n1317) );
  NAND2_X4 U1286 ( .A1(n820), .A2(n824), .ZN(n1115) );
  NAND3_X2 U1287 ( .A1(n1676), .A2(n1744), .A3(n1711), .ZN(n885) );
  OAI21_X4 U1288 ( .B1(n1443), .B2(n1208), .A(n1207), .ZN(n1209) );
  OAI211_X4 U1289 ( .C1(n1206), .C2(n1297), .A(n1205), .B(n1204), .ZN(n1207)
         );
  AOI22_X1 U1290 ( .A1(busA[23]), .A2(fp), .B1(n852), .B2(n2023), .ZN(n2024)
         );
  AOI21_X1 U1291 ( .B1(n785), .B2(n1780), .A(n846), .ZN(n1782) );
  NAND2_X1 U1292 ( .A1(n1973), .A2(n1780), .ZN(n882) );
  OAI21_X1 U1293 ( .B1(n1443), .B2(n1442), .A(n1441), .ZN(n1445) );
  NAND2_X1 U1294 ( .A1(n822), .A2(n1066), .ZN(n1068) );
  NAND2_X1 U1295 ( .A1(n822), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1296 ( .A1(n822), .A2(n1651), .ZN(n1656) );
  NAND2_X1 U1297 ( .A1(n822), .A2(n1533), .ZN(n1535) );
  NAND2_X1 U1298 ( .A1(n822), .A2(n1559), .ZN(n1561) );
  NAND2_X1 U1299 ( .A1(n822), .A2(n1620), .ZN(n1622) );
  XNOR2_X1 U1300 ( .A(n1344), .B(n1343), .ZN(n1684) );
  OAI21_X1 U1301 ( .B1(n1386), .B2(n1385), .A(n1384), .ZN(n1388) );
  OAI21_X1 U1302 ( .B1(n1386), .B2(n1347), .A(n1384), .ZN(n1349) );
  NAND2_X4 U1303 ( .A1(n1179), .A2(n1178), .ZN(n1344) );
  NAND2_X1 U1304 ( .A1(n1526), .A2(n822), .ZN(n1470) );
  INV_X2 U1305 ( .A(n1384), .ZN(n1174) );
  NAND3_X2 U1306 ( .A1(n1384), .A2(n1171), .A3(n1380), .ZN(n1348) );
  NAND2_X1 U1307 ( .A1(n1520), .A2(n822), .ZN(n958) );
  AOI21_X1 U1308 ( .B1(n785), .B2(n818), .A(n846), .ZN(n1553) );
  NAND2_X1 U1309 ( .A1(n2143), .A2(n2142), .ZN(n2144) );
  OAI221_X1 U1310 ( .B1(n1478), .B2(n1022), .C1(n1021), .C2(n783), .A(n1020), 
        .ZN(n2105) );
  OAI211_X4 U1311 ( .C1(n1002), .C2(n1022), .A(n797), .B(n811), .ZN(n2142) );
  AOI21_X1 U1312 ( .B1(n1460), .B2(n1458), .A(n1306), .ZN(n1451) );
  AOI21_X1 U1313 ( .B1(n1461), .B2(n1460), .A(setInv), .ZN(n1462) );
  NAND2_X1 U1314 ( .A1(n1331), .A2(n1330), .ZN(n1440) );
  NAND2_X1 U1315 ( .A1(n1002), .A2(n1027), .ZN(n1849) );
  INV_X8 U1316 ( .A(n1027), .ZN(n1059) );
  NAND2_X4 U1317 ( .A1(n1114), .A2(n1113), .ZN(n1320) );
  NAND3_X1 U1318 ( .A1(n1342), .A2(n1335), .A3(n1334), .ZN(n1338) );
  INV_X8 U1319 ( .A(n1460), .ZN(n1457) );
  NAND2_X4 U1320 ( .A1(n2155), .A2(n2165), .ZN(n1460) );
  INV_X2 U1321 ( .A(n1453), .ZN(n1456) );
  OAI21_X1 U1322 ( .B1(n1413), .B2(n1287), .A(n1232), .ZN(n1234) );
  OAI21_X1 U1323 ( .B1(n1413), .B2(n1290), .A(n1295), .ZN(n1291) );
  OAI21_X1 U1324 ( .B1(n1413), .B2(n1402), .A(n1401), .ZN(n1403) );
  OAI21_X1 U1325 ( .B1(n1413), .B2(n1412), .A(n1435), .ZN(n1414) );
  NAND3_X1 U1326 ( .A1(n1440), .A2(n1428), .A3(n1437), .ZN(n1332) );
  XNOR2_X1 U1327 ( .A(n1416), .B(n1415), .ZN(n1789) );
  AOI21_X1 U1328 ( .B1(n1438), .B2(n1437), .A(n1436), .ZN(n1439) );
  NAND3_X1 U1329 ( .A1(n820), .A2(n1419), .A3(n1415), .ZN(n1263) );
  AOI21_X1 U1330 ( .B1(n1261), .B2(n1415), .A(n1260), .ZN(n1262) );
  NAND3_X1 U1331 ( .A1(n1415), .A2(n1320), .A3(n1319), .ZN(n1323) );
  OAI21_X1 U1332 ( .B1(n1251), .B2(n1415), .A(n1250), .ZN(n1252) );
  NAND2_X4 U1333 ( .A1(n1217), .A2(n1437), .ZN(n1413) );
  INV_X4 U1334 ( .A(busB[1]), .ZN(n855) );
  INV_X4 U1335 ( .A(imm32[1]), .ZN(n854) );
  MUX2_X2 U1336 ( .A(n855), .B(n854), .S(aluSrc), .Z(n1002) );
  INV_X4 U1337 ( .A(n1002), .ZN(n1478) );
  INV_X4 U1338 ( .A(busB[2]), .ZN(n857) );
  INV_X4 U1339 ( .A(imm32[2]), .ZN(n856) );
  MUX2_X2 U1340 ( .A(n857), .B(n856), .S(aluSrc), .Z(n1027) );
  INV_X4 U1341 ( .A(busB[4]), .ZN(n859) );
  INV_X4 U1342 ( .A(imm32[4]), .ZN(n858) );
  MUX2_X2 U1343 ( .A(n859), .B(n858), .S(aluSrc), .Z(n1520) );
  INV_X4 U1344 ( .A(busB[3]), .ZN(n861) );
  INV_X4 U1345 ( .A(imm32[3]), .ZN(n860) );
  MUX2_X2 U1346 ( .A(n861), .B(n860), .S(aluSrc), .Z(n1652) );
  INV_X4 U1347 ( .A(n1470), .ZN(n993) );
  INV_X4 U1348 ( .A(busB[9]), .ZN(n863) );
  INV_X4 U1349 ( .A(imm32[9]), .ZN(n862) );
  MUX2_X2 U1350 ( .A(n863), .B(n862), .S(aluSrc), .Z(n1676) );
  INV_X4 U1351 ( .A(busB[11]), .ZN(n865) );
  INV_X4 U1352 ( .A(imm32[11]), .ZN(n864) );
  MUX2_X2 U1353 ( .A(n865), .B(n864), .S(aluSrc), .Z(n1744) );
  INV_X4 U1354 ( .A(busB[10]), .ZN(n867) );
  INV_X4 U1355 ( .A(imm32[10]), .ZN(n866) );
  MUX2_X2 U1356 ( .A(n867), .B(n866), .S(aluSrc), .Z(n1711) );
  INV_X4 U1357 ( .A(busB[17]), .ZN(n869) );
  INV_X4 U1358 ( .A(imm32[17]), .ZN(n868) );
  MUX2_X2 U1359 ( .A(n869), .B(n868), .S(aluSrc), .Z(n1901) );
  INV_X4 U1360 ( .A(busB[16]), .ZN(n871) );
  INV_X4 U1361 ( .A(imm32[16]), .ZN(n870) );
  MUX2_X2 U1362 ( .A(n871), .B(n870), .S(aluSrc), .Z(n1102) );
  INV_X4 U1363 ( .A(busB[18]), .ZN(n873) );
  INV_X4 U1364 ( .A(imm32[18]), .ZN(n872) );
  MUX2_X2 U1365 ( .A(n873), .B(n872), .S(aluSrc), .Z(n1919) );
  INV_X4 U1366 ( .A(busB[22]), .ZN(n875) );
  INV_X4 U1367 ( .A(imm32[22]), .ZN(n874) );
  MUX2_X2 U1368 ( .A(n875), .B(n874), .S(aluSrc), .Z(n1992) );
  INV_X4 U1369 ( .A(busB[20]), .ZN(n877) );
  INV_X4 U1370 ( .A(imm32[20]), .ZN(n876) );
  MUX2_X2 U1371 ( .A(n877), .B(n876), .S(aluSrc), .Z(n1140) );
  NAND2_X2 U1372 ( .A1(n1992), .A2(n1140), .ZN(n883) );
  INV_X4 U1373 ( .A(busB[21]), .ZN(n879) );
  INV_X4 U1374 ( .A(imm32[21]), .ZN(n878) );
  MUX2_X2 U1375 ( .A(n879), .B(n878), .S(aluSrc), .Z(n1973) );
  INV_X4 U1376 ( .A(busB[12]), .ZN(n881) );
  INV_X4 U1377 ( .A(imm32[12]), .ZN(n880) );
  MUX2_X2 U1378 ( .A(n881), .B(n880), .S(aluSrc), .Z(n1780) );
  NOR4_X2 U1379 ( .A1(n885), .A2(n884), .A3(n883), .A4(n882), .ZN(n929) );
  INV_X4 U1380 ( .A(busB[13]), .ZN(n887) );
  INV_X4 U1381 ( .A(imm32[13]), .ZN(n886) );
  MUX2_X2 U1382 ( .A(n887), .B(n886), .S(aluSrc), .Z(n1807) );
  INV_X4 U1383 ( .A(busB[15]), .ZN(n889) );
  NAND2_X2 U1384 ( .A1(imm32[15]), .A2(aluSrc), .ZN(n888) );
  INV_X4 U1385 ( .A(busB[14]), .ZN(n891) );
  INV_X4 U1386 ( .A(imm32[14]), .ZN(n890) );
  MUX2_X2 U1387 ( .A(n891), .B(n890), .S(aluSrc), .Z(n1839) );
  INV_X4 U1388 ( .A(n1839), .ZN(n1845) );
  INV_X4 U1389 ( .A(busB[31]), .ZN(n893) );
  NAND2_X2 U1390 ( .A1(imm32[31]), .A2(aluSrc), .ZN(n892) );
  NOR4_X2 U1391 ( .A1(n1813), .A2(n1879), .A3(n1845), .A4(n2161), .ZN(n928) );
  INV_X4 U1392 ( .A(busB[8]), .ZN(n895) );
  INV_X4 U1393 ( .A(imm32[8]), .ZN(n894) );
  MUX2_X2 U1394 ( .A(n895), .B(n894), .S(aluSrc), .Z(n1642) );
  INV_X4 U1395 ( .A(busB[30]), .ZN(n897) );
  INV_X4 U1396 ( .A(imm32[30]), .ZN(n896) );
  MUX2_X2 U1397 ( .A(n897), .B(n896), .S(aluSrc), .Z(n1145) );
  INV_X4 U1398 ( .A(busB[5]), .ZN(n899) );
  INV_X4 U1399 ( .A(imm32[5]), .ZN(n898) );
  MUX2_X2 U1400 ( .A(n899), .B(n898), .S(aluSrc), .Z(n1551) );
  NAND3_X4 U1401 ( .A1(n1642), .A2(n1145), .A3(n818), .ZN(n917) );
  INV_X4 U1402 ( .A(busB[24]), .ZN(n901) );
  INV_X4 U1403 ( .A(imm32[24]), .ZN(n900) );
  MUX2_X2 U1404 ( .A(n901), .B(n900), .S(aluSrc), .Z(n2031) );
  INV_X4 U1405 ( .A(busB[23]), .ZN(n903) );
  INV_X4 U1406 ( .A(imm32[23]), .ZN(n902) );
  MUX2_X2 U1407 ( .A(n903), .B(n902), .S(aluSrc), .Z(n2011) );
  INV_X4 U1408 ( .A(busB[25]), .ZN(n905) );
  INV_X4 U1409 ( .A(imm32[25]), .ZN(n904) );
  MUX2_X2 U1410 ( .A(n905), .B(n904), .S(aluSrc), .Z(n2048) );
  NAND3_X4 U1411 ( .A1(n2031), .A2(n2011), .A3(n2048), .ZN(n916) );
  INV_X4 U1412 ( .A(busB[29]), .ZN(n907) );
  INV_X4 U1413 ( .A(imm32[29]), .ZN(n906) );
  MUX2_X2 U1414 ( .A(n907), .B(n906), .S(aluSrc), .Z(n1144) );
  INV_X4 U1415 ( .A(busB[27]), .ZN(n909) );
  INV_X4 U1416 ( .A(imm32[27]), .ZN(n908) );
  MUX2_X2 U1417 ( .A(n909), .B(n908), .S(aluSrc), .Z(n2081) );
  NAND2_X2 U1418 ( .A1(n1144), .A2(n2081), .ZN(n915) );
  INV_X4 U1419 ( .A(busB[28]), .ZN(n911) );
  INV_X4 U1420 ( .A(imm32[28]), .ZN(n910) );
  MUX2_X2 U1421 ( .A(n911), .B(n910), .S(aluSrc), .Z(n2098) );
  INV_X4 U1422 ( .A(busB[19]), .ZN(n913) );
  INV_X4 U1423 ( .A(imm32[19]), .ZN(n912) );
  MUX2_X2 U1424 ( .A(n913), .B(n912), .S(aluSrc), .Z(n1081) );
  NAND2_X2 U1425 ( .A1(n2098), .A2(n1081), .ZN(n914) );
  NOR4_X2 U1426 ( .A1(n917), .A2(n916), .A3(n915), .A4(n914), .ZN(n927) );
  INV_X4 U1427 ( .A(busB[6]), .ZN(n919) );
  INV_X4 U1428 ( .A(imm32[6]), .ZN(n918) );
  MUX2_X2 U1429 ( .A(n919), .B(n918), .S(aluSrc), .Z(n1579) );
  INV_X4 U1430 ( .A(n1579), .ZN(n925) );
  INV_X4 U1431 ( .A(busB[7]), .ZN(n921) );
  INV_X4 U1432 ( .A(imm32[7]), .ZN(n920) );
  MUX2_X2 U1433 ( .A(n921), .B(n920), .S(aluSrc), .Z(n1612) );
  INV_X4 U1434 ( .A(n1612), .ZN(n924) );
  INV_X4 U1435 ( .A(busB[26]), .ZN(n923) );
  INV_X4 U1436 ( .A(imm32[26]), .ZN(n922) );
  MUX2_X2 U1437 ( .A(n923), .B(n922), .S(aluSrc), .Z(n1146) );
  NAND4_X2 U1438 ( .A1(n929), .A2(n928), .A3(n927), .A4(n926), .ZN(n931) );
  NAND2_X2 U1439 ( .A1(busA[20]), .A2(n955), .ZN(n1141) );
  NAND2_X2 U1440 ( .A1(busA[11]), .A2(n955), .ZN(n1745) );
  NAND2_X2 U1441 ( .A1(busA[31]), .A2(n836), .ZN(n1080) );
  INV_X4 U1442 ( .A(n1080), .ZN(n2162) );
  NAND2_X2 U1443 ( .A1(aluCtrl[0]), .A2(n2162), .ZN(n2156) );
  INV_X4 U1444 ( .A(n2156), .ZN(n2160) );
  NAND2_X2 U1445 ( .A1(n2160), .A2(n931), .ZN(n997) );
  OAI221_X2 U1446 ( .B1(n829), .B2(n1141), .C1(n831), .C2(n1745), .A(n837), 
        .ZN(n1735) );
  NAND2_X2 U1447 ( .A1(n993), .A2(n1735), .ZN(n936) );
  NAND2_X2 U1448 ( .A1(busA[28]), .A2(n955), .ZN(n2099) );
  NAND2_X2 U1449 ( .A1(busA[3]), .A2(n836), .ZN(n1063) );
  NAND2_X2 U1450 ( .A1(n1736), .A2(n1526), .ZN(n933) );
  NAND2_X2 U1451 ( .A1(busA[12]), .A2(n836), .ZN(n1781) );
  INV_X4 U1452 ( .A(n1781), .ZN(n1767) );
  NAND2_X2 U1453 ( .A1(busA[19]), .A2(n955), .ZN(n1120) );
  INV_X4 U1454 ( .A(n1120), .ZN(n1942) );
  AOI22_X2 U1455 ( .A1(n786), .A2(n1767), .B1(n789), .B2(n1942), .ZN(n932) );
  NAND3_X2 U1456 ( .A1(n933), .A2(n838), .A3(n932), .ZN(n1559) );
  NAND2_X2 U1457 ( .A1(n1559), .A2(n1591), .ZN(n935) );
  NAND2_X2 U1458 ( .A1(n1770), .A2(n830), .ZN(n973) );
  NAND2_X2 U1459 ( .A1(busA[27]), .A2(n955), .ZN(n2082) );
  INV_X4 U1460 ( .A(n2082), .ZN(n2078) );
  NAND2_X2 U1461 ( .A1(n1770), .A2(n828), .ZN(n972) );
  INV_X4 U1462 ( .A(n972), .ZN(n1472) );
  NAND2_X2 U1463 ( .A1(busA[4]), .A2(n955), .ZN(n1521) );
  INV_X4 U1464 ( .A(n1521), .ZN(n1513) );
  AOI221_X2 U1465 ( .B1(n1474), .B2(n2078), .C1(n1472), .C2(n1513), .A(n839), 
        .ZN(n934) );
  NAND2_X2 U1466 ( .A1(busA[5]), .A2(n836), .ZN(n1552) );
  NAND2_X2 U1467 ( .A1(busA[26]), .A2(n836), .ZN(n1195) );
  NAND2_X2 U1468 ( .A1(n1753), .A2(n1526), .ZN(n938) );
  NAND2_X2 U1469 ( .A1(busA[21]), .A2(n836), .ZN(n1974) );
  INV_X4 U1470 ( .A(n1974), .ZN(n1970) );
  NAND2_X2 U1471 ( .A1(busA[10]), .A2(n836), .ZN(n1712) );
  INV_X4 U1472 ( .A(n1712), .ZN(n1700) );
  AOI22_X2 U1473 ( .A1(n789), .A2(n1970), .B1(n786), .B2(n1700), .ZN(n937) );
  NAND3_X2 U1474 ( .A1(n938), .A2(n838), .A3(n937), .ZN(n1066) );
  NAND2_X2 U1475 ( .A1(n1066), .A2(n1591), .ZN(n941) );
  NAND2_X2 U1476 ( .A1(busA[18]), .A2(n836), .ZN(n1920) );
  NAND2_X2 U1477 ( .A1(busA[13]), .A2(n836), .ZN(n1808) );
  NAND2_X2 U1478 ( .A1(n993), .A2(n1752), .ZN(n940) );
  NAND2_X2 U1479 ( .A1(busA[2]), .A2(n836), .ZN(n1038) );
  INV_X4 U1480 ( .A(n1038), .ZN(n1061) );
  NAND2_X2 U1481 ( .A1(busA[29]), .A2(n836), .ZN(n1184) );
  INV_X4 U1482 ( .A(n1184), .ZN(n2117) );
  AOI22_X2 U1483 ( .A1(n1472), .A2(n1061), .B1(n1474), .B2(n2117), .ZN(n939)
         );
  NAND4_X2 U1484 ( .A1(n941), .A2(n837), .A3(n940), .A4(n939), .ZN(n947) );
  NAND2_X2 U1485 ( .A1(busA[30]), .A2(n836), .ZN(n1182) );
  NAND2_X2 U1486 ( .A1(busA[1]), .A2(n836), .ZN(n1008) );
  OAI221_X2 U1487 ( .B1(n829), .B2(n1182), .C1(n831), .C2(n1008), .A(n837), 
        .ZN(n1669) );
  NAND2_X2 U1488 ( .A1(n1669), .A2(n1526), .ZN(n943) );
  NAND2_X2 U1489 ( .A1(busA[14]), .A2(n836), .ZN(n1840) );
  NAND2_X2 U1490 ( .A1(busA[17]), .A2(n836), .ZN(n1902) );
  INV_X4 U1491 ( .A(n1902), .ZN(n1898) );
  AOI22_X2 U1492 ( .A1(n786), .A2(n1829), .B1(n789), .B2(n1898), .ZN(n942) );
  NAND3_X2 U1493 ( .A1(n943), .A2(n838), .A3(n942), .ZN(n1620) );
  NAND2_X2 U1494 ( .A1(n1620), .A2(n1591), .ZN(n946) );
  NAND2_X2 U1495 ( .A1(busA[22]), .A2(n836), .ZN(n1993) );
  NAND2_X2 U1496 ( .A1(busA[9]), .A2(n955), .ZN(n1677) );
  OAI221_X2 U1497 ( .B1(n829), .B2(n1993), .C1(n831), .C2(n1677), .A(n837), 
        .ZN(n1668) );
  NAND2_X2 U1498 ( .A1(n993), .A2(n1668), .ZN(n945) );
  NAND2_X2 U1499 ( .A1(busA[6]), .A2(n836), .ZN(n1580) );
  INV_X4 U1500 ( .A(n1580), .ZN(n1571) );
  NAND2_X2 U1501 ( .A1(busA[25]), .A2(n955), .ZN(n2049) );
  INV_X4 U1502 ( .A(n2049), .ZN(n2045) );
  AOI22_X2 U1503 ( .A1(n1472), .A2(n1571), .B1(n1474), .B2(n2045), .ZN(n944)
         );
  NAND4_X2 U1504 ( .A1(n946), .A2(n837), .A3(n945), .A4(n944), .ZN(n1562) );
  MUX2_X2 U1505 ( .A(n947), .B(n1562), .S(n1059), .Z(n1479) );
  NAND2_X2 U1506 ( .A1(busA[7]), .A2(n836), .ZN(n1613) );
  NAND2_X2 U1507 ( .A1(busA[24]), .A2(n836), .ZN(n2032) );
  OAI221_X2 U1508 ( .B1(n831), .B2(n1613), .C1(n829), .C2(n2032), .A(n837), 
        .ZN(n1687) );
  NAND2_X2 U1509 ( .A1(n1687), .A2(n1526), .ZN(n949) );
  INV_X4 U1510 ( .A(n1643), .ZN(n1632) );
  NAND2_X2 U1511 ( .A1(busA[23]), .A2(n836), .ZN(n2012) );
  INV_X4 U1512 ( .A(n2012), .ZN(n2008) );
  AOI22_X2 U1513 ( .A1(n786), .A2(n1632), .B1(n789), .B2(n2008), .ZN(n948) );
  NAND3_X2 U1514 ( .A1(n949), .A2(n838), .A3(n948), .ZN(n1473) );
  INV_X4 U1515 ( .A(n1473), .ZN(n951) );
  NAND2_X2 U1516 ( .A1(busA[16]), .A2(n955), .ZN(n1089) );
  NAND2_X2 U1517 ( .A1(busA[15]), .A2(n955), .ZN(n1084) );
  NAND2_X2 U1518 ( .A1(n799), .A2(n1688), .ZN(n950) );
  NAND2_X2 U1519 ( .A1(n2160), .A2(n1526), .ZN(n1773) );
  INV_X4 U1520 ( .A(n1773), .ZN(n1634) );
  NAND2_X2 U1521 ( .A1(n1634), .A2(n1591), .ZN(n1655) );
  OAI211_X2 U1522 ( .C1(n951), .C2(n1591), .A(n950), .B(n1655), .ZN(n1619) );
  NAND2_X2 U1523 ( .A1(n954), .A2(n1092), .ZN(n1489) );
  INV_X4 U1524 ( .A(n1489), .ZN(n1003) );
  INV_X4 U1525 ( .A(busB[0]), .ZN(n953) );
  INV_X4 U1526 ( .A(imm32[0]), .ZN(n952) );
  MUX2_X2 U1527 ( .A(n953), .B(n952), .S(aluSrc), .Z(n1500) );
  INV_X4 U1528 ( .A(n1500), .ZN(n1503) );
  NAND2_X2 U1529 ( .A1(n1003), .A2(n1503), .ZN(n1529) );
  NAND2_X2 U1530 ( .A1(n804), .A2(n1503), .ZN(n1491) );
  INV_X4 U1531 ( .A(n1491), .ZN(n1527) );
  NAND2_X2 U1532 ( .A1(n2160), .A2(n958), .ZN(n959) );
  INV_X4 U1533 ( .A(n959), .ZN(n1607) );
  NAND2_X2 U1534 ( .A1(busA[0]), .A2(n836), .ZN(n1499) );
  INV_X4 U1535 ( .A(n1499), .ZN(n1471) );
  NAND2_X2 U1536 ( .A1(n830), .A2(n1471), .ZN(n957) );
  NAND2_X2 U1537 ( .A1(n959), .A2(n958), .ZN(n1606) );
  MUX2_X2 U1538 ( .A(n2156), .B(n1034), .S(n1868), .Z(n2171) );
  INV_X4 U1539 ( .A(n2171), .ZN(n1497) );
  NAND2_X2 U1540 ( .A1(n1527), .A2(n1497), .ZN(n967) );
  INV_X4 U1541 ( .A(aluCtrl[3]), .ZN(n962) );
  NAND2_X2 U1542 ( .A1(aluCtrl[2]), .A2(n962), .ZN(n1493) );
  INV_X4 U1543 ( .A(n1493), .ZN(n1528) );
  OAI22_X2 U1544 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n960) );
  XNOR2_X2 U1545 ( .A(n960), .B(n1008), .ZN(n961) );
  XNOR2_X2 U1546 ( .A(n961), .B(n1002), .ZN(n1026) );
  INV_X4 U1547 ( .A(n1026), .ZN(n1057) );
  OAI22_X2 U1548 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n963) );
  XNOR2_X2 U1549 ( .A(n963), .B(n1499), .ZN(n964) );
  XNOR2_X2 U1550 ( .A(n964), .B(n1500), .ZN(n1377) );
  INV_X4 U1551 ( .A(n1377), .ZN(n965) );
  NAND2_X2 U1552 ( .A1(n965), .A2(n835), .ZN(n1169) );
  NAND2_X2 U1553 ( .A1(n1166), .A2(n1169), .ZN(n1346) );
  INV_X4 U1554 ( .A(n1346), .ZN(n1025) );
  XNOR2_X2 U1555 ( .A(n1057), .B(n1025), .ZN(n1372) );
  NAND2_X2 U1556 ( .A1(n1528), .A2(n1372), .ZN(n966) );
  OAI211_X2 U1557 ( .C1(n2152), .C2(n1529), .A(n967), .B(n966), .ZN(n1016) );
  INV_X4 U1558 ( .A(n1141), .ZN(n1957) );
  INV_X4 U1559 ( .A(n1745), .ZN(n1733) );
  AOI22_X2 U1560 ( .A1(n789), .A2(n1957), .B1(n786), .B2(n1733), .ZN(n968) );
  NAND3_X2 U1561 ( .A1(n969), .A2(n838), .A3(n968), .ZN(n1533) );
  NAND2_X2 U1562 ( .A1(n1533), .A2(n1591), .ZN(n970) );
  INV_X4 U1563 ( .A(n970), .ZN(n977) );
  OAI221_X2 U1564 ( .B1(n831), .B2(n1781), .C1(n829), .C2(n1120), .A(n837), 
        .ZN(n1769) );
  INV_X4 U1565 ( .A(n1769), .ZN(n971) );
  NOR4_X2 U1566 ( .A1(n977), .A2(n976), .A3(n975), .A4(n974), .ZN(n984) );
  OAI221_X2 U1567 ( .B1(n831), .B2(n1643), .C1(n829), .C2(n2012), .A(n837), 
        .ZN(n1653) );
  NAND2_X2 U1568 ( .A1(n993), .A2(n1653), .ZN(n982) );
  NAND2_X2 U1569 ( .A1(n1635), .A2(n1526), .ZN(n979) );
  INV_X4 U1570 ( .A(n1084), .ZN(n1875) );
  NAND2_X2 U1571 ( .A1(n1651), .A2(n1591), .ZN(n981) );
  INV_X4 U1572 ( .A(n2032), .ZN(n2028) );
  INV_X4 U1573 ( .A(n1613), .ZN(n1603) );
  AOI221_X2 U1574 ( .B1(n1474), .B2(n2028), .C1(n1472), .C2(n1603), .A(n839), 
        .ZN(n980) );
  NAND3_X4 U1575 ( .A1(n982), .A2(n981), .A3(n980), .ZN(n1586) );
  INV_X4 U1576 ( .A(n1586), .ZN(n983) );
  MUX2_X2 U1577 ( .A(n984), .B(n983), .S(n1059), .Z(n1022) );
  OAI221_X2 U1578 ( .B1(n831), .B2(n1580), .C1(n829), .C2(n2049), .A(n837), 
        .ZN(n1720) );
  NAND2_X2 U1579 ( .A1(n1720), .A2(n1526), .ZN(n986) );
  INV_X4 U1580 ( .A(n1993), .ZN(n1989) );
  INV_X4 U1581 ( .A(n1677), .ZN(n1666) );
  AOI22_X2 U1582 ( .A1(n789), .A2(n1989), .B1(n786), .B2(n1666), .ZN(n985) );
  NAND3_X2 U1583 ( .A1(n986), .A2(n838), .A3(n985), .ZN(n1017) );
  INV_X4 U1584 ( .A(n1182), .ZN(n2138) );
  INV_X4 U1585 ( .A(n1008), .ZN(n1058) );
  NAND2_X2 U1586 ( .A1(n1472), .A2(n1058), .ZN(n987) );
  NAND2_X2 U1587 ( .A1(n988), .A2(n987), .ZN(n991) );
  INV_X4 U1588 ( .A(n1719), .ZN(n989) );
  OAI221_X2 U1589 ( .B1(n829), .B2(n1974), .C1(n831), .C2(n1712), .A(n837), 
        .ZN(n1702) );
  NAND2_X2 U1590 ( .A1(n993), .A2(n1702), .ZN(n1001) );
  OAI221_X2 U1591 ( .B1(n831), .B2(n1038), .C1(n829), .C2(n1184), .A(n837), 
        .ZN(n1703) );
  NAND2_X2 U1592 ( .A1(n1703), .A2(n1526), .ZN(n998) );
  INV_X4 U1593 ( .A(n1920), .ZN(n1917) );
  INV_X4 U1594 ( .A(n1808), .ZN(n1800) );
  AOI22_X2 U1595 ( .A1(n789), .A2(n1917), .B1(n786), .B2(n1800), .ZN(n996) );
  NAND3_X2 U1596 ( .A1(n998), .A2(n838), .A3(n996), .ZN(n1588) );
  NAND2_X2 U1597 ( .A1(n1588), .A2(n1591), .ZN(n1000) );
  INV_X4 U1598 ( .A(n1195), .ZN(n2068) );
  INV_X4 U1599 ( .A(n1552), .ZN(n1544) );
  AOI221_X2 U1600 ( .B1(n1474), .B2(n2068), .C1(n1472), .C2(n1544), .A(n839), 
        .ZN(n999) );
  INV_X4 U1601 ( .A(n1531), .ZN(n1021) );
  NAND2_X2 U1602 ( .A1(n1003), .A2(n1500), .ZN(n2139) );
  NAND2_X2 U1603 ( .A1(n804), .A2(n1500), .ZN(n1054) );
  INV_X4 U1604 ( .A(n1054), .ZN(n2143) );
  MUX2_X2 U1605 ( .A(n2156), .B(n1047), .S(n1868), .Z(n2140) );
  INV_X4 U1606 ( .A(n2140), .ZN(n1023) );
  NAND2_X2 U1607 ( .A1(n2143), .A2(n1023), .ZN(n1013) );
  NAND2_X2 U1608 ( .A1(aluCtrl[1]), .A2(aluCtrl[3]), .ZN(n1216) );
  INV_X4 U1609 ( .A(n1216), .ZN(n1005) );
  NAND2_X2 U1610 ( .A1(n1005), .A2(n1004), .ZN(n2135) );
  NAND2_X2 U1611 ( .A1(aluCtrl[3]), .A2(n1092), .ZN(n1466) );
  INV_X4 U1612 ( .A(n1466), .ZN(n1006) );
  INV_X4 U1613 ( .A(aluCtrl[2]), .ZN(n1465) );
  NAND2_X2 U1614 ( .A1(n1006), .A2(n1465), .ZN(n1498) );
  MUX2_X2 U1615 ( .A(n2135), .B(n1498), .S(n1478), .Z(n1007) );
  INV_X4 U1616 ( .A(n1498), .ZN(n2130) );
  NAND2_X2 U1617 ( .A1(aluCtrl[0]), .A2(n2130), .ZN(n2134) );
  NAND2_X2 U1618 ( .A1(n1007), .A2(n2134), .ZN(n1011) );
  INV_X4 U1619 ( .A(n2134), .ZN(n2133) );
  INV_X4 U1620 ( .A(n2135), .ZN(n2131) );
  INV_X4 U1621 ( .A(n1009), .ZN(n1010) );
  OAI211_X2 U1622 ( .C1(n1014), .C2(n2139), .A(n1013), .B(n1012), .ZN(n1015)
         );
  NOR2_X2 U1623 ( .A1(n1016), .A2(n1015), .ZN(n439) );
  NAND2_X2 U1624 ( .A1(n799), .A2(n1719), .ZN(n1018) );
  NAND2_X2 U1625 ( .A1(n1866), .A2(n1650), .ZN(n1020) );
  INV_X4 U1626 ( .A(n2105), .ZN(n2114) );
  NAND2_X2 U1627 ( .A1(n1527), .A2(n1023), .ZN(n1032) );
  XNOR2_X2 U1628 ( .A(n1478), .B(n840), .ZN(n1024) );
  NAND2_X2 U1629 ( .A1(n1058), .A2(n1024), .ZN(n1170) );
  XNOR2_X2 U1630 ( .A(n1038), .B(n835), .ZN(n1028) );
  XNOR2_X2 U1631 ( .A(n1029), .B(n1056), .ZN(n1374) );
  INV_X4 U1632 ( .A(n1374), .ZN(n1030) );
  NAND2_X2 U1633 ( .A1(n1528), .A2(n1030), .ZN(n1031) );
  OAI211_X2 U1634 ( .C1(n2114), .C2(n1529), .A(n1032), .B(n1031), .ZN(n1045)
         );
  INV_X4 U1635 ( .A(n1033), .ZN(n1638) );
  INV_X4 U1636 ( .A(n1034), .ZN(n1573) );
  NAND2_X2 U1637 ( .A1(n1573), .A2(n1864), .ZN(n1035) );
  NAND2_X2 U1638 ( .A1(n1036), .A2(n1035), .ZN(n2123) );
  INV_X4 U1639 ( .A(n2123), .ZN(n1043) );
  MUX2_X2 U1640 ( .A(n2135), .B(n1498), .S(n1059), .Z(n1037) );
  NAND2_X2 U1641 ( .A1(n1037), .A2(n2134), .ZN(n1041) );
  INV_X4 U1642 ( .A(n1039), .ZN(n1040) );
  OAI221_X2 U1643 ( .B1(n1043), .B2(n1054), .C1(n2152), .C2(n2139), .A(n1042), 
        .ZN(n1044) );
  NOR2_X2 U1644 ( .A1(n1045), .A2(n1044), .ZN(n299) );
  INV_X4 U1645 ( .A(n1046), .ZN(n1672) );
  INV_X4 U1646 ( .A(n1047), .ZN(n1605) );
  NAND2_X2 U1647 ( .A1(n1605), .A2(n1864), .ZN(n1048) );
  NAND2_X2 U1648 ( .A1(n1049), .A2(n1048), .ZN(n2107) );
  INV_X4 U1649 ( .A(n2107), .ZN(n1055) );
  INV_X4 U1650 ( .A(n1063), .ZN(n1165) );
  MUX2_X2 U1651 ( .A(n2135), .B(n1498), .S(n1165), .Z(n1050) );
  NAND2_X2 U1652 ( .A1(n1050), .A2(n2134), .ZN(n1052) );
  OAI221_X2 U1653 ( .B1(n1055), .B2(n1054), .C1(n2114), .C2(n2139), .A(n1053), 
        .ZN(n1079) );
  INV_X4 U1654 ( .A(n1170), .ZN(n1345) );
  XNOR2_X2 U1655 ( .A(n1059), .B(n840), .ZN(n1060) );
  XNOR2_X2 U1656 ( .A(n1063), .B(n835), .ZN(n1064) );
  XNOR2_X2 U1657 ( .A(n1064), .B(n822), .ZN(n1381) );
  XNOR2_X2 U1658 ( .A(n1065), .B(n1381), .ZN(n1375) );
  NAND2_X2 U1659 ( .A1(n799), .A2(n1752), .ZN(n1067) );
  NAND2_X2 U1660 ( .A1(n1866), .A2(n1692), .ZN(n1074) );
  INV_X4 U1661 ( .A(n1619), .ZN(n1069) );
  INV_X4 U1662 ( .A(n1070), .ZN(n1481) );
  INV_X4 U1663 ( .A(n2088), .ZN(n2097) );
  NAND2_X2 U1664 ( .A1(n1527), .A2(n2123), .ZN(n1076) );
  NOR3_X2 U1665 ( .A1(n1079), .A2(n1078), .A3(n1077), .ZN(n267) );
  XNOR2_X2 U1666 ( .A(n1503), .B(n1471), .ZN(n1215) );
  XNOR2_X2 U1667 ( .A(n2161), .B(n1080), .ZN(n1211) );
  XNOR2_X2 U1668 ( .A(n835), .B(n1211), .ZN(n1210) );
  INV_X4 U1669 ( .A(n1081), .ZN(n1941) );
  XNOR2_X2 U1670 ( .A(n1941), .B(n840), .ZN(n1121) );
  NAND2_X2 U1671 ( .A1(n1942), .A2(n1121), .ZN(n1336) );
  INV_X4 U1672 ( .A(n1676), .ZN(n1682) );
  XNOR2_X2 U1673 ( .A(n1682), .B(n840), .ZN(n1150) );
  NAND2_X2 U1674 ( .A1(n1666), .A2(n1150), .ZN(n1243) );
  XNOR2_X2 U1675 ( .A(n1925), .B(n840), .ZN(n1098) );
  INV_X4 U1676 ( .A(n1132), .ZN(n1423) );
  XNOR2_X2 U1677 ( .A(n1907), .B(n840), .ZN(n1082) );
  NAND2_X2 U1678 ( .A1(n1898), .A2(n1082), .ZN(n1321) );
  XNOR2_X2 U1679 ( .A(n1154), .B(n1808), .ZN(n1083) );
  XNOR2_X2 U1680 ( .A(n1083), .B(n1807), .ZN(n1328) );
  INV_X4 U1681 ( .A(n1328), .ZN(n1250) );
  OAI22_X2 U1682 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n1086) );
  XNOR2_X2 U1683 ( .A(n1086), .B(n1084), .ZN(n1085) );
  XNOR2_X2 U1684 ( .A(n1085), .B(n1879), .ZN(n1265) );
  INV_X4 U1685 ( .A(n1265), .ZN(n1088) );
  XNOR2_X2 U1686 ( .A(n1086), .B(n1879), .ZN(n1087) );
  NAND2_X2 U1687 ( .A1(n1875), .A2(n1087), .ZN(n1282) );
  OAI22_X2 U1688 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n1103) );
  XNOR2_X2 U1689 ( .A(n1103), .B(n1089), .ZN(n1090) );
  XNOR2_X2 U1690 ( .A(n1090), .B(n1102), .ZN(n1285) );
  INV_X4 U1691 ( .A(n1285), .ZN(n1266) );
  OAI22_X2 U1692 ( .A1(aluCtrl[3]), .A2(n1092), .B1(aluCtrl[0]), .B2(
        aluCtrl[3]), .ZN(n1094) );
  XNOR2_X2 U1693 ( .A(n1845), .B(n1094), .ZN(n1093) );
  XNOR2_X2 U1694 ( .A(n1094), .B(n1840), .ZN(n1095) );
  XNOR2_X2 U1695 ( .A(n1095), .B(n1839), .ZN(n1276) );
  NAND3_X2 U1696 ( .A1(n1264), .A2(n1282), .A3(n1276), .ZN(n1112) );
  NAND2_X2 U1697 ( .A1(n1111), .A2(n1112), .ZN(n1126) );
  NAND2_X2 U1698 ( .A1(n1321), .A2(n1126), .ZN(n1133) );
  XNOR2_X2 U1699 ( .A(n1902), .B(n835), .ZN(n1096) );
  XNOR2_X2 U1700 ( .A(n1096), .B(n1901), .ZN(n1319) );
  INV_X4 U1701 ( .A(n1319), .ZN(n1107) );
  XNOR2_X2 U1702 ( .A(n1786), .B(n1767), .ZN(n1097) );
  INV_X4 U1703 ( .A(n1134), .ZN(n1099) );
  XNOR2_X2 U1704 ( .A(n1750), .B(n840), .ZN(n1124) );
  XNOR2_X2 U1705 ( .A(n1124), .B(n1745), .ZN(n1418) );
  XNOR2_X2 U1706 ( .A(n1098), .B(n1920), .ZN(n1420) );
  OAI21_X4 U1707 ( .B1(n1099), .B2(n1115), .A(n1132), .ZN(n1100) );
  NAND2_X2 U1708 ( .A1(n1800), .A2(n1101), .ZN(n1253) );
  INV_X4 U1709 ( .A(n1110), .ZN(n1271) );
  INV_X4 U1710 ( .A(n1102), .ZN(n1891) );
  XNOR2_X2 U1711 ( .A(n1891), .B(n1103), .ZN(n1104) );
  NAND2_X2 U1712 ( .A1(n1886), .A2(n1104), .ZN(n1270) );
  INV_X4 U1713 ( .A(n1270), .ZN(n1260) );
  NAND2_X2 U1714 ( .A1(n1767), .A2(n1105), .ZN(n1326) );
  INV_X4 U1715 ( .A(n1326), .ZN(n1251) );
  OAI21_X4 U1716 ( .B1(n1271), .B2(n1107), .A(n1106), .ZN(n1135) );
  NAND4_X2 U1717 ( .A1(n1110), .A2(n1109), .A3(n1108), .A4(n1266), .ZN(n1114)
         );
  INV_X4 U1718 ( .A(n1115), .ZN(n1116) );
  NAND3_X2 U1719 ( .A1(n1135), .A2(n1320), .A3(n1116), .ZN(n1117) );
  XNOR2_X2 U1720 ( .A(n1121), .B(n1120), .ZN(n1417) );
  INV_X4 U1721 ( .A(n1711), .ZN(n1717) );
  XNOR2_X2 U1722 ( .A(n1717), .B(n840), .ZN(n1123) );
  XNOR2_X2 U1723 ( .A(n1123), .B(n1712), .ZN(n1341) );
  NAND2_X2 U1724 ( .A1(n1417), .A2(n1341), .ZN(n1333) );
  OAI21_X4 U1725 ( .B1(n1137), .B2(n1333), .A(n1336), .ZN(n1330) );
  INV_X4 U1726 ( .A(n1330), .ZN(n1122) );
  AOI21_X4 U1727 ( .B1(n1336), .B2(n1243), .A(n1122), .ZN(n1143) );
  NAND2_X2 U1728 ( .A1(n1700), .A2(n1123), .ZN(n1247) );
  NAND2_X2 U1729 ( .A1(n1733), .A2(n1124), .ZN(n1316) );
  NAND2_X2 U1730 ( .A1(n1316), .A2(n1321), .ZN(n1127) );
  NAND3_X2 U1731 ( .A1(n1271), .A2(n1126), .A3(n1125), .ZN(n1131) );
  INV_X4 U1732 ( .A(n1135), .ZN(n1129) );
  INV_X4 U1733 ( .A(n1127), .ZN(n1128) );
  NAND2_X2 U1734 ( .A1(n1136), .A2(n1322), .ZN(n1424) );
  INV_X4 U1735 ( .A(n1424), .ZN(n1138) );
  OAI21_X4 U1736 ( .B1(n1138), .B2(n1421), .A(n1137), .ZN(n1335) );
  NAND3_X4 U1737 ( .A1(n1139), .A2(n1417), .A3(n1335), .ZN(n1337) );
  INV_X4 U1738 ( .A(n1140), .ZN(n1956) );
  XNOR2_X2 U1739 ( .A(n1956), .B(n840), .ZN(n1148) );
  XNOR2_X2 U1740 ( .A(n1148), .B(n1141), .ZN(n1339) );
  OAI21_X4 U1741 ( .B1(n1143), .B2(n1142), .A(n1339), .ZN(n1437) );
  INV_X4 U1742 ( .A(n1144), .ZN(n2116) );
  XNOR2_X2 U1743 ( .A(n2116), .B(n840), .ZN(n1185) );
  NAND2_X2 U1744 ( .A1(n2117), .A2(n1185), .ZN(n1297) );
  INV_X4 U1745 ( .A(n1145), .ZN(n2136) );
  XNOR2_X2 U1746 ( .A(n2136), .B(n840), .ZN(n1183) );
  NAND2_X2 U1747 ( .A1(n2138), .A2(n1183), .ZN(n1204) );
  INV_X4 U1748 ( .A(n1146), .ZN(n2067) );
  XNOR2_X2 U1749 ( .A(n2067), .B(n840), .ZN(n1196) );
  NAND2_X2 U1750 ( .A1(n2068), .A2(n1196), .ZN(n1433) );
  INV_X4 U1751 ( .A(n2048), .ZN(n2054) );
  XNOR2_X2 U1752 ( .A(n2054), .B(n840), .ZN(n1194) );
  NAND2_X2 U1753 ( .A1(n2045), .A2(n1194), .ZN(n1409) );
  NAND2_X2 U1754 ( .A1(n1433), .A2(n1409), .ZN(n1221) );
  INV_X4 U1755 ( .A(n2081), .ZN(n2087) );
  XNOR2_X2 U1756 ( .A(n2087), .B(n840), .ZN(n1197) );
  NAND2_X2 U1757 ( .A1(n2078), .A2(n1197), .ZN(n1230) );
  INV_X4 U1758 ( .A(n1230), .ZN(n1218) );
  INV_X4 U1759 ( .A(n2099), .ZN(n2095) );
  INV_X4 U1760 ( .A(n2098), .ZN(n2104) );
  XNOR2_X2 U1761 ( .A(n2104), .B(n841), .ZN(n1201) );
  NAND2_X2 U1762 ( .A1(n2095), .A2(n1201), .ZN(n1288) );
  NAND2_X2 U1763 ( .A1(n1970), .A2(n1147), .ZN(n1220) );
  NAND2_X2 U1764 ( .A1(n1957), .A2(n1148), .ZN(n1428) );
  NAND2_X2 U1765 ( .A1(n1220), .A2(n1428), .ZN(n1307) );
  INV_X4 U1766 ( .A(n1307), .ZN(n1398) );
  INV_X4 U1767 ( .A(n1992), .ZN(n1998) );
  XNOR2_X2 U1768 ( .A(n1998), .B(n841), .ZN(n1308) );
  NAND2_X2 U1769 ( .A1(n1989), .A2(n1308), .ZN(n1399) );
  NAND2_X2 U1770 ( .A1(n1398), .A2(n1399), .ZN(n1312) );
  INV_X4 U1771 ( .A(n1312), .ZN(n1405) );
  INV_X4 U1772 ( .A(n2031), .ZN(n2037) );
  XNOR2_X2 U1773 ( .A(n2037), .B(n840), .ZN(n1186) );
  NAND2_X2 U1774 ( .A1(n2028), .A2(n1186), .ZN(n1407) );
  INV_X4 U1775 ( .A(n2011), .ZN(n2017) );
  XNOR2_X2 U1776 ( .A(n2017), .B(n841), .ZN(n1191) );
  NAND2_X2 U1777 ( .A1(n2008), .A2(n1191), .ZN(n1400) );
  INV_X4 U1778 ( .A(n1292), .ZN(n1181) );
  XNOR2_X2 U1779 ( .A(n1150), .B(n1677), .ZN(n1343) );
  XNOR2_X2 U1780 ( .A(n924), .B(n841), .ZN(n1159) );
  NAND2_X2 U1781 ( .A1(n1603), .A2(n1159), .ZN(n1356) );
  INV_X4 U1782 ( .A(n818), .ZN(n1557) );
  XNOR2_X2 U1783 ( .A(n1557), .B(n1154), .ZN(n1151) );
  INV_X4 U1784 ( .A(n1364), .ZN(n1350) );
  XNOR2_X2 U1785 ( .A(n1580), .B(n1154), .ZN(n1152) );
  XNOR2_X2 U1786 ( .A(n1152), .B(n1579), .ZN(n1362) );
  INV_X4 U1787 ( .A(n1362), .ZN(n1353) );
  NAND2_X2 U1788 ( .A1(n1350), .A2(n1353), .ZN(n1157) );
  NAND2_X2 U1789 ( .A1(n1571), .A2(n1153), .ZN(n1366) );
  XNOR2_X2 U1790 ( .A(n1155), .B(n818), .ZN(n1378) );
  INV_X4 U1791 ( .A(n1378), .ZN(n1351) );
  NAND3_X2 U1792 ( .A1(n1157), .A2(n1366), .A3(n1156), .ZN(n1176) );
  XNOR2_X2 U1793 ( .A(n1526), .B(n840), .ZN(n1158) );
  NAND2_X2 U1794 ( .A1(n1513), .A2(n1158), .ZN(n1365) );
  NAND3_X2 U1795 ( .A1(n1364), .A2(n1366), .A3(n1365), .ZN(n1160) );
  XNOR2_X2 U1796 ( .A(n1159), .B(n1613), .ZN(n1370) );
  INV_X4 U1797 ( .A(n1642), .ZN(n1648) );
  XNOR2_X2 U1798 ( .A(n1648), .B(n841), .ZN(n1161) );
  AOI21_X4 U1799 ( .B1(n1356), .B2(n1357), .A(n826), .ZN(n1163) );
  NAND2_X2 U1800 ( .A1(n1632), .A2(n1161), .ZN(n1236) );
  INV_X4 U1801 ( .A(n1236), .ZN(n1162) );
  XNOR2_X2 U1802 ( .A(n1591), .B(n841), .ZN(n1164) );
  NAND2_X2 U1803 ( .A1(n1165), .A2(n1164), .ZN(n1384) );
  INV_X4 U1804 ( .A(n1166), .ZN(n1167) );
  NOR2_X4 U1805 ( .A1(n1382), .A2(n1167), .ZN(n1168) );
  NAND4_X2 U1806 ( .A1(n1170), .A2(n1169), .A3(n1384), .A4(n1168), .ZN(n1172)
         );
  INV_X4 U1807 ( .A(n1359), .ZN(n1235) );
  XNOR2_X2 U1808 ( .A(n1521), .B(n835), .ZN(n1173) );
  INV_X4 U1809 ( .A(n1175), .ZN(n1354) );
  NAND2_X2 U1810 ( .A1(n1370), .A2(n1176), .ZN(n1177) );
  INV_X4 U1811 ( .A(n1177), .ZN(n1355) );
  NAND4_X2 U1812 ( .A1(n1235), .A2(n1354), .A3(n1355), .A4(n1360), .ZN(n1178)
         );
  NAND4_X2 U1813 ( .A1(n1297), .A2(n1204), .A3(n1181), .A4(n1217), .ZN(n1208)
         );
  XNOR2_X2 U1814 ( .A(n1183), .B(n1182), .ZN(n1300) );
  INV_X4 U1815 ( .A(n1300), .ZN(n1206) );
  XNOR2_X2 U1816 ( .A(n1185), .B(n1184), .ZN(n1294) );
  XNOR2_X2 U1817 ( .A(n1186), .B(n2032), .ZN(n1404) );
  XNOR2_X2 U1818 ( .A(n841), .B(n1993), .ZN(n1187) );
  XNOR2_X2 U1819 ( .A(n1998), .B(n1187), .ZN(n1190) );
  XNOR2_X2 U1820 ( .A(n1979), .B(n1970), .ZN(n1188) );
  INV_X4 U1821 ( .A(n1399), .ZN(n1189) );
  AOI21_X4 U1822 ( .B1(n1190), .B2(n1311), .A(n1189), .ZN(n1192) );
  OAI21_X4 U1823 ( .B1(n1192), .B2(n791), .A(n1400), .ZN(n1401) );
  XNOR2_X2 U1824 ( .A(n1194), .B(n2049), .ZN(n1444) );
  INV_X4 U1825 ( .A(n1444), .ZN(n1410) );
  NAND2_X2 U1826 ( .A1(n1410), .A2(n1409), .ZN(n1228) );
  XNOR2_X2 U1827 ( .A(n1196), .B(n1195), .ZN(n1434) );
  NAND2_X2 U1828 ( .A1(n1228), .A2(n1434), .ZN(n1198) );
  AOI21_X4 U1829 ( .B1(n1200), .B2(n1199), .A(n1218), .ZN(n1203) );
  XNOR2_X2 U1830 ( .A(n1201), .B(n2099), .ZN(n1233) );
  INV_X4 U1831 ( .A(n1233), .ZN(n1202) );
  OAI21_X4 U1832 ( .B1(n1203), .B2(n1202), .A(n1288), .ZN(n1295) );
  NAND3_X4 U1833 ( .A1(n1300), .A2(n1294), .A3(n1295), .ZN(n1205) );
  XNOR2_X2 U1834 ( .A(n1210), .B(n1209), .ZN(n2155) );
  INV_X4 U1835 ( .A(n1211), .ZN(n2165) );
  NAND2_X2 U1836 ( .A1(n1211), .A2(n2161), .ZN(n1305) );
  INV_X4 U1837 ( .A(n1305), .ZN(n1459) );
  NOR2_X4 U1838 ( .A1(n1457), .A2(n1459), .ZN(n1213) );
  INV_X4 U1839 ( .A(setInv), .ZN(n1212) );
  XNOR2_X2 U1840 ( .A(n1213), .B(n1212), .ZN(n1214) );
  MUX2_X2 U1841 ( .A(n1215), .B(n1214), .S(aluCtrl[2]), .Z(n1512) );
  INV_X4 U1842 ( .A(n1428), .ZN(n1219) );
  NAND2_X2 U1843 ( .A1(n1399), .A2(n1220), .ZN(n1429) );
  INV_X4 U1844 ( .A(n1429), .ZN(n1223) );
  INV_X4 U1845 ( .A(n1221), .ZN(n1222) );
  NAND4_X2 U1846 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n803), .ZN(n1287)
         );
  INV_X4 U1847 ( .A(n1434), .ZN(n1225) );
  INV_X4 U1848 ( .A(n1433), .ZN(n1227) );
  XNOR2_X2 U1849 ( .A(n1234), .B(n1233), .ZN(n2106) );
  NAND2_X2 U1850 ( .A1(n1236), .A2(n826), .ZN(n1237) );
  NAND3_X2 U1851 ( .A1(n1355), .A2(n1237), .A3(n1343), .ZN(n1246) );
  INV_X4 U1852 ( .A(n1357), .ZN(n1242) );
  NAND2_X2 U1853 ( .A1(n1236), .A2(n1356), .ZN(n1241) );
  INV_X4 U1854 ( .A(n1237), .ZN(n1239) );
  INV_X4 U1855 ( .A(n1343), .ZN(n1238) );
  INV_X4 U1856 ( .A(n1342), .ZN(n1249) );
  INV_X4 U1857 ( .A(n1341), .ZN(n1248) );
  OAI21_X4 U1858 ( .B1(n1249), .B2(n1248), .A(n1247), .ZN(n1419) );
  INV_X4 U1859 ( .A(n1252), .ZN(n1256) );
  NAND2_X2 U1860 ( .A1(n1254), .A2(n1253), .ZN(n1281) );
  INV_X4 U1861 ( .A(n1281), .ZN(n1257) );
  NAND2_X2 U1862 ( .A1(n1316), .A2(n1326), .ZN(n1255) );
  NAND2_X2 U1863 ( .A1(n1256), .A2(n1255), .ZN(n1278) );
  INV_X4 U1864 ( .A(n1277), .ZN(n1258) );
  OAI21_X4 U1865 ( .B1(n1276), .B2(n1258), .A(n1264), .ZN(n1259) );
  INV_X4 U1866 ( .A(n1316), .ZN(n1261) );
  NAND4_X2 U1867 ( .A1(n1271), .A2(n1263), .A3(n1326), .A4(n1262), .ZN(n1274)
         );
  INV_X4 U1868 ( .A(n1282), .ZN(n1268) );
  INV_X4 U1869 ( .A(n1264), .ZN(n1280) );
  INV_X4 U1870 ( .A(n1283), .ZN(n1267) );
  NAND2_X2 U1871 ( .A1(n1269), .A2(n1270), .ZN(n1273) );
  NAND3_X2 U1872 ( .A1(n1274), .A2(n1273), .A3(n1272), .ZN(n1275) );
  XNOR2_X2 U1873 ( .A(n1275), .B(n1319), .ZN(n1912) );
  INV_X4 U1874 ( .A(n1278), .ZN(n1279) );
  XNOR2_X2 U1875 ( .A(n1286), .B(n1285), .ZN(n1893) );
  INV_X4 U1876 ( .A(n1287), .ZN(n1289) );
  NAND2_X2 U1877 ( .A1(n1289), .A2(n1288), .ZN(n1290) );
  XNOR2_X2 U1878 ( .A(n1291), .B(n1294), .ZN(n2127) );
  INV_X4 U1879 ( .A(n1297), .ZN(n1293) );
  XNOR2_X2 U1880 ( .A(n1301), .B(n1206), .ZN(n2149) );
  NAND3_X4 U1881 ( .A1(n1304), .A2(n1303), .A3(n1302), .ZN(n1464) );
  INV_X4 U1882 ( .A(n1464), .ZN(n1452) );
  NAND2_X2 U1883 ( .A1(setInv), .A2(n1305), .ZN(n1306) );
  XNOR2_X2 U1884 ( .A(n1308), .B(n1993), .ZN(n1310) );
  XNOR2_X2 U1885 ( .A(n1309), .B(n1310), .ZN(n2003) );
  INV_X4 U1886 ( .A(n2003), .ZN(n1397) );
  AOI21_X4 U1887 ( .B1(n1399), .B2(n1314), .A(n1313), .ZN(n1315) );
  XNOR2_X2 U1888 ( .A(n1315), .B(n791), .ZN(n2023) );
  INV_X4 U1889 ( .A(n2023), .ZN(n1396) );
  OAI21_X4 U1890 ( .B1(n1318), .B2(n1317), .A(n1316), .ZN(n1416) );
  INV_X4 U1891 ( .A(n1416), .ZN(n1327) );
  OAI211_X2 U1892 ( .C1(n1327), .C2(n1323), .A(n1322), .B(n1321), .ZN(n1324)
         );
  XNOR2_X2 U1893 ( .A(n1324), .B(n824), .ZN(n1325) );
  INV_X4 U1894 ( .A(n1325), .ZN(n1930) );
  XNOR2_X2 U1895 ( .A(n816), .B(n1332), .ZN(n1984) );
  INV_X4 U1896 ( .A(n1333), .ZN(n1334) );
  INV_X4 U1897 ( .A(n1381), .ZN(n1347) );
  NAND2_X2 U1898 ( .A1(n1363), .A2(n1365), .ZN(n1379) );
  AOI21_X2 U1899 ( .B1(n1379), .B2(n1351), .A(n1350), .ZN(n1352) );
  XNOR2_X2 U1900 ( .A(n1353), .B(n1352), .ZN(n1585) );
  NAND2_X2 U1901 ( .A1(n1355), .A2(n1354), .ZN(n1358) );
  INV_X4 U1902 ( .A(n1366), .ZN(n1367) );
  XNOR2_X2 U1903 ( .A(n1371), .B(n1370), .ZN(n1618) );
  INV_X4 U1904 ( .A(n1372), .ZN(n1373) );
  NAND3_X2 U1905 ( .A1(n1375), .A2(n1374), .A3(n1373), .ZN(n1389) );
  XNOR2_X2 U1906 ( .A(n1377), .B(n835), .ZN(n1492) );
  XNOR2_X2 U1907 ( .A(n1379), .B(n1378), .ZN(n1558) );
  INV_X4 U1908 ( .A(n1380), .ZN(n1383) );
  NOR4_X2 U1909 ( .A1(n1389), .A2(n1492), .A3(n1558), .A4(n792), .ZN(n1390) );
  NAND4_X2 U1910 ( .A1(n1392), .A2(n1684), .A3(n1391), .A4(n1390), .ZN(n1393)
         );
  XNOR2_X2 U1911 ( .A(n1404), .B(n1403), .ZN(n2040) );
  INV_X4 U1912 ( .A(n2040), .ZN(n1449) );
  NAND2_X2 U1913 ( .A1(n803), .A2(n1409), .ZN(n1430) );
  INV_X4 U1914 ( .A(n1430), .ZN(n1406) );
  NAND2_X2 U1915 ( .A1(n1406), .A2(n1405), .ZN(n1412) );
  INV_X4 U1916 ( .A(n1441), .ZN(n1411) );
  XNOR2_X2 U1917 ( .A(n1414), .B(n1434), .ZN(n2062) );
  INV_X4 U1918 ( .A(n2062), .ZN(n1448) );
  INV_X4 U1919 ( .A(n1417), .ZN(n1427) );
  NAND2_X2 U1920 ( .A1(n1422), .A2(n1421), .ZN(n1425) );
  XNOR2_X2 U1921 ( .A(n1427), .B(n1426), .ZN(n1935) );
  NAND2_X2 U1922 ( .A1(n1789), .A2(n1935), .ZN(n1446) );
  NAND2_X2 U1923 ( .A1(n1433), .A2(n1428), .ZN(n1431) );
  NOR4_X2 U1924 ( .A1(n1432), .A2(n1431), .A3(n1430), .A4(n1429), .ZN(n1438)
         );
  XNOR2_X2 U1925 ( .A(n1439), .B(n787), .ZN(n2090) );
  XNOR2_X2 U1926 ( .A(n1445), .B(n1444), .ZN(n2057) );
  NAND3_X2 U1927 ( .A1(n1449), .A2(n1448), .A3(n1447), .ZN(n1454) );
  OAI211_X2 U1928 ( .C1(n1452), .C2(n1460), .A(n1451), .B(n1450), .ZN(n1469)
         );
  INV_X4 U1929 ( .A(n1454), .ZN(n1455) );
  NAND3_X2 U1930 ( .A1(n1469), .A2(n1468), .A3(n1467), .ZN(n1511) );
  AOI22_X2 U1931 ( .A1(n1688), .A2(n993), .B1(n1472), .B2(n1471), .ZN(n1477)
         );
  NAND2_X2 U1932 ( .A1(n1473), .A2(n1591), .ZN(n1476) );
  INV_X4 U1933 ( .A(n833), .ZN(n1484) );
  NAND2_X2 U1934 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  INV_X4 U1935 ( .A(n1480), .ZN(n1483) );
  MUX2_X2 U1936 ( .A(n1487), .B(n1486), .S(n1503), .Z(n1488) );
  INV_X4 U1937 ( .A(n1488), .ZN(n2174) );
  INV_X4 U1938 ( .A(n2174), .ZN(n1490) );
  INV_X4 U1939 ( .A(n1492), .ZN(n1494) );
  NAND2_X2 U1940 ( .A1(n1500), .A2(n1499), .ZN(n1502) );
  NAND2_X2 U1941 ( .A1(busA[0]), .A2(fp), .ZN(n1505) );
  INV_X4 U1942 ( .A(n1505), .ZN(n1501) );
  AOI221_X2 U1943 ( .B1(n1504), .B2(n1503), .C1(n2133), .C2(n1502), .A(n1501), 
        .ZN(n1506) );
  AOI21_X4 U1944 ( .B1(n1509), .B2(n853), .A(n1508), .ZN(n1510) );
  OAI211_X2 U1945 ( .C1(n1512), .C2(n813), .A(n1511), .B(n1510), .ZN(aluRes[0]) );
  NAND2_X2 U1946 ( .A1(n2130), .A2(n853), .ZN(n2163) );
  MUX2_X2 U1947 ( .A(n851), .B(n2163), .S(n1513), .Z(n1514) );
  NAND2_X2 U1948 ( .A1(n2133), .A2(n853), .ZN(n2158) );
  NAND2_X2 U1949 ( .A1(n1514), .A2(n847), .ZN(n1525) );
  NAND2_X2 U1950 ( .A1(n2143), .A2(n853), .ZN(n2113) );
  NAND2_X2 U1951 ( .A1(n1638), .A2(n1864), .ZN(n1518) );
  INV_X4 U1952 ( .A(n1515), .ZN(n1706) );
  NAND2_X2 U1953 ( .A1(n1706), .A2(n1868), .ZN(n1517) );
  INV_X4 U1954 ( .A(n2089), .ZN(n1519) );
  NAND2_X2 U1955 ( .A1(n1527), .A2(n853), .ZN(n2151) );
  NAND2_X2 U1956 ( .A1(n845), .A2(n2107), .ZN(n1542) );
  NAND2_X2 U1957 ( .A1(n1528), .A2(n853), .ZN(n1788) );
  AOI22_X2 U1958 ( .A1(fp), .A2(busA[4]), .B1(n852), .B2(n792), .ZN(n1541) );
  INV_X4 U1959 ( .A(n1529), .ZN(n1530) );
  INV_X4 U1960 ( .A(n833), .ZN(n1532) );
  NAND2_X2 U1961 ( .A1(n1532), .A2(n1531), .ZN(n1539) );
  NAND2_X2 U1962 ( .A1(n1587), .A2(n1586), .ZN(n1538) );
  NAND2_X2 U1963 ( .A1(n1862), .A2(n1650), .ZN(n1537) );
  NAND2_X2 U1964 ( .A1(n799), .A2(n1769), .ZN(n1534) );
  NAND2_X2 U1965 ( .A1(n1866), .A2(n1649), .ZN(n1536) );
  NAND4_X2 U1966 ( .A1(n1539), .A2(n1538), .A3(n1537), .A4(n1536), .ZN(n2064)
         );
  AOI22_X2 U1967 ( .A1(n2108), .A2(n2064), .B1(n2124), .B2(n2088), .ZN(n1540)
         );
  NAND4_X2 U1968 ( .A1(n1543), .A2(n1542), .A3(n1541), .A4(n1540), .ZN(
        aluRes[4]) );
  MUX2_X2 U1969 ( .A(n851), .B(n2163), .S(n1544), .Z(n1545) );
  NAND2_X2 U1970 ( .A1(n1545), .A2(n847), .ZN(n1556) );
  NAND2_X2 U1971 ( .A1(n1672), .A2(n1864), .ZN(n1549) );
  INV_X4 U1972 ( .A(n1546), .ZN(n1739) );
  NAND2_X2 U1973 ( .A1(n1739), .A2(n1868), .ZN(n1548) );
  INV_X4 U1974 ( .A(n2063), .ZN(n1550) );
  NAND2_X2 U1975 ( .A1(n845), .A2(n2089), .ZN(n1569) );
  AOI22_X2 U1976 ( .A1(fp), .A2(busA[5]), .B1(n852), .B2(n1558), .ZN(n1568) );
  NAND2_X2 U1977 ( .A1(n1862), .A2(n1692), .ZN(n1566) );
  NAND2_X2 U1978 ( .A1(n799), .A2(n1735), .ZN(n1560) );
  NAND2_X2 U1979 ( .A1(n1816), .A2(n1691), .ZN(n1565) );
  NAND2_X2 U1980 ( .A1(n1864), .A2(n1619), .ZN(n1563) );
  NAND4_X2 U1981 ( .A1(n1566), .A2(n1565), .A3(n1564), .A4(n1563), .ZN(n2047)
         );
  AOI22_X2 U1982 ( .A1(n2108), .A2(n2047), .B1(n2124), .B2(n2064), .ZN(n1567)
         );
  NAND4_X2 U1983 ( .A1(n1570), .A2(n1569), .A3(n1568), .A4(n1567), .ZN(
        aluRes[5]) );
  MUX2_X2 U1984 ( .A(n851), .B(n2163), .S(n1571), .Z(n1572) );
  NAND2_X2 U1985 ( .A1(n1572), .A2(n847), .ZN(n1584) );
  NAND2_X2 U1986 ( .A1(n1573), .A2(n1866), .ZN(n1577) );
  NAND2_X2 U1987 ( .A1(n1638), .A2(n1862), .ZN(n1576) );
  NAND2_X2 U1988 ( .A1(n1706), .A2(n1864), .ZN(n1575) );
  INV_X4 U1989 ( .A(n1775), .ZN(n1707) );
  NAND2_X2 U1990 ( .A1(n1707), .A2(n1868), .ZN(n1574) );
  NAND4_X2 U1991 ( .A1(n1577), .A2(n1576), .A3(n1575), .A4(n1574), .ZN(n2056)
         );
  INV_X4 U1992 ( .A(n2056), .ZN(n1578) );
  NAND2_X2 U1993 ( .A1(n845), .A2(n2063), .ZN(n1601) );
  AOI22_X2 U1994 ( .A1(fp), .A2(busA[6]), .B1(n852), .B2(n1585), .ZN(n1600) );
  NAND2_X2 U1995 ( .A1(n1586), .A2(n1484), .ZN(n1598) );
  INV_X4 U1996 ( .A(n783), .ZN(n1587) );
  NAND2_X2 U1997 ( .A1(n1587), .A2(n1650), .ZN(n1597) );
  INV_X4 U1998 ( .A(n1649), .ZN(n1724) );
  INV_X4 U1999 ( .A(n1588), .ZN(n1592) );
  INV_X4 U2000 ( .A(n1655), .ZN(n1589) );
  AOI21_X2 U2001 ( .B1(n799), .B2(n1702), .A(n1589), .ZN(n1590) );
  INV_X4 U2002 ( .A(n1593), .ZN(n1795) );
  AOI22_X2 U2003 ( .A1(n2108), .A2(n2055), .B1(n2124), .B2(n2047), .ZN(n1599)
         );
  NAND4_X2 U2004 ( .A1(n1602), .A2(n1601), .A3(n1600), .A4(n1599), .ZN(
        aluRes[6]) );
  MUX2_X2 U2005 ( .A(n851), .B(n2163), .S(n1603), .Z(n1604) );
  NAND2_X2 U2006 ( .A1(n1604), .A2(n847), .ZN(n1617) );
  NAND2_X2 U2007 ( .A1(n1605), .A2(n1866), .ZN(n1611) );
  NAND2_X2 U2008 ( .A1(n1672), .A2(n1862), .ZN(n1610) );
  NAND2_X2 U2009 ( .A1(n1739), .A2(n1864), .ZN(n1609) );
  INV_X4 U2010 ( .A(n1802), .ZN(n1740) );
  NAND2_X2 U2011 ( .A1(n1740), .A2(n1868), .ZN(n1608) );
  NAND4_X2 U2012 ( .A1(n1611), .A2(n1610), .A3(n1609), .A4(n1608), .ZN(n2039)
         );
  INV_X4 U2013 ( .A(n2039), .ZN(n2020) );
  NAND2_X2 U2014 ( .A1(n845), .A2(n2056), .ZN(n1630) );
  AOI22_X2 U2015 ( .A1(fp), .A2(busA[7]), .B1(n852), .B2(n1618), .ZN(n1629) );
  NAND2_X2 U2016 ( .A1(n1484), .A2(n1619), .ZN(n1627) );
  NAND2_X2 U2017 ( .A1(n1692), .A2(n1587), .ZN(n1626) );
  NAND2_X2 U2018 ( .A1(n799), .A2(n1668), .ZN(n1621) );
  INV_X4 U2019 ( .A(n1817), .ZN(n1761) );
  INV_X4 U2020 ( .A(n1691), .ZN(n1762) );
  AOI22_X2 U2021 ( .A1(n2108), .A2(n2038), .B1(n2124), .B2(n2055), .ZN(n1628)
         );
  NAND4_X2 U2022 ( .A1(n1631), .A2(n1630), .A3(n1629), .A4(n1628), .ZN(
        aluRes[7]) );
  MUX2_X2 U2023 ( .A(n851), .B(n2163), .S(n1632), .Z(n1633) );
  NAND2_X2 U2024 ( .A1(n1633), .A2(n847), .ZN(n1647) );
  NAND2_X2 U2025 ( .A1(n1707), .A2(n1864), .ZN(n1641) );
  AOI21_X2 U2026 ( .B1(n1770), .B2(n1653), .A(n1634), .ZN(n1637) );
  NAND2_X2 U2027 ( .A1(n799), .A2(n1635), .ZN(n1636) );
  NAND2_X2 U2028 ( .A1(n1637), .A2(n1636), .ZN(n1831) );
  NAND2_X2 U2029 ( .A1(n1868), .A2(n1831), .ZN(n1640) );
  AOI22_X2 U2030 ( .A1(n1706), .A2(n1862), .B1(n1638), .B2(n1866), .ZN(n1639)
         );
  INV_X4 U2031 ( .A(n1683), .ZN(n2019) );
  NAND2_X2 U2032 ( .A1(n845), .A2(n2039), .ZN(n1664) );
  AOI22_X2 U2033 ( .A1(fp), .A2(busA[8]), .B1(n852), .B2(n793), .ZN(n1663) );
  NAND2_X2 U2034 ( .A1(n1587), .A2(n1649), .ZN(n1661) );
  NAND2_X2 U2035 ( .A1(n1650), .A2(n1532), .ZN(n1660) );
  NAND2_X2 U2036 ( .A1(n799), .A2(n1653), .ZN(n1654) );
  INV_X4 U2037 ( .A(n1850), .ZN(n1794) );
  AOI22_X2 U2038 ( .A1(n2108), .A2(n2018), .B1(n2124), .B2(n2038), .ZN(n1662)
         );
  NAND4_X2 U2039 ( .A1(n1665), .A2(n1664), .A3(n1663), .A4(n1662), .ZN(
        aluRes[8]) );
  MUX2_X2 U2040 ( .A(n851), .B(n2163), .S(n1666), .Z(n1667) );
  NAND2_X2 U2041 ( .A1(n1667), .A2(n847), .ZN(n1681) );
  NAND2_X2 U2042 ( .A1(n1770), .A2(n1668), .ZN(n1671) );
  INV_X4 U2043 ( .A(n1865), .ZN(n1675) );
  NAND2_X2 U2044 ( .A1(n1740), .A2(n1864), .ZN(n1674) );
  AOI22_X2 U2045 ( .A1(n1739), .A2(n1862), .B1(n1672), .B2(n1866), .ZN(n1673)
         );
  OAI211_X2 U2046 ( .C1(n1675), .C2(n833), .A(n1674), .B(n1673), .ZN(n1718) );
  INV_X4 U2047 ( .A(n1718), .ZN(n2000) );
  NAND2_X2 U2048 ( .A1(n845), .A2(n1683), .ZN(n1698) );
  NAND2_X2 U2049 ( .A1(n799), .A2(n1687), .ZN(n1690) );
  NAND2_X2 U2050 ( .A1(n1770), .A2(n1688), .ZN(n1689) );
  AOI22_X2 U2051 ( .A1(n1723), .A2(n1867), .B1(n1862), .B2(n1817), .ZN(n1695)
         );
  NAND2_X2 U2052 ( .A1(n1864), .A2(n1691), .ZN(n1694) );
  NAND2_X2 U2053 ( .A1(n1868), .A2(n1692), .ZN(n1693) );
  AOI22_X2 U2054 ( .A1(n2108), .A2(n1999), .B1(n2124), .B2(n2018), .ZN(n1696)
         );
  NAND4_X2 U2055 ( .A1(n1699), .A2(n1698), .A3(n1697), .A4(n1696), .ZN(
        aluRes[9]) );
  MUX2_X2 U2056 ( .A(n851), .B(n2163), .S(n1700), .Z(n1701) );
  NAND2_X2 U2057 ( .A1(n1701), .A2(n847), .ZN(n1716) );
  NAND2_X2 U2058 ( .A1(n1864), .A2(n1831), .ZN(n1710) );
  NAND2_X2 U2059 ( .A1(n1770), .A2(n1702), .ZN(n1705) );
  NAND2_X2 U2060 ( .A1(n799), .A2(n1703), .ZN(n1704) );
  NAND2_X2 U2061 ( .A1(n1868), .A2(n1847), .ZN(n1709) );
  AOI22_X2 U2062 ( .A1(n1707), .A2(n1862), .B1(n1706), .B2(n1866), .ZN(n1708)
         );
  NAND3_X2 U2063 ( .A1(n1710), .A2(n1709), .A3(n1708), .ZN(n1751) );
  INV_X4 U2064 ( .A(n1751), .ZN(n1981) );
  NAND2_X2 U2065 ( .A1(n845), .A2(n1718), .ZN(n1731) );
  AOI22_X2 U2066 ( .A1(fp), .A2(busA[10]), .B1(n852), .B2(n788), .ZN(n1730) );
  INV_X4 U2067 ( .A(n798), .ZN(n1723) );
  NAND2_X2 U2068 ( .A1(n1770), .A2(n1719), .ZN(n1722) );
  NAND2_X2 U2069 ( .A1(n799), .A2(n1720), .ZN(n1721) );
  AOI22_X2 U2070 ( .A1(n1723), .A2(n1851), .B1(n1862), .B2(n1850), .ZN(n1728)
         );
  NAND2_X2 U2071 ( .A1(n1728), .A2(n1727), .ZN(n1980) );
  AOI22_X2 U2072 ( .A1(n2108), .A2(n1980), .B1(n2124), .B2(n1999), .ZN(n1729)
         );
  NAND4_X2 U2073 ( .A1(n1732), .A2(n1731), .A3(n1730), .A4(n1729), .ZN(
        aluRes[10]) );
  MUX2_X2 U2074 ( .A(n851), .B(n2163), .S(n1733), .Z(n1734) );
  NAND2_X2 U2075 ( .A1(n1734), .A2(n847), .ZN(n1749) );
  NAND2_X2 U2076 ( .A1(n1864), .A2(n1865), .ZN(n1743) );
  NAND2_X2 U2077 ( .A1(n1770), .A2(n1735), .ZN(n1738) );
  NAND2_X2 U2078 ( .A1(n799), .A2(n1736), .ZN(n1737) );
  NAND2_X2 U2079 ( .A1(n1868), .A2(n1861), .ZN(n1742) );
  AOI22_X2 U2080 ( .A1(n1740), .A2(n1862), .B1(n1739), .B2(n1866), .ZN(n1741)
         );
  NAND3_X2 U2081 ( .A1(n1743), .A2(n1742), .A3(n1741), .ZN(n1787) );
  INV_X4 U2082 ( .A(n1787), .ZN(n1966) );
  NAND2_X2 U2083 ( .A1(n845), .A2(n1751), .ZN(n1765) );
  AOI22_X2 U2084 ( .A1(fp), .A2(busA[11]), .B1(n852), .B2(n795), .ZN(n1764) );
  NAND2_X2 U2085 ( .A1(n1770), .A2(n1752), .ZN(n1755) );
  NAND2_X2 U2086 ( .A1(n799), .A2(n1753), .ZN(n1754) );
  INV_X4 U2087 ( .A(n1863), .ZN(n1756) );
  INV_X4 U2088 ( .A(n1867), .ZN(n1757) );
  OAI221_X2 U2089 ( .B1(n1762), .B2(n833), .C1(n1761), .C2(n783), .A(n1760), 
        .ZN(n1946) );
  AOI22_X2 U2090 ( .A1(n2108), .A2(n1946), .B1(n2124), .B2(n1980), .ZN(n1763)
         );
  NAND4_X2 U2091 ( .A1(n1766), .A2(n1765), .A3(n1764), .A4(n1763), .ZN(
        aluRes[11]) );
  MUX2_X2 U2092 ( .A(n851), .B(n2163), .S(n1767), .Z(n1768) );
  NAND2_X2 U2093 ( .A1(n1768), .A2(n847), .ZN(n1785) );
  NAND2_X2 U2094 ( .A1(n1864), .A2(n1847), .ZN(n1779) );
  NAND2_X2 U2095 ( .A1(n1770), .A2(n1769), .ZN(n1774) );
  NAND2_X2 U2096 ( .A1(n1868), .A2(n1848), .ZN(n1778) );
  INV_X4 U2097 ( .A(n1814), .ZN(n1937) );
  NAND2_X2 U2098 ( .A1(n845), .A2(n1787), .ZN(n1798) );
  INV_X4 U2099 ( .A(n1848), .ZN(n1833) );
  INV_X4 U2100 ( .A(n1851), .ZN(n1832) );
  OAI221_X2 U2101 ( .B1(n1795), .B2(n833), .C1(n1794), .C2(n783), .A(n1793), 
        .ZN(n1815) );
  AOI22_X2 U2102 ( .A1(n2108), .A2(n1815), .B1(n2124), .B2(n1946), .ZN(n1796)
         );
  NAND4_X2 U2103 ( .A1(n1799), .A2(n1798), .A3(n1797), .A4(n1796), .ZN(
        aluRes[12]) );
  MUX2_X2 U2104 ( .A(n851), .B(n2163), .S(n1800), .Z(n1801) );
  NAND2_X2 U2105 ( .A1(n1801), .A2(n847), .ZN(n1812) );
  NAND2_X2 U2106 ( .A1(n1864), .A2(n1861), .ZN(n1806) );
  NAND2_X2 U2107 ( .A1(n1868), .A2(n1863), .ZN(n1805) );
  INV_X4 U2108 ( .A(n1846), .ZN(n1927) );
  NAND2_X2 U2109 ( .A1(n845), .A2(n1814), .ZN(n1827) );
  INV_X4 U2110 ( .A(n1815), .ZN(n1947) );
  INV_X4 U2111 ( .A(n798), .ZN(n1816) );
  NAND2_X2 U2112 ( .A1(n1861), .A2(n1816), .ZN(n1821) );
  NAND2_X2 U2113 ( .A1(n1862), .A2(n1863), .ZN(n1820) );
  NAND2_X2 U2114 ( .A1(n1484), .A2(n1817), .ZN(n1819) );
  NAND2_X2 U2115 ( .A1(n1864), .A2(n1867), .ZN(n1818) );
  NAND4_X2 U2116 ( .A1(n1821), .A2(n1820), .A3(n1819), .A4(n1818), .ZN(n1926)
         );
  INV_X4 U2117 ( .A(n1926), .ZN(n1900) );
  NAND4_X2 U2118 ( .A1(n1828), .A2(n1827), .A3(n1826), .A4(n1825), .ZN(
        aluRes[13]) );
  MUX2_X2 U2119 ( .A(n851), .B(n2163), .S(n1829), .Z(n1830) );
  NAND2_X2 U2120 ( .A1(n1830), .A2(n847), .ZN(n1844) );
  NAND2_X2 U2121 ( .A1(n1831), .A2(n1723), .ZN(n1838) );
  NAND2_X2 U2122 ( .A1(n1862), .A2(n1847), .ZN(n1837) );
  INV_X4 U2123 ( .A(n1892), .ZN(n1909) );
  NAND2_X2 U2124 ( .A1(n845), .A2(n1846), .ZN(n1859) );
  NAND2_X2 U2125 ( .A1(n1847), .A2(n1816), .ZN(n1855) );
  NAND2_X2 U2126 ( .A1(n1862), .A2(n1848), .ZN(n1854) );
  NAND2_X2 U2127 ( .A1(n1532), .A2(n1850), .ZN(n1853) );
  NAND2_X2 U2128 ( .A1(n1864), .A2(n1851), .ZN(n1852) );
  NAND4_X2 U2129 ( .A1(n1855), .A2(n1854), .A3(n1853), .A4(n1852), .ZN(n1908)
         );
  AOI22_X2 U2130 ( .A1(n2108), .A2(n1908), .B1(n2124), .B2(n1926), .ZN(n1858)
         );
  AOI22_X2 U2131 ( .A1(busA[14]), .A2(fp), .B1(n852), .B2(n1856), .ZN(n1857)
         );
  NAND4_X2 U2132 ( .A1(n1860), .A2(n1859), .A3(n1858), .A4(n1857), .ZN(
        aluRes[14]) );
  NAND2_X2 U2133 ( .A1(n1862), .A2(n1861), .ZN(n1872) );
  NAND2_X2 U2134 ( .A1(n1864), .A2(n1863), .ZN(n1871) );
  NAND2_X2 U2135 ( .A1(n1866), .A2(n1865), .ZN(n1870) );
  NAND2_X2 U2136 ( .A1(n1868), .A2(n1867), .ZN(n1869) );
  MUX2_X2 U2137 ( .A(n851), .B(n2163), .S(n1875), .Z(n1876) );
  NAND2_X2 U2138 ( .A1(n1876), .A2(n847), .ZN(n1878) );
  NAND2_X2 U2139 ( .A1(busA[15]), .A2(fp), .ZN(n1881) );
  AOI22_X2 U2140 ( .A1(n852), .A2(n800), .B1(n2124), .B2(n1908), .ZN(n1880) );
  NAND4_X2 U2141 ( .A1(n1883), .A2(n1882), .A3(n1881), .A4(n1880), .ZN(
        aluRes[15]) );
  MUX2_X2 U2142 ( .A(n851), .B(n2163), .S(n1886), .Z(n1887) );
  NAND2_X2 U2143 ( .A1(n1887), .A2(n847), .ZN(n1890) );
  INV_X4 U2144 ( .A(n1908), .ZN(n1888) );
  NAND2_X2 U2145 ( .A1(busA[16]), .A2(fp), .ZN(n1895) );
  AOI22_X2 U2146 ( .A1(n852), .A2(n1893), .B1(n2108), .B2(n1892), .ZN(n1894)
         );
  NAND4_X2 U2147 ( .A1(n1897), .A2(n1896), .A3(n1895), .A4(n1894), .ZN(
        aluRes[16]) );
  MUX2_X2 U2148 ( .A(n851), .B(n2163), .S(n1898), .Z(n1899) );
  NAND2_X2 U2149 ( .A1(n1899), .A2(n847), .ZN(n1906) );
  NAND2_X2 U2150 ( .A1(n845), .A2(n1908), .ZN(n1915) );
  AOI22_X2 U2151 ( .A1(busA[17]), .A2(fp), .B1(n852), .B2(n1912), .ZN(n1913)
         );
  NAND4_X2 U2152 ( .A1(n1916), .A2(n1915), .A3(n1914), .A4(n1913), .ZN(
        aluRes[17]) );
  MUX2_X2 U2153 ( .A(n851), .B(n2163), .S(n1917), .Z(n1918) );
  NAND2_X2 U2154 ( .A1(n1918), .A2(n847), .ZN(n1924) );
  NAND2_X2 U2155 ( .A1(n845), .A2(n1926), .ZN(n1933) );
  AOI22_X2 U2156 ( .A1(busA[18]), .A2(fp), .B1(n852), .B2(n1930), .ZN(n1931)
         );
  NAND4_X2 U2157 ( .A1(n1934), .A2(n1933), .A3(n1932), .A4(n1931), .ZN(
        aluRes[18]) );
  NAND2_X2 U2158 ( .A1(busA[19]), .A2(fp), .ZN(n1954) );
  INV_X4 U2159 ( .A(n1935), .ZN(n1936) );
  NAND2_X2 U2160 ( .A1(n852), .A2(n1936), .ZN(n1953) );
  MUX2_X2 U2161 ( .A(n785), .B(n849), .S(n1942), .Z(n1940) );
  NAND2_X2 U2162 ( .A1(n1945), .A2(n1944), .ZN(n1950) );
  INV_X4 U2163 ( .A(n1946), .ZN(n1962) );
  NAND4_X2 U2164 ( .A1(n1954), .A2(n1953), .A3(n1952), .A4(n1951), .ZN(
        aluRes[19]) );
  MUX2_X2 U2165 ( .A(n785), .B(n849), .S(n1957), .Z(n1955) );
  NAND2_X2 U2166 ( .A1(n1960), .A2(n1959), .ZN(n1965) );
  INV_X4 U2167 ( .A(n1980), .ZN(n1961) );
  OAI22_X2 U2168 ( .A1(n1981), .A2(n2157), .B1(n1966), .B2(n2170), .ZN(n1967)
         );
  NAND2_X2 U2169 ( .A1(n1969), .A2(n1968), .ZN(aluRes[20]) );
  MUX2_X2 U2170 ( .A(n851), .B(n2163), .S(n1970), .Z(n1971) );
  NAND2_X2 U2171 ( .A1(n1971), .A2(n847), .ZN(n1978) );
  INV_X4 U2172 ( .A(n1999), .ZN(n1972) );
  NAND2_X2 U2173 ( .A1(n845), .A2(n1980), .ZN(n1987) );
  AOI22_X2 U2174 ( .A1(busA[21]), .A2(fp), .B1(n852), .B2(n1984), .ZN(n1985)
         );
  NAND4_X2 U2175 ( .A1(n1988), .A2(n1987), .A3(n1986), .A4(n1985), .ZN(
        aluRes[21]) );
  MUX2_X2 U2176 ( .A(n851), .B(n2163), .S(n1989), .Z(n1990) );
  NAND2_X2 U2177 ( .A1(n1990), .A2(n847), .ZN(n1997) );
  INV_X4 U2178 ( .A(n2018), .ZN(n1991) );
  NAND2_X2 U2179 ( .A1(n845), .A2(n1999), .ZN(n2006) );
  AOI22_X2 U2180 ( .A1(busA[22]), .A2(fp), .B1(n852), .B2(n2003), .ZN(n2004)
         );
  NAND4_X2 U2181 ( .A1(n2007), .A2(n2006), .A3(n2005), .A4(n2004), .ZN(
        aluRes[22]) );
  MUX2_X2 U2182 ( .A(n851), .B(n2163), .S(n2008), .Z(n2009) );
  NAND2_X2 U2183 ( .A1(n2009), .A2(n847), .ZN(n2016) );
  INV_X4 U2184 ( .A(n2038), .ZN(n2010) );
  NAND2_X2 U2185 ( .A1(n845), .A2(n2018), .ZN(n2026) );
  NAND4_X2 U2186 ( .A1(n2027), .A2(n2026), .A3(n2025), .A4(n2024), .ZN(
        aluRes[23]) );
  MUX2_X2 U2187 ( .A(n851), .B(n2163), .S(n2028), .Z(n2029) );
  NAND2_X2 U2188 ( .A1(n2029), .A2(n847), .ZN(n2036) );
  INV_X4 U2189 ( .A(n2055), .ZN(n2030) );
  NAND2_X2 U2190 ( .A1(n845), .A2(n2038), .ZN(n2043) );
  AOI22_X2 U2191 ( .A1(n2108), .A2(n2056), .B1(n2124), .B2(n2039), .ZN(n2042)
         );
  AOI22_X2 U2192 ( .A1(busA[24]), .A2(fp), .B1(n852), .B2(n2040), .ZN(n2041)
         );
  NAND4_X2 U2193 ( .A1(n2044), .A2(n2043), .A3(n2042), .A4(n2041), .ZN(
        aluRes[24]) );
  MUX2_X2 U2194 ( .A(n851), .B(n2163), .S(n2045), .Z(n2046) );
  NAND2_X2 U2195 ( .A1(n2046), .A2(n847), .ZN(n2053) );
  INV_X4 U2196 ( .A(n2047), .ZN(n2065) );
  NAND2_X2 U2197 ( .A1(n845), .A2(n2055), .ZN(n2060) );
  AOI22_X2 U2198 ( .A1(n2108), .A2(n2063), .B1(n2124), .B2(n2056), .ZN(n2059)
         );
  AOI22_X2 U2199 ( .A1(busA[25]), .A2(fp), .B1(n852), .B2(n2057), .ZN(n2058)
         );
  NAND4_X2 U2200 ( .A1(n2061), .A2(n2060), .A3(n2059), .A4(n2058), .ZN(
        aluRes[25]) );
  NAND2_X2 U2201 ( .A1(busA[26]), .A2(fp), .ZN(n2077) );
  NAND2_X2 U2202 ( .A1(n852), .A2(n2062), .ZN(n2076) );
  AOI22_X2 U2203 ( .A1(n2124), .A2(n2063), .B1(n2108), .B2(n2089), .ZN(n2075)
         );
  INV_X4 U2204 ( .A(n2064), .ZN(n2080) );
  OAI22_X2 U2205 ( .A1(n2065), .A2(n2151), .B1(n2080), .B2(n843), .ZN(n2073)
         );
  MUX2_X2 U2206 ( .A(n785), .B(n849), .S(n2068), .Z(n2066) );
  NAND2_X2 U2207 ( .A1(n2071), .A2(n2070), .ZN(n2072) );
  NAND4_X2 U2208 ( .A1(n2077), .A2(n2076), .A3(n2075), .A4(n2074), .ZN(
        aluRes[26]) );
  MUX2_X2 U2209 ( .A(n851), .B(n2163), .S(n2078), .Z(n2079) );
  NAND2_X2 U2210 ( .A1(n2079), .A2(n847), .ZN(n2086) );
  NAND2_X2 U2211 ( .A1(n844), .A2(n2088), .ZN(n2093) );
  AOI22_X2 U2212 ( .A1(n2108), .A2(n2107), .B1(n2124), .B2(n2089), .ZN(n2092)
         );
  NAND4_X2 U2213 ( .A1(n2094), .A2(n2093), .A3(n2092), .A4(n2091), .ZN(
        aluRes[27]) );
  MUX2_X2 U2214 ( .A(n851), .B(n2163), .S(n2095), .Z(n2096) );
  NAND2_X2 U2215 ( .A1(n2096), .A2(n847), .ZN(n2103) );
  NAND2_X2 U2216 ( .A1(n844), .A2(n2105), .ZN(n2111) );
  AOI22_X2 U2217 ( .A1(busA[28]), .A2(fp), .B1(n852), .B2(n2106), .ZN(n2110)
         );
  AOI22_X2 U2218 ( .A1(n2108), .A2(n2123), .B1(n2124), .B2(n2107), .ZN(n2109)
         );
  NAND4_X2 U2219 ( .A1(n2112), .A2(n2111), .A3(n2110), .A4(n2109), .ZN(
        aluRes[28]) );
  OAI22_X2 U2220 ( .A1(n2114), .A2(n2151), .B1(n2152), .B2(n2113), .ZN(n2122)
         );
  MUX2_X2 U2221 ( .A(n785), .B(n849), .S(n2117), .Z(n2115) );
  NAND2_X2 U2222 ( .A1(n2120), .A2(n2119), .ZN(n2121) );
  NAND2_X2 U2223 ( .A1(n2124), .A2(n2123), .ZN(n2125) );
  AOI211_X2 U2224 ( .C1(n852), .C2(n2127), .A(n2126), .B(n814), .ZN(n2128) );
  NAND2_X2 U2225 ( .A1(n2129), .A2(n2128), .ZN(aluRes[29]) );
  MUX2_X2 U2226 ( .A(n2131), .B(n2130), .S(n2138), .Z(n2132) );
  NAND2_X2 U2227 ( .A1(n2138), .A2(n2137), .ZN(n2146) );
  INV_X4 U2228 ( .A(n2139), .ZN(n2141) );
  NAND2_X2 U2229 ( .A1(n2141), .A2(n1023), .ZN(n2145) );
  NAND4_X2 U2230 ( .A1(n2147), .A2(n2146), .A3(n2145), .A4(n2144), .ZN(n2148)
         );
  MUX2_X2 U2231 ( .A(n2148), .B(busA[30]), .S(fp), .Z(n2154) );
  OAI221_X2 U2232 ( .B1(n2152), .B2(n2151), .C1(n2171), .C2(n2157), .A(n2150), 
        .ZN(n2153) );
  INV_X4 U2233 ( .A(n2161), .ZN(n2159) );
  OAI22_X2 U2234 ( .A1(n2165), .A2(n851), .B1(n2164), .B2(n2163), .ZN(n2166)
         );
  NAND2_X2 U2235 ( .A1(n804), .A2(n2174), .ZN(n2176) );
  INV_X4 U2236 ( .A(busA[31]), .ZN(n2175) );
  MUX2_X2 U2237 ( .A(n2176), .B(n2175), .S(fp), .Z(n2177) );
  NAND2_X2 U2238 ( .A1(n2178), .A2(n2177), .ZN(aluRes[31]) );
endmodule

