
module pipeline ( clk, rst, initPC, instruction, iAddr, memAddr, memRdData, 
        memWrData, dSize, memWr, busA, busB, busFP, rs1, rs2, rd, regWrData, 
        regWr, fp );
  input [31:0] initPC;
  input [31:0] instruction;
  output [31:0] iAddr;
  output [31:0] memAddr;
  input [31:0] memRdData;
  output [31:0] memWrData;
  output [1:0] dSize;
  input [31:0] busA;
  input [31:0] busB;
  input [31:0] busFP;
  output [4:0] rs1;
  output [4:0] rs2;
  output [4:0] rd;
  output [31:0] regWrData;
  input clk, rst;
  output memWr, regWr, fp;
  wire   not_trap_3, op0_1, valid_2, valid_3, setInv_2, op0_2, zeroExt_2,
         link_3, op0_3, fp_3, \id_ex/N44 , \id_ex/N42 , \id_ex/N41 ,
         \id_ex/N40 , \id_ex/N39 , \id_ex/N38 , \id_ex/N37 , \id_ex/N36 ,
         \id_ex/N33 , \id_ex/N31 , \id_ex/N30 , \id_ex/N4 , \ex_mem/N247 ,
         \ex_mem/N246 , \ex_mem/N245 , \ex_mem/N244 , \ex_mem/N243 ,
         \ex_mem/N242 , \ex_mem/N241 , \ex_mem/N240 , \ex_mem/N239 ,
         \ex_mem/N237 , \ex_mem/N236 , \ex_mem/N235 , \ex_mem/N234 ,
         \ex_mem/N233 , \ex_mem/N232 , \ex_mem/N231 , \ex_mem/N230 ,
         \ex_mem/N229 , \ex_mem/N227 , \ex_mem/N226 , \ex_mem/N225 ,
         \ex_mem/N224 , \ex_mem/N223 , \ex_mem/N222 , \ex_mem/N221 ,
         \ex_mem/N220 , \ex_mem/N219 , \ex_mem/N218 , \ex_mem/N217 ,
         \ex_mem/N216 , \ex_mem/N215 , \ex_mem/N214 , \ex_mem/N213 ,
         \ex_mem/N212 , \ex_mem/N211 , \ex_mem/N210 , \ex_mem/N209 ,
         \ex_mem/N208 , \ex_mem/N207 , \ex_mem/N206 , \ex_mem/N205 ,
         \ex_mem/N204 , \ex_mem/N203 , \ex_mem/N202 , \ex_mem/N200 ,
         \ex_mem/N199 , \ex_mem/N198 , \ex_mem/N197 , \ex_mem/N196 ,
         \ex_mem/N162 , \ex_mem/N161 , \ex_mem/N160 , \ex_mem/N159 ,
         \ex_mem/N158 , \ex_mem/N157 , \ex_mem/N156 , \ex_mem/N155 ,
         \ex_mem/N154 , \ex_mem/N153 , \ex_mem/N152 , \ex_mem/N151 ,
         \ex_mem/N150 , \ex_mem/N149 , \ex_mem/N148 , \ex_mem/N147 ,
         \ex_mem/N146 , \ex_mem/N145 , \ex_mem/N144 , \ex_mem/N143 ,
         \ex_mem/N142 , \ex_mem/N141 , \ex_mem/N140 , \ex_mem/N139 ,
         \ex_mem/N138 , \ex_mem/N137 , \ex_mem/N136 , \ex_mem/N135 ,
         \ex_mem/N134 , \ex_mem/N133 , \ex_mem/N132 , \ex_mem/N131 ,
         \ex_mem/N130 , \ex_mem/N129 , \ex_mem/N128 , \ex_mem/N127 ,
         \ex_mem/N126 , \ex_mem/N125 , \ex_mem/N124 , \ex_mem/N123 ,
         \ex_mem/N122 , \ex_mem/N121 , \ex_mem/N120 , \ex_mem/N119 ,
         \ex_mem/N118 , \ex_mem/N117 , \ex_mem/N116 , \ex_mem/N115 ,
         \ex_mem/N114 , \ex_mem/N113 , \ex_mem/N112 , \ex_mem/N111 ,
         \ex_mem/N110 , \ex_mem/N109 , \ex_mem/N108 , \ex_mem/N107 ,
         \ex_mem/N106 , \ex_mem/N105 , \ex_mem/N104 , \ex_mem/N103 ,
         \ex_mem/N102 , \ex_mem/N101 , \ex_mem/N100 , \ex_mem/N99 ,
         \ex_mem/N66 , \ex_mem/N65 , \ex_mem/N64 , \ex_mem/N63 , \ex_mem/N62 ,
         \ex_mem/N61 , \ex_mem/N60 , \ex_mem/N59 , \ex_mem/N58 , \ex_mem/N57 ,
         \ex_mem/N56 , \ex_mem/N55 , \ex_mem/N54 , \ex_mem/N53 , \ex_mem/N52 ,
         \ex_mem/N51 , \ex_mem/N50 , \ex_mem/N49 , \ex_mem/N48 , \ex_mem/N47 ,
         \ex_mem/N46 , \ex_mem/N45 , \ex_mem/N44 , \ex_mem/N43 , \ex_mem/N42 ,
         \ex_mem/N41 , \ex_mem/N40 , \ex_mem/N39 , \ex_mem/N38 , \ex_mem/N37 ,
         \ex_mem/N36 , \ex_mem/N35 , \mem_wb/N41 , \mem_wb/N36 ,
         \mem/addImm/mux_map1/M1/M3/z2[31] , n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1950, n1952,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1986, n1990,
         n1992, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2083, n2084, n2086, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2116,
         n2118, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2133, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2220, n2222, n2223, n2224, n2225, n2227, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2528, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2544, n2545, n2546, n2547, n2548, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         \hazard_detect/eq_83/A[0] , \hazard_detect/eq_83/A[1] ,
         \hazard_detect/eq_83/A[2] , \hazard_detect/eq_83/A[3] ,
         \hazard_detect/eq_83/A[4] , n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3112, n3113, n3114, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3136, n3137,
         n3138, n3139, n3140, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6752, n6753, n6756, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777;
  wire   [27:0] instr_2;
  wire   [4:0] rd_2;
  wire   [4:0] rd_3;
  wire   [1:0] reg31Val_3;
  wire   [31:0] reg31Val_0;
  wire   [31:0] \wb/dsize_reg/z2 ;
  assign \mem_wb/N41  = rst;
  assign rs2[0] = \hazard_detect/eq_83/A[0] ;
  assign rs2[1] = \hazard_detect/eq_83/A[1] ;
  assign rs2[2] = \hazard_detect/eq_83/A[2] ;
  assign rs2[3] = \hazard_detect/eq_83/A[3] ;
  assign rs2[4] = \hazard_detect/eq_83/A[4] ;

  DFFR_X1 \ex_mem/aluRes_q_reg[0]  ( .D(n6111), .CK(clk), .RN(n3252), .Q(
        memAddr[0]), .QN(n6300) );
  DFFR_X1 \ex_mem/aluRes_q_reg[16]  ( .D(\ex_mem/N212 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[16]), .QN(n6299) );
  DFFR_X1 \ex_mem/aluRes_q_reg[21]  ( .D(\ex_mem/N217 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[21]), .QN(n6298) );
  DFFR_X1 \ex_mem/aluRes_q_reg[22]  ( .D(\ex_mem/N218 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[22]), .QN(n6297) );
  DFFR_X1 \ex_mem/aluRes_q_reg[23]  ( .D(\ex_mem/N219 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[23]), .QN(n6296) );
  DFFR_X1 \ex_mem/aluRes_q_reg[24]  ( .D(\ex_mem/N220 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[24]), .QN(n6295) );
  DFFR_X1 \ex_mem/aluRes_q_reg[25]  ( .D(\ex_mem/N221 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[25]), .QN(n6294) );
  DFFR_X1 \ex_mem/aluRes_q_reg[31]  ( .D(\ex_mem/N227 ), .CK(clk), .RN(n3252), 
        .Q(memAddr[31]), .QN(n6293) );
  DFFR_X1 \ex_mem/aluRes_q_reg[4]  ( .D(\ex_mem/N199 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[4]), .QN(n6292) );
  DFFR_X1 \ex_mem/aluRes_q_reg[9]  ( .D(\ex_mem/N205 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[9]), .QN(n6291) );
  DFFR_X1 \ex_mem/aluRes_q_reg[2]  ( .D(\ex_mem/N197 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[2]), .QN(n6290) );
  DFFR_X1 \ex_mem/aluRes_q_reg[1]  ( .D(\ex_mem/N196 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[1]), .QN(n6289) );
  DFFR_X1 \ex_mem/aluRes_q_reg[3]  ( .D(\ex_mem/N198 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[3]), .QN(n6288) );
  DFFR_X1 \ex_mem/aluRes_q_reg[6]  ( .D(\ex_mem/N202 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[6]), .QN(n6287) );
  DFFR_X1 \ex_mem/aluRes_q_reg[11]  ( .D(\ex_mem/N207 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[11]), .QN(n6286) );
  DFFR_X1 \ex_mem/aluRes_q_reg[7]  ( .D(\ex_mem/N203 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[7]), .QN(n6285) );
  DFFR_X1 \ex_mem/aluRes_q_reg[29]  ( .D(\ex_mem/N225 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[29]), .QN(n6284) );
  DFFR_X1 \ex_mem/aluRes_q_reg[8]  ( .D(\ex_mem/N204 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[8]), .QN(n6283) );
  DFFR_X1 \ex_mem/aluRes_q_reg[12]  ( .D(\ex_mem/N208 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[12]), .QN(n6282) );
  DFFR_X1 \ex_mem/aluRes_q_reg[13]  ( .D(\ex_mem/N209 ), .CK(clk), .RN(n3251), 
        .Q(memAddr[13]), .QN(n6281) );
  DFFR_X1 \ex_mem/aluRes_q_reg[10]  ( .D(\ex_mem/N206 ), .CK(clk), .RN(n3250), 
        .Q(memAddr[10]), .QN(n6280) );
  DFFR_X1 \ex_mem/busA_q_reg[10]  ( .D(n2761), .CK(clk), .RN(n3250), .Q(n2624)
         );
  DFFR_X1 \ex_mem/incPC_q_reg[13]  ( .D(\ex_mem/N48 ), .CK(clk), .RN(n3250), 
        .Q(n2684), .QN(n6277) );
  DFFR_X1 \ex_mem/incPC_q_reg[14]  ( .D(\ex_mem/N49 ), .CK(clk), .RN(n3250), 
        .Q(n2691), .QN(n6276) );
  DFFR_X1 \ex_mem/incPC_q_reg[15]  ( .D(\ex_mem/N50 ), .CK(clk), .RN(n3250), 
        .Q(n2682), .QN(n6275) );
  DFFR_X1 \ex_mem/incPC_q_reg[18]  ( .D(\ex_mem/N53 ), .CK(clk), .RN(n3250), 
        .Q(n2697), .QN(n6272) );
  DFFR_X1 \ex_mem/incPC_q_reg[19]  ( .D(\ex_mem/N54 ), .CK(clk), .RN(n3250), 
        .Q(n2824), .QN(n6271) );
  DFFR_X1 \ex_mem/incPC_q_reg[20]  ( .D(\ex_mem/N55 ), .CK(clk), .RN(n3249), 
        .Q(n2826), .QN(n6270) );
  DFFR_X1 \ex_mem/incPC_q_reg[21]  ( .D(\ex_mem/N56 ), .CK(clk), .RN(n3249), 
        .Q(n2821), .QN(n6269) );
  DFFR_X1 \ex_mem/incPC_q_reg[22]  ( .D(\ex_mem/N57 ), .CK(clk), .RN(n3249), 
        .Q(n2825), .QN(n6268) );
  DFFR_X1 \ex_mem/incPC_q_reg[23]  ( .D(\ex_mem/N58 ), .CK(clk), .RN(n3249), 
        .Q(n2810), .QN(n6267) );
  DFFR_X1 \ex_mem/incPC_q_reg[24]  ( .D(\ex_mem/N59 ), .CK(clk), .RN(n3249), 
        .Q(n2689), .QN(n6266) );
  DFFR_X1 \ex_mem/incPC_q_reg[25]  ( .D(\ex_mem/N60 ), .CK(clk), .RN(n3249), 
        .Q(n2681), .QN(n6265) );
  DFFR_X1 \ex_mem/incPC_q_reg[26]  ( .D(\ex_mem/N61 ), .CK(clk), .RN(n3249), 
        .Q(n2696), .QN(n6264) );
  DFFR_X1 \ex_mem/incPC_q_reg[27]  ( .D(\ex_mem/N62 ), .CK(clk), .RN(n3249), 
        .Q(n2823), .QN(n6263) );
  DFFR_X1 \ex_mem/incPC_q_reg[28]  ( .D(\ex_mem/N63 ), .CK(clk), .RN(n3249), 
        .Q(n2688), .QN(n6262) );
  DFFR_X1 \ex_mem/incPC_q_reg[29]  ( .D(\ex_mem/N64 ), .CK(clk), .RN(n3249), 
        .Q(n2822), .QN(n6261) );
  DFFR_X1 \ex_mem/incPC_q_reg[30]  ( .D(\ex_mem/N65 ), .CK(clk), .RN(n3249), 
        .QN(n6260) );
  DFFR_X1 \ex_mem/aluRes_q_reg[30]  ( .D(\ex_mem/N226 ), .CK(clk), .RN(n3249), 
        .Q(memAddr[30]), .QN(n6259) );
  DFFR_X1 \ex_mem/aluRes_q_reg[19]  ( .D(\ex_mem/N215 ), .CK(clk), .RN(n3248), 
        .Q(memAddr[19]), .QN(n6258) );
  DFFR_X1 \ex_mem/isZero_q_reg  ( .D(\ex_mem/N232 ), .CK(clk), .RN(n3248), 
        .QN(n6257) );
  DFFR_X1 \ex_mem/fp_q_reg  ( .D(n3225), .CK(clk), .RN(n3248), .Q(fp_3) );
  DFFR_X1 \ex_mem/rd_q_reg[1]  ( .D(\ex_mem/N244 ), .CK(clk), .RN(n3248), .Q(
        rd_3[1]), .QN(n2785) );
  DFFR_X1 \ex_mem/rd_q_reg[2]  ( .D(\ex_mem/N245 ), .CK(clk), .RN(n3248), .Q(
        rd_3[2]), .QN(n2784) );
  DFFR_X1 \id_ex/instr_q_reg[5]  ( .D(n6129), .CK(clk), .RN(n3248), .Q(
        instr_2[5]) );
  DFFR_X1 \id_ex/instr_q_reg[3]  ( .D(n6126), .CK(clk), .RN(n3248), .QN(n6256)
         );
  DFFR_X1 \id_ex/instr_q_reg[1]  ( .D(n6125), .CK(clk), .RN(n3248), .QN(n6255)
         );
  DFFR_X1 \id_ex/zeroExt_q_reg  ( .D(n6131), .CK(clk), .RN(n3248), .Q(
        zeroExt_2), .QN(n3041) );
  DFFR_X1 \id_ex/busA_sel_q_reg[0]  ( .D(\id_ex/N38 ), .CK(clk), .RN(n3248), 
        .QN(n6254) );
  DFFR_X1 \id_ex/memWr_q_reg  ( .D(\id_ex/N36 ), .CK(clk), .RN(n3248), .QN(
        n6253) );
  DFFR_X1 \id_ex/instr_q_reg[30]  ( .D(n6137), .CK(clk), .RN(n3248), .Q(n2846), 
        .QN(n6252) );
  DFFR_X1 \id_ex/instr_q_reg[29]  ( .D(\id_ex/N33 ), .CK(clk), .RN(n3247), .Q(
        n2797), .QN(n6251) );
  DFFR_X1 \id_ex/instr_q_reg[28]  ( .D(n6128), .CK(clk), .RN(n3247), .QN(n6250) );
  DFFR_X1 \id_ex/instr_q_reg[27]  ( .D(\id_ex/N31 ), .CK(clk), .RN(n3247), .Q(
        instr_2[27]) );
  DFFR_X1 \id_ex/instr_q_reg[26]  ( .D(\id_ex/N30 ), .CK(clk), .RN(n3247), .Q(
        instr_2[26]) );
  DFFR_X1 \id_ex/instr_q_reg[25]  ( .D(n6121), .CK(clk), .RN(n3247), .QN(n6249) );
  DFFR_X1 \id_ex/instr_q_reg[24]  ( .D(n6127), .CK(clk), .RN(n3247), .QN(n6248) );
  DFFR_X1 \id_ex/instr_q_reg[23]  ( .D(n6120), .CK(clk), .RN(n3247), .QN(n6247) );
  DFFR_X1 \id_ex/instr_q_reg[22]  ( .D(n6119), .CK(clk), .RN(n3247), .QN(n6246) );
  DFFR_X1 \id_ex/instr_q_reg[21]  ( .D(n6118), .CK(clk), .RN(n3247), .QN(n6245) );
  DFFR_X1 \id_ex/instr_q_reg[20]  ( .D(n2960), .CK(clk), .RN(n3247), .QN(n6244) );
  DFFR_X1 \id_ex/instr_q_reg[19]  ( .D(n2764), .CK(clk), .RN(n3247), .Q(
        instr_2[19]) );
  DFFR_X1 \id_ex/instr_q_reg[18]  ( .D(n2763), .CK(clk), .RN(n3247), .Q(
        instr_2[18]) );
  DFFR_X1 \id_ex/instr_q_reg[17]  ( .D(n2762), .CK(clk), .RN(n3246), .Q(
        instr_2[17]) );
  DFFR_X1 \id_ex/instr_q_reg[16]  ( .D(n2981), .CK(clk), .RN(n3246), .Q(
        instr_2[16]) );
  DFFR_X1 \id_ex/instr_q_reg[15]  ( .D(n6134), .CK(clk), .RN(n3246), .QN(n6243) );
  DFFR_X1 \id_ex/instr_q_reg[14]  ( .D(n6124), .CK(clk), .RN(n3246), .QN(n6242) );
  DFFR_X1 \id_ex/instr_q_reg[13]  ( .D(n6123), .CK(clk), .RN(n3246), .QN(n6241) );
  DFFR_X1 \id_ex/instr_q_reg[12]  ( .D(n6122), .CK(clk), .RN(n3246), .QN(n6240) );
  DFFR_X1 \id_ex/instr_q_reg[11]  ( .D(n6117), .CK(clk), .RN(n3246), .QN(n6239) );
  DFFR_X1 \id_ex/instr_q_reg[10]  ( .D(n6116), .CK(clk), .RN(n3246), .QN(n6238) );
  DFFR_X1 \id_ex/instr_q_reg[9]  ( .D(n6115), .CK(clk), .RN(n3246), .Q(
        instr_2[9]) );
  DFFR_X1 \id_ex/instr_q_reg[8]  ( .D(n6114), .CK(clk), .RN(n3246), .Q(
        instr_2[8]) );
  DFFR_X1 \id_ex/instr_q_reg[7]  ( .D(n6113), .CK(clk), .RN(n3246), .Q(
        instr_2[7]) );
  DFFR_X1 \id_ex/instr_q_reg[6]  ( .D(n6112), .CK(clk), .RN(n3246), .Q(
        instr_2[6]) );
  DFFR_X1 \id_ex/valid_q_reg  ( .D(\id_ex/N44 ), .CK(clk), .RN(n3267), .Q(
        valid_2), .QN(n2786) );
  DFFR_X1 \id_ex/instr_q_reg[31]  ( .D(n6130), .CK(clk), .RN(n3266), .Q(n2841), 
        .QN(n6236) );
  DFFR_X1 \ex_mem/rd_q_reg[0]  ( .D(\ex_mem/N243 ), .CK(clk), .RN(n3256), .Q(
        rd_3[0]), .QN(n2633) );
  DFFR_X1 \id_ex/regWr_q_reg  ( .D(\id_ex/N37 ), .CK(clk), .RN(n3264), .QN(
        n6235) );
  DFFR_X1 \ex_mem/busB_q_reg[0]  ( .D(\ex_mem/N99 ), .CK(clk), .RN(n3249), 
        .QN(n6234) );
  DFFR_X1 \ex_mem/rd_q_reg[4]  ( .D(\ex_mem/N247 ), .CK(clk), .RN(n3257), .Q(
        rd_3[4]), .QN(n2632) );
  DFFR_X1 \ex_mem/rd_q_reg[3]  ( .D(\ex_mem/N246 ), .CK(clk), .RN(n3263), .Q(
        rd_3[3]), .QN(n2598) );
  DFFR_X1 \ex_mem/valid_q_reg  ( .D(\ex_mem/N241 ), .CK(clk), .RN(n3248), .Q(
        valid_3) );
  DFFR_X1 \id_ex/memWrData_sel_q_reg[0]  ( .D(\id_ex/N42 ), .CK(clk), .RN(
        n3251), .QN(n6233) );
  DFFR_X1 \id_ex/busA_sel_q_reg[1]  ( .D(\id_ex/N39 ), .CK(clk), .RN(n3250), 
        .Q(n2888), .QN(n6231) );
  DFFR_X1 \ex_mem/memWrData_sel_q_reg[0]  ( .D(\ex_mem/N239 ), .CK(clk), .RN(
        n3265), .Q(n2664), .QN(n6230) );
  DFFR_X1 \ex_mem/op0_q_reg  ( .D(\ex_mem/N237 ), .CK(clk), .RN(n3265), .Q(
        op0_3) );
  DFFR_X1 \ex_mem/link_q_reg  ( .D(\ex_mem/N236 ), .CK(clk), .RN(n3265), .Q(
        link_3) );
  DFFR_X1 \ex_mem/jr_q_reg  ( .D(\ex_mem/N235 ), .CK(clk), .RN(n3265), .Q(
        n2596), .QN(n6229) );
  DFFR_X1 \ex_mem/branch_q_reg  ( .D(\ex_mem/N234 ), .CK(clk), .RN(n3265), 
        .QN(n6228) );
  DFFR_X1 \ex_mem/jump_q_reg  ( .D(\ex_mem/N233 ), .CK(clk), .RN(n3265), .QN(
        n6227) );
  DFFR_X1 \ex_mem/regWr_q_reg  ( .D(\ex_mem/N231 ), .CK(clk), .RN(n3265), .Q(
        \mem_wb/N36 ) );
  DFFR_X1 \ex_mem/memWr_q_reg  ( .D(\ex_mem/N230 ), .CK(clk), .RN(n3265), .Q(
        memWr) );
  DFFR_X1 \ex_mem/memRd_q_reg  ( .D(\ex_mem/N229 ), .CK(clk), .RN(n3265), .Q(
        n2635) );
  DFFR_X1 \id_ex/memWrData_sel_q_reg[1]  ( .D(n6765), .CK(clk), .RN(n3265), 
        .QN(n6226) );
  DFFR_X1 \ex_mem/memWrData_sel_q_reg[1]  ( .D(\ex_mem/N240 ), .CK(clk), .RN(
        n3264), .Q(n2601), .QN(n6225) );
  DFFR_X1 \ex_mem/busA_q_reg[31]  ( .D(n2530), .CK(clk), .RN(n3264), .QN(n6224) );
  DFFR_X1 \ex_mem/busA_q_reg[30]  ( .D(n2544), .CK(clk), .RN(n3264), .Q(n3020)
         );
  DFFR_X1 \ex_mem/busA_q_reg[29]  ( .D(n2533), .CK(clk), .RN(n3264), .Q(n3019)
         );
  DFFR_X1 \ex_mem/busA_q_reg[13]  ( .D(n2531), .CK(clk), .RN(n3264), .Q(n3005)
         );
  DFFR_X1 \ex_mem/busA_q_reg[12]  ( .D(n2553), .CK(clk), .RN(n3264), .QN(n6223) );
  DFFR_X1 \ex_mem/busA_q_reg[11]  ( .D(n2554), .CK(clk), .RN(n3264), .Q(n3006)
         );
  DFFR_X1 \ex_mem/busA_q_reg[9]  ( .D(n2539), .CK(clk), .RN(n3264), .Q(n3011)
         );
  DFFR_X1 \ex_mem/busA_q_reg[8]  ( .D(n2546), .CK(clk), .RN(n3264), .Q(n3009)
         );
  DFFR_X1 \ex_mem/busA_q_reg[7]  ( .D(n2551), .CK(clk), .RN(n3264), .Q(n3010)
         );
  DFFR_X1 \ex_mem/busA_q_reg[6]  ( .D(n2542), .CK(clk), .RN(n3264), .Q(n3007)
         );
  DFFR_X1 \ex_mem/imm32_q_reg[31]  ( .D(\ex_mem/N162 ), .CK(clk), .RN(n3264), 
        .Q(\mem/addImm/mux_map1/M1/M3/z2[31] ) );
  DFFR_X1 \ex_mem/imm32_q_reg[30]  ( .D(\ex_mem/N161 ), .CK(clk), .RN(n3263), 
        .QN(n6222) );
  DFFR_X1 \ex_mem/imm32_q_reg[29]  ( .D(\ex_mem/N160 ), .CK(clk), .RN(n3263), 
        .QN(n6221) );
  DFFR_X1 \ex_mem/imm32_q_reg[28]  ( .D(\ex_mem/N159 ), .CK(clk), .RN(n3263), 
        .Q(n2909), .QN(n6220) );
  DFFR_X1 \ex_mem/imm32_q_reg[27]  ( .D(\ex_mem/N158 ), .CK(clk), .RN(n3263), 
        .QN(n6219) );
  DFFR_X1 \ex_mem/imm32_q_reg[26]  ( .D(\ex_mem/N157 ), .CK(clk), .RN(n3263), 
        .Q(n2910), .QN(n6218) );
  DFFR_X1 \ex_mem/imm32_q_reg[25]  ( .D(\ex_mem/N156 ), .CK(clk), .RN(n3263), 
        .Q(n2911), .QN(n6217) );
  DFFR_X1 \ex_mem/imm32_q_reg[24]  ( .D(\ex_mem/N155 ), .CK(clk), .RN(n3263), 
        .Q(n2912), .QN(n6216) );
  DFFR_X1 \ex_mem/imm32_q_reg[23]  ( .D(\ex_mem/N154 ), .CK(clk), .RN(n3263), 
        .QN(n6215) );
  DFFR_X1 \ex_mem/imm32_q_reg[22]  ( .D(\ex_mem/N153 ), .CK(clk), .RN(n3263), 
        .QN(n6214) );
  DFFR_X1 \ex_mem/imm32_q_reg[21]  ( .D(\ex_mem/N152 ), .CK(clk), .RN(n3263), 
        .QN(n6213) );
  DFFR_X1 \ex_mem/imm32_q_reg[20]  ( .D(\ex_mem/N151 ), .CK(clk), .RN(n3263), 
        .QN(n6212) );
  DFFR_X1 \ex_mem/imm32_q_reg[19]  ( .D(\ex_mem/N150 ), .CK(clk), .RN(n3263), 
        .QN(n6211) );
  DFFR_X1 \ex_mem/imm32_q_reg[18]  ( .D(\ex_mem/N149 ), .CK(clk), .RN(n3262), 
        .Q(n2913), .QN(n6210) );
  DFFR_X1 \ex_mem/imm32_q_reg[15]  ( .D(\ex_mem/N146 ), .CK(clk), .RN(n3262), 
        .Q(n2914), .QN(n6207) );
  DFFR_X1 \ex_mem/imm32_q_reg[14]  ( .D(\ex_mem/N145 ), .CK(clk), .RN(n3262), 
        .Q(n2921), .QN(n6206) );
  DFFR_X1 \ex_mem/imm32_q_reg[13]  ( .D(\ex_mem/N144 ), .CK(clk), .RN(n3262), 
        .Q(n2920), .QN(n6205) );
  DFFR_X1 \ex_mem/imm32_q_reg[12]  ( .D(\ex_mem/N143 ), .CK(clk), .RN(n3262), 
        .Q(n2917), .QN(n6204) );
  DFFR_X1 \ex_mem/imm32_q_reg[9]  ( .D(\ex_mem/N140 ), .CK(clk), .RN(n3262), 
        .Q(n2916), .QN(n6201) );
  DFFR_X1 \ex_mem/imm32_q_reg[8]  ( .D(\ex_mem/N139 ), .CK(clk), .RN(n3262), 
        .Q(n2918), .QN(n6200) );
  DFFR_X1 \ex_mem/imm32_q_reg[7]  ( .D(\ex_mem/N138 ), .CK(clk), .RN(n3262), 
        .Q(n2919), .QN(n6199) );
  DFFR_X1 \ex_mem/imm32_q_reg[6]  ( .D(\ex_mem/N137 ), .CK(clk), .RN(n3261), 
        .Q(n2952), .QN(n6198) );
  DFFR_X1 \ex_mem/imm32_q_reg[5]  ( .D(\ex_mem/N136 ), .CK(clk), .RN(n3261), 
        .Q(n2951), .QN(n6197) );
  DFFR_X1 \ex_mem/imm32_q_reg[4]  ( .D(\ex_mem/N135 ), .CK(clk), .RN(n3261), 
        .QN(n6196) );
  DFFR_X1 \ex_mem/imm32_q_reg[3]  ( .D(\ex_mem/N134 ), .CK(clk), .RN(n3261), 
        .Q(n2915), .QN(n6195) );
  DFFR_X1 \ex_mem/imm32_q_reg[2]  ( .D(\ex_mem/N133 ), .CK(clk), .RN(n3261), 
        .QN(n6194) );
  DFFR_X1 \ex_mem/imm32_q_reg[1]  ( .D(\ex_mem/N132 ), .CK(clk), .RN(n3261), 
        .Q(n2953), .QN(n6193) );
  DFFR_X1 \ex_mem/imm32_q_reg[0]  ( .D(\ex_mem/N131 ), .CK(clk), .RN(n3261), 
        .Q(n2840) );
  DFFR_X1 \ex_mem/busA_q_reg[0]  ( .D(n6733), .CK(clk), .RN(n3261), .QN(n6192)
         );
  DFFR_X1 \ex_mem/busA_q_reg[1]  ( .D(n6734), .CK(clk), .RN(n3261), .QN(n6191)
         );
  DFFR_X1 \ex_mem/busA_q_reg[2]  ( .D(n2534), .CK(clk), .RN(n3260), .Q(n2903)
         );
  DFFR_X1 \ex_mem/busA_q_reg[3]  ( .D(n2558), .CK(clk), .RN(n3260), .Q(n2902)
         );
  DFFR_X1 \ex_mem/busA_q_reg[4]  ( .D(n2557), .CK(clk), .RN(n3260), .Q(n2901)
         );
  DFFR_X1 \ex_mem/incPC_q_reg[8]  ( .D(\ex_mem/N43 ), .CK(clk), .RN(n3260), 
        .Q(n2690), .QN(n6185) );
  DFFR_X1 \ex_mem/incPC_q_reg[9]  ( .D(\ex_mem/N44 ), .CK(clk), .RN(n3260), 
        .QN(n6184) );
  DFFR_X1 \ex_mem/incPC_q_reg[12]  ( .D(\ex_mem/N47 ), .CK(clk), .RN(n3260), 
        .Q(n2698), .QN(n6183) );
  DFFR_X1 \ex_mem/aluRes_q_reg[28]  ( .D(\ex_mem/N224 ), .CK(clk), .RN(n3260), 
        .Q(memAddr[28]), .QN(n6182) );
  DFFR_X1 \ex_mem/busA_q_reg[28]  ( .D(n2559), .CK(clk), .RN(n3259), .Q(n3018)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[27]  ( .D(\ex_mem/N223 ), .CK(clk), .RN(n3259), 
        .Q(memAddr[27]), .QN(n6181) );
  DFFR_X1 \ex_mem/busA_q_reg[27]  ( .D(n2556), .CK(clk), .RN(n3259), .Q(n3017)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[26]  ( .D(\ex_mem/N222 ), .CK(clk), .RN(n3259), 
        .Q(memAddr[26]), .QN(n6180) );
  DFFR_X1 \ex_mem/busA_q_reg[26]  ( .D(n2535), .CK(clk), .RN(n3259), .QN(n6179) );
  DFFR_X1 \ex_mem/aluRes_q_reg[5]  ( .D(\ex_mem/N200 ), .CK(clk), .RN(n3259), 
        .Q(memAddr[5]), .QN(n6178) );
  DFFR_X1 \ex_mem/busA_q_reg[5]  ( .D(n2536), .CK(clk), .RN(n3259), .Q(n3008)
         );
  DFFR_X1 \ex_mem/busA_q_reg[25]  ( .D(n2541), .CK(clk), .RN(n3259), .Q(n3002)
         );
  DFFR_X1 \ex_mem/busA_q_reg[24]  ( .D(n2550), .CK(clk), .RN(n3259), .Q(n3000)
         );
  DFFR_X1 \ex_mem/busA_q_reg[23]  ( .D(n2545), .CK(clk), .RN(n3259), .Q(n3001)
         );
  DFFR_X1 \ex_mem/busA_q_reg[22]  ( .D(n2540), .CK(clk), .RN(n3259), .Q(n3012)
         );
  DFFR_X1 \ex_mem/busA_q_reg[21]  ( .D(n2528), .CK(clk), .RN(n3258), .Q(n3015)
         );
  DFFR_X1 \ex_mem/busA_q_reg[16]  ( .D(n2548), .CK(clk), .RN(n3258), .Q(n2999)
         );
  DFFR_X1 \ex_mem/busA_q_reg[14]  ( .D(n2538), .CK(clk), .RN(n3258), .Q(n3004)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[20]  ( .D(\ex_mem/N216 ), .CK(clk), .RN(n3258), 
        .Q(memAddr[20]), .QN(n6175) );
  DFFR_X1 \ex_mem/busA_q_reg[20]  ( .D(n2555), .CK(clk), .RN(n3258), .Q(n3013)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[15]  ( .D(\ex_mem/N211 ), .CK(clk), .RN(n3258), 
        .Q(memAddr[15]), .QN(n6174) );
  DFFR_X1 \ex_mem/busA_q_reg[15]  ( .D(n2547), .CK(clk), .RN(n3258), .Q(n3003)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[18]  ( .D(\ex_mem/N214 ), .CK(clk), .RN(n3258), 
        .Q(memAddr[18]), .QN(n6173) );
  DFFR_X1 \ex_mem/busA_q_reg[18]  ( .D(n2532), .CK(clk), .RN(n3258), .Q(n3014)
         );
  DFFR_X1 \ex_mem/aluRes_q_reg[17]  ( .D(\ex_mem/N213 ), .CK(clk), .RN(n3258), 
        .Q(memAddr[17]), .QN(n6172) );
  DFFR_X1 \ex_mem/busA_q_reg[17]  ( .D(n2537), .CK(clk), .RN(n3258), .Q(n3016)
         );
  DFFR_X1 \ex_mem/busB_q_reg[28]  ( .D(\ex_mem/N127 ), .CK(clk), .RN(n3257), 
        .QN(n6171) );
  DFFR_X1 \ex_mem/busB_q_reg[27]  ( .D(\ex_mem/N126 ), .CK(clk), .RN(n3257), 
        .QN(n6170) );
  DFFR_X1 \ex_mem/busB_q_reg[26]  ( .D(\ex_mem/N125 ), .CK(clk), .RN(n3257), 
        .QN(n6169) );
  DFFR_X1 \ex_mem/busB_q_reg[20]  ( .D(\ex_mem/N119 ), .CK(clk), .RN(n3257), 
        .QN(n6168) );
  DFFR_X1 \ex_mem/busB_q_reg[18]  ( .D(\ex_mem/N117 ), .CK(clk), .RN(n3257), 
        .QN(n6167) );
  DFFR_X1 \ex_mem/busB_q_reg[17]  ( .D(\ex_mem/N116 ), .CK(clk), .RN(n3257), 
        .QN(n6166) );
  DFFR_X1 \ex_mem/busB_q_reg[15]  ( .D(\ex_mem/N114 ), .CK(clk), .RN(n3257), 
        .QN(n6165) );
  DFFR_X1 \ex_mem/busB_q_reg[14]  ( .D(\ex_mem/N113 ), .CK(clk), .RN(n3257), 
        .QN(n6164) );
  DFFR_X1 \ex_mem/busB_q_reg[5]  ( .D(\ex_mem/N104 ), .CK(clk), .RN(n3257), 
        .QN(n6163) );
  DFFR_X1 \ex_mem/busA_q_reg[19]  ( .D(n2552), .CK(clk), .RN(n3257), .QN(n6162) );
  DFFR_X1 \ex_mem/busB_q_reg[19]  ( .D(\ex_mem/N118 ), .CK(clk), .RN(n3257), 
        .QN(n6161) );
  DFFR_X1 \ex_mem/busB_q_reg[30]  ( .D(\ex_mem/N129 ), .CK(clk), .RN(n3257), 
        .QN(n6160) );
  DFFR_X1 \ex_mem/incPC_q_reg[31]  ( .D(\ex_mem/N66 ), .CK(clk), .RN(n3256), 
        .QN(n6159) );
  DFFR_X1 \ex_mem/busB_q_reg[10]  ( .D(\ex_mem/N109 ), .CK(clk), .RN(n3256), 
        .QN(n6158) );
  DFFR_X1 \ex_mem/busB_q_reg[13]  ( .D(\ex_mem/N112 ), .CK(clk), .RN(n3256), 
        .QN(n6157) );
  DFFR_X1 \ex_mem/busB_q_reg[12]  ( .D(\ex_mem/N111 ), .CK(clk), .RN(n3256), 
        .QN(n6156) );
  DFFR_X1 \ex_mem/busB_q_reg[8]  ( .D(\ex_mem/N107 ), .CK(clk), .RN(n3256), 
        .QN(n6155) );
  DFFR_X1 \ex_mem/busB_q_reg[29]  ( .D(\ex_mem/N128 ), .CK(clk), .RN(n3256), 
        .QN(n6154) );
  DFFR_X1 \ex_mem/busB_q_reg[11]  ( .D(\ex_mem/N110 ), .CK(clk), .RN(n3256), 
        .QN(n6153) );
  DFFR_X1 \ex_mem/busB_q_reg[6]  ( .D(\ex_mem/N105 ), .CK(clk), .RN(n3256), 
        .QN(n6152) );
  DFFR_X1 \ex_mem/busB_q_reg[3]  ( .D(\ex_mem/N102 ), .CK(clk), .RN(n3256), 
        .QN(n6151) );
  DFFR_X1 \ex_mem/busB_q_reg[1]  ( .D(\ex_mem/N100 ), .CK(clk), .RN(n3256), 
        .QN(n6150) );
  DFFR_X1 \ex_mem/busB_q_reg[2]  ( .D(\ex_mem/N101 ), .CK(clk), .RN(n3256), 
        .QN(n6149) );
  DFFR_X1 \ex_mem/busB_q_reg[9]  ( .D(\ex_mem/N108 ), .CK(clk), .RN(n3256), 
        .QN(n6148) );
  DFFR_X1 \ex_mem/busB_q_reg[4]  ( .D(\ex_mem/N103 ), .CK(clk), .RN(n3255), 
        .QN(n6147) );
  DFFR_X1 \ex_mem/busB_q_reg[31]  ( .D(\ex_mem/N130 ), .CK(clk), .RN(n3255), 
        .QN(n6146) );
  DFFR_X1 \ex_mem/busB_q_reg[25]  ( .D(\ex_mem/N124 ), .CK(clk), .RN(n3255), 
        .QN(n6145) );
  DFFR_X1 \ex_mem/busB_q_reg[24]  ( .D(\ex_mem/N123 ), .CK(clk), .RN(n3255), 
        .QN(n6144) );
  DFFR_X1 \ex_mem/busB_q_reg[23]  ( .D(\ex_mem/N122 ), .CK(clk), .RN(n3255), 
        .QN(n6143) );
  DFFR_X1 \ex_mem/busB_q_reg[22]  ( .D(\ex_mem/N121 ), .CK(clk), .RN(n3255), 
        .QN(n6142) );
  DFFR_X1 \ex_mem/busB_q_reg[21]  ( .D(\ex_mem/N120 ), .CK(clk), .RN(n3260), 
        .QN(n6141) );
  DFFR_X1 \ex_mem/busB_q_reg[16]  ( .D(\ex_mem/N115 ), .CK(clk), .RN(n3252), 
        .QN(n6140) );
  DFFR_X1 \ex_mem/busB_q_reg[7]  ( .D(\ex_mem/N106 ), .CK(clk), .RN(n3255), 
        .QN(n6139) );
  DFFR_X1 \if_id/incPC_q_reg[10]  ( .D(n2214), .CK(clk), .RN(n3255), .Q(n2949)
         );
  DFFR_X1 \id_ex/incPC_q_reg[10]  ( .D(n2213), .CK(clk), .RN(n3270), .Q(n2756), 
        .QN(n6548) );
  DFFR_X1 \if_id/incPC_q_reg[11]  ( .D(n2212), .CK(clk), .RN(n3268), .Q(n2948)
         );
  DFFR_X1 \id_ex/incPC_q_reg[11]  ( .D(n2211), .CK(clk), .RN(n3273), .Q(n2755), 
        .QN(n6547) );
  DFFR_X1 \if_id/incPC_q_reg[13]  ( .D(n2210), .CK(clk), .RN(n3268), .Q(n2947)
         );
  DFFR_X1 \id_ex/incPC_q_reg[13]  ( .D(n2209), .CK(clk), .RN(n3273), .Q(n2754), 
        .QN(n6546) );
  DFFR_X1 \if_id/incPC_q_reg[14]  ( .D(n2208), .CK(clk), .RN(n3255), .Q(n2946)
         );
  DFFR_X1 \id_ex/incPC_q_reg[14]  ( .D(n2207), .CK(clk), .RN(n3269), .Q(n2753), 
        .QN(n6545) );
  DFFR_X1 \if_id/incPC_q_reg[15]  ( .D(n2206), .CK(clk), .RN(n3268), .Q(n2945)
         );
  DFFR_X1 \id_ex/incPC_q_reg[15]  ( .D(n2205), .CK(clk), .RN(n3273), .Q(n2752), 
        .QN(n6544) );
  DFFR_X1 \if_id/incPC_q_reg[16]  ( .D(n2204), .CK(clk), .RN(n3255), .Q(n2944)
         );
  DFFR_X1 \id_ex/incPC_q_reg[16]  ( .D(n2203), .CK(clk), .RN(n3269), .Q(n2751), 
        .QN(n6543) );
  DFFR_X1 \if_id/incPC_q_reg[17]  ( .D(n2202), .CK(clk), .RN(n3267), .Q(n2943)
         );
  DFFR_X1 \id_ex/incPC_q_reg[17]  ( .D(n2201), .CK(clk), .RN(n3273), .Q(n2750), 
        .QN(n6542) );
  DFFR_X1 \if_id/incPC_q_reg[18]  ( .D(n2200), .CK(clk), .RN(n3254), .Q(n2942)
         );
  DFFR_X1 \id_ex/incPC_q_reg[18]  ( .D(n2199), .CK(clk), .RN(n3269), .Q(n2749), 
        .QN(n6541) );
  DFFR_X1 \if_id/incPC_q_reg[19]  ( .D(n2198), .CK(clk), .RN(n3267), .Q(n2941)
         );
  DFFR_X1 \id_ex/incPC_q_reg[19]  ( .D(n2197), .CK(clk), .RN(n3273), .Q(n2748), 
        .QN(n6540) );
  DFFR_X1 \if_id/incPC_q_reg[20]  ( .D(n2196), .CK(clk), .RN(n3267), .Q(n2759)
         );
  DFFR_X1 \id_ex/incPC_q_reg[20]  ( .D(n2195), .CK(clk), .RN(n3273), .Q(n2899), 
        .QN(n6539) );
  DFFR_X1 \if_id/incPC_q_reg[21]  ( .D(n2194), .CK(clk), .RN(n3254), .Q(n2940)
         );
  DFFR_X1 \id_ex/incPC_q_reg[21]  ( .D(n2193), .CK(clk), .RN(n3269), .Q(n2747), 
        .QN(n6538) );
  DFFR_X1 \if_id/incPC_q_reg[22]  ( .D(n2192), .CK(clk), .RN(n3267), .Q(n2939)
         );
  DFFR_X1 \id_ex/incPC_q_reg[22]  ( .D(n2191), .CK(clk), .RN(n3273), .Q(n2746), 
        .QN(n6537) );
  DFFR_X1 \if_id/incPC_q_reg[23]  ( .D(n2190), .CK(clk), .RN(n3254), .Q(n2938)
         );
  DFFR_X1 \id_ex/incPC_q_reg[23]  ( .D(n2189), .CK(clk), .RN(n3269), .Q(n2745), 
        .QN(n6536) );
  DFFR_X1 \if_id/incPC_q_reg[24]  ( .D(n2188), .CK(clk), .RN(n3267), .Q(n2937)
         );
  DFFR_X1 \id_ex/incPC_q_reg[24]  ( .D(n2187), .CK(clk), .RN(n3273), .Q(n2744), 
        .QN(n6535) );
  DFFR_X1 \if_id/incPC_q_reg[25]  ( .D(n2186), .CK(clk), .RN(n3254), .Q(n2936)
         );
  DFFR_X1 \id_ex/incPC_q_reg[25]  ( .D(n2185), .CK(clk), .RN(n3269), .Q(n2743), 
        .QN(n6534) );
  DFFR_X1 \if_id/incPC_q_reg[26]  ( .D(n2184), .CK(clk), .RN(n3267), .Q(n2935)
         );
  DFFR_X1 \id_ex/incPC_q_reg[26]  ( .D(n2183), .CK(clk), .RN(n3273), .Q(n2742), 
        .QN(n6533) );
  DFFR_X1 \if_id/incPC_q_reg[27]  ( .D(n2182), .CK(clk), .RN(n3254), .Q(n2934)
         );
  DFFR_X1 \id_ex/incPC_q_reg[27]  ( .D(n2181), .CK(clk), .RN(n3269), .Q(n2741), 
        .QN(n6532) );
  DFFR_X1 \if_id/incPC_q_reg[28]  ( .D(n2180), .CK(clk), .RN(n3267), .Q(n2933)
         );
  DFFR_X1 \id_ex/incPC_q_reg[28]  ( .D(n2179), .CK(clk), .RN(n3273), .Q(n2740), 
        .QN(n6531) );
  DFFR_X1 \if_id/incPC_q_reg[29]  ( .D(n2178), .CK(clk), .RN(n3254), .Q(n2932)
         );
  DFFR_X1 \id_ex/incPC_q_reg[29]  ( .D(n2177), .CK(clk), .RN(n3269), .Q(n2739), 
        .QN(n6530) );
  DFFR_X1 \if_id/incPC_q_reg[30]  ( .D(n2176), .CK(clk), .RN(n3254), .Q(n2931)
         );
  DFFR_X1 \id_ex/incPC_q_reg[30]  ( .D(n2175), .CK(clk), .RN(n3269), .Q(n2738), 
        .QN(n6529) );
  DFFR_X1 \if_id/instr_q_reg[31]  ( .D(n2170), .CK(clk), .RN(n3266), .Q(n2662), 
        .QN(n6588) );
  DFFR_X1 \if_id/instr_q_reg[30]  ( .D(n2169), .CK(clk), .RN(n3253), .Q(n2650), 
        .QN(n6594) );
  DFFR_X1 \if_id/instr_q_reg[29]  ( .D(n2168), .CK(clk), .RN(n3253), .Q(n2780), 
        .QN(n6590) );
  DFFR_X1 \if_id/instr_q_reg[28]  ( .D(n2167), .CK(clk), .RN(n3266), .Q(n2597), 
        .QN(n6587) );
  DFFR_X1 \if_id/instr_q_reg[26]  ( .D(n2165), .CK(clk), .RN(n3266), .Q(op0_1), 
        .QN(n2630) );
  DFFR_X1 \if_id/instr_q_reg[25]  ( .D(n2164), .CK(clk), .RN(n3253), .Q(rs1[4]), .QN(n2831) );
  DFFR_X1 \if_id/instr_q_reg[24]  ( .D(n2163), .CK(clk), .RN(n3266), .Q(rs1[3]), .QN(n2709) );
  DFFR_X1 \if_id/instr_q_reg[23]  ( .D(n2162), .CK(clk), .RN(n3253), .Q(rs1[2]), .QN(n2834) );
  DFFR_X1 \if_id/instr_q_reg[22]  ( .D(n2161), .CK(clk), .RN(n3266), .Q(rs1[1]), .QN(n2835) );
  DFFR_X1 \if_id/instr_q_reg[21]  ( .D(n2160), .CK(clk), .RN(n3253), .Q(rs1[0]), .QN(n2832) );
  DFFR_X1 \if_id/instr_q_reg[20]  ( .D(n2159), .CK(clk), .RN(n3266), .Q(n2661), 
        .QN(n6528) );
  DFFR_X1 \if_id/instr_q_reg[19]  ( .D(n2158), .CK(clk), .RN(n3266), .Q(n2972)
         );
  DFFR_X1 \if_id/instr_q_reg[18]  ( .D(n2157), .CK(clk), .RN(n3253), .Q(n2973)
         );
  DFFR_X1 \if_id/instr_q_reg[17]  ( .D(n2156), .CK(clk), .RN(n3266), .Q(n2974)
         );
  DFFR_X1 \if_id/instr_q_reg[16]  ( .D(n2155), .CK(clk), .RN(n3253), .Q(n2975)
         );
  DFFR_X1 \if_id/instr_q_reg[15]  ( .D(n2154), .CK(clk), .RN(n3266), .Q(n2679), 
        .QN(n6553) );
  DFFR_X1 \if_id/instr_q_reg[14]  ( .D(n2153), .CK(clk), .RN(n3253), .Q(n2883)
         );
  DFFR_X1 \if_id/instr_q_reg[13]  ( .D(n2152), .CK(clk), .RN(n3266), .Q(n2884)
         );
  DFFR_X1 \if_id/instr_q_reg[12]  ( .D(n2151), .CK(clk), .RN(n3253), .Q(n2885)
         );
  DFFR_X1 \if_id/instr_q_reg[11]  ( .D(n2150), .CK(clk), .RN(n3266), .Q(n2886)
         );
  DFFR_X1 \if_id/instr_q_reg[10]  ( .D(n2149), .CK(clk), .RN(n3253), .Q(n2678), 
        .QN(n6527) );
  DFFR_X1 \if_id/instr_q_reg[9]  ( .D(n2148), .CK(clk), .RN(n3252), .Q(n2955), 
        .QN(n6549) );
  DFFR_X1 \if_id/instr_q_reg[8]  ( .D(n2147), .CK(clk), .RN(n3265), .Q(n2956), 
        .QN(n6550) );
  DFFR_X1 \if_id/instr_q_reg[7]  ( .D(n2146), .CK(clk), .RN(n3252), .Q(n2957), 
        .QN(n6551) );
  DFFR_X1 \if_id/instr_q_reg[6]  ( .D(n2145), .CK(clk), .RN(n3266), .Q(n2958), 
        .QN(n6552) );
  DFFR_X1 \if_id/instr_q_reg[5]  ( .D(n2144), .CK(clk), .RN(n3252), .Q(n2604), 
        .QN(n6591) );
  DFFR_X1 \if_id/instr_q_reg[3]  ( .D(n2142), .CK(clk), .RN(n3252), .Q(n2649), 
        .QN(n6593) );
  DFFR_X1 \if_id/instr_q_reg[1]  ( .D(n2140), .CK(clk), .RN(n3253), .Q(n2636), 
        .QN(n6592) );
  DFFR_X1 \id_ex/rd_q_reg[0]  ( .D(n2138), .CK(clk), .RN(n3268), .Q(rd_2[0]), 
        .QN(n2781) );
  DFFR_X1 \id_ex/aluCtrl_q_reg[3]  ( .D(n2137), .CK(clk), .RN(n3278), .Q(n2595), .QN(n6618) );
  DFFR_X1 \id_ex/setInv_q_reg  ( .D(n2135), .CK(clk), .RN(n3255), .Q(setInv_2)
         );
  DFFR_X1 \id_ex/memRd_q_reg  ( .D(n6772), .CK(clk), .RN(n3268), .QN(n6598) );
  DFFR_X1 \id_ex/branch_q_reg  ( .D(n2133), .CK(clk), .RN(n3278), .QN(n6526)
         );
  DFFR_X1 \id_ex/jr_q_reg  ( .D(n6771), .CK(clk), .RN(n3272), .QN(n6597) );
  DFFR_X1 \id_ex/jump_q_reg  ( .D(n2131), .CK(clk), .RN(n3268), .Q(n2737), 
        .QN(n6525) );
  DFFR_X1 \id_ex/link_q_reg  ( .D(n2130), .CK(clk), .RN(n3272), .Q(n2798), 
        .QN(n6524) );
  DFFR_X1 \id_ex/fp_q_reg  ( .D(n2129), .CK(clk), .RN(n3270), .Q(n2872), .QN(
        n6599) );
  DFFR_X1 \id_ex/op0_q_reg  ( .D(n2127), .CK(clk), .RN(n3272), .Q(op0_2), .QN(
        n2878) );
  DFFR_X1 \id_ex/dSize_q_reg[0]  ( .D(n2126), .CK(clk), .RN(n3270), .Q(n2758)
         );
  DFFR_X1 \id_ex/dSize_q_reg[1]  ( .D(n2123), .CK(clk), .RN(n3275), .Q(n2757)
         );
  DFFR_X1 \id_ex/imm32_q_reg[0]  ( .D(n2120), .CK(clk), .RN(n3275), .QN(n6616)
         );
  DFFR_X1 \id_ex/imm32_q_reg[1]  ( .D(n6775), .CK(clk), .RN(n3268), .QN(n6636)
         );
  DFFR_X1 \id_ex/imm32_q_reg[2]  ( .D(n2118), .CK(clk), .RN(n3274), .Q(n2833), 
        .QN(n6601) );
  DFFR_X1 \id_ex/imm32_q_reg[3]  ( .D(n6777), .CK(clk), .RN(n3269), .QN(n6635)
         );
  DFFR_X1 \id_ex/imm32_q_reg[4]  ( .D(n2116), .CK(clk), .RN(n3274), .Q(n2838), 
        .QN(n6602) );
  DFFR_X1 \id_ex/imm32_q_reg[5]  ( .D(n6773), .CK(clk), .RN(n3253), .QN(n6634)
         );
  DFFR_X1 \id_ex/imm32_q_reg[6]  ( .D(n6766), .CK(clk), .RN(n3274), .QN(n6633)
         );
  DFFR_X1 \id_ex/imm32_q_reg[7]  ( .D(n6767), .CK(clk), .RN(n3276), .Q(n2839), 
        .QN(n6632) );
  DFFR_X1 \id_ex/imm32_q_reg[8]  ( .D(n6768), .CK(clk), .RN(n3273), .QN(n6631)
         );
  DFFR_X1 \id_ex/imm32_q_reg[9]  ( .D(n6769), .CK(clk), .RN(n3258), .QN(n6630)
         );
  DFFR_X1 \id_ex/imm32_q_reg[10]  ( .D(n6770), .CK(clk), .RN(n3270), .QN(n6629) );
  DFFR_X1 \id_ex/imm32_q_reg[11]  ( .D(n2109), .CK(clk), .RN(n3275), .Q(n2855), 
        .QN(n6606) );
  DFFR_X1 \id_ex/imm32_q_reg[12]  ( .D(n2108), .CK(clk), .RN(n3270), .QN(n6607) );
  DFFR_X1 \id_ex/imm32_q_reg[13]  ( .D(n2107), .CK(clk), .RN(n3275), .QN(n6604) );
  DFFR_X1 \id_ex/imm32_q_reg[14]  ( .D(n2106), .CK(clk), .RN(n3270), .Q(n2854), 
        .QN(n6608) );
  DFFR_X1 \id_ex/imm32_q_reg[15]  ( .D(n2105), .CK(clk), .RN(n3274), .QN(n6609) );
  DFFR_X1 \id_ex/imm32_q_reg[16]  ( .D(n2104), .CK(clk), .RN(n3270), .Q(n2861), 
        .QN(n6628) );
  DFFR_X1 \id_ex/imm32_q_reg[17]  ( .D(n2103), .CK(clk), .RN(n3274), .Q(n2866), 
        .QN(n6627) );
  DFFR_X1 \id_ex/imm32_q_reg[18]  ( .D(n2102), .CK(clk), .RN(n3270), .Q(n2860), 
        .QN(n6626) );
  DFFR_X1 \id_ex/imm32_q_reg[19]  ( .D(n2101), .CK(clk), .RN(n3274), .Q(n2862), 
        .QN(n6625) );
  DFFR_X1 \id_ex/imm32_q_reg[20]  ( .D(n2100), .CK(clk), .RN(n3274), .Q(n2868), 
        .QN(n6624) );
  DFFR_X1 \id_ex/imm32_q_reg[21]  ( .D(n2099), .CK(clk), .RN(n3277), .Q(n2865), 
        .QN(n6623) );
  DFFR_X1 \id_ex/imm32_q_reg[22]  ( .D(n2098), .CK(clk), .RN(n3274), .Q(n2873), 
        .QN(n6622) );
  DFFR_X1 \id_ex/imm32_q_reg[23]  ( .D(n2097), .CK(clk), .RN(n3273), .Q(n2716), 
        .QN(n6621) );
  DFFR_X1 \id_ex/imm32_q_reg[24]  ( .D(n2096), .CK(clk), .RN(n3274), .Q(n2867), 
        .QN(n6620) );
  DFFR_X1 \id_ex/imm32_q_reg[25]  ( .D(n2095), .CK(clk), .RN(n3272), .Q(n2863), 
        .QN(n6619) );
  DFFR_X1 \id_ex/imm32_q_reg[26]  ( .D(n2094), .CK(clk), .RN(n3274), .Q(n2859), 
        .QN(n6611) );
  DFFR_X1 \id_ex/imm32_q_reg[27]  ( .D(n2093), .CK(clk), .RN(n3275), .Q(n2869), 
        .QN(n6610) );
  DFFR_X1 \id_ex/imm32_q_reg[28]  ( .D(n2092), .CK(clk), .RN(n3274), .Q(n2858), 
        .QN(n6613) );
  DFFR_X1 \id_ex/imm32_q_reg[29]  ( .D(n2091), .CK(clk), .RN(n3271), .Q(n2864), 
        .QN(n6614) );
  DFFR_X1 \id_ex/imm32_q_reg[30]  ( .D(n2090), .CK(clk), .RN(n3274), .Q(n2713), 
        .QN(n6612) );
  DFFR_X1 \id_ex/imm32_q_reg[31]  ( .D(n2089), .CK(clk), .RN(n3274), .QN(n6605) );
  DFFR_X1 \id_ex/rd_q_reg[1]  ( .D(n2088), .CK(clk), .RN(n3272), .Q(rd_2[1]), 
        .QN(n2628) );
  DFFR_X1 \id_ex/rd_q_reg[2]  ( .D(n2086), .CK(clk), .RN(n3268), .Q(rd_2[2]), 
        .QN(n2629) );
  DFFR_X1 \id_ex/rd_q_reg[3]  ( .D(n2084), .CK(clk), .RN(n3275), .Q(rd_2[3]), 
        .QN(n2593) );
  DFFR_X1 \id_ex/rd_q_reg[4]  ( .D(n2083), .CK(clk), .RN(n3268), .Q(rd_2[4]), 
        .QN(n2782) );
  DFFR_X1 \id_ex/busA_q_reg[0]  ( .D(n6700), .CK(clk), .RN(n3278), .Q(n2648)
         );
  DFFR_X1 \id_ex/busA_q_reg[1]  ( .D(n6699), .CK(clk), .RN(n3277), .Q(n2647)
         );
  DFFR_X1 \id_ex/busA_q_reg[2]  ( .D(n6698), .CK(clk), .RN(n3279), .Q(n2646)
         );
  DFFR_X1 \id_ex/busA_q_reg[3]  ( .D(n6697), .CK(clk), .RN(n3277), .Q(n2809), 
        .QN(n6572) );
  DFFR_X1 \id_ex/busA_q_reg[4]  ( .D(n6696), .CK(clk), .RN(n3272), .Q(n2796), 
        .QN(n6571) );
  DFFR_X1 \id_ex/busA_q_reg[5]  ( .D(n6695), .CK(clk), .RN(n3276), .Q(n2791), 
        .QN(n6570) );
  DFFR_X1 \id_ex/busA_q_reg[6]  ( .D(n6694), .CK(clk), .RN(n3272), .Q(n2795), 
        .QN(n6569) );
  DFFR_X1 \id_ex/busA_q_reg[7]  ( .D(n6693), .CK(clk), .RN(n3276), .Q(n2794), 
        .QN(n6568) );
  DFFR_X1 \id_ex/busA_q_reg[8]  ( .D(n6692), .CK(clk), .RN(n3271), .Q(n2793), 
        .QN(n6567) );
  DFFR_X1 \id_ex/busA_q_reg[9]  ( .D(n6691), .CK(clk), .RN(n3276), .Q(n2600)
         );
  DFFR_X1 \id_ex/busA_q_reg[10]  ( .D(n6690), .CK(clk), .RN(n3278), .Q(n2645)
         );
  DFFR_X1 \id_ex/busA_q_reg[11]  ( .D(n6689), .CK(clk), .RN(n3278), .Q(n2644)
         );
  DFFR_X1 \id_ex/busA_q_reg[12]  ( .D(n6688), .CK(clk), .RN(n3277), .Q(n2643)
         );
  DFFR_X1 \id_ex/busA_q_reg[13]  ( .D(n6687), .CK(clk), .RN(n3278), .Q(n2642)
         );
  DFFR_X1 \id_ex/busA_q_reg[14]  ( .D(n6686), .CK(clk), .RN(n3277), .Q(n2641)
         );
  DFFR_X1 \id_ex/busA_q_reg[15]  ( .D(n6685), .CK(clk), .RN(n3278), .Q(n2808), 
        .QN(n6586) );
  DFFR_X1 \id_ex/busA_q_reg[16]  ( .D(n6684), .CK(clk), .RN(n3277), .Q(n2599)
         );
  DFFR_X1 \id_ex/busA_q_reg[17]  ( .D(n6683), .CK(clk), .RN(n3278), .Q(n2792), 
        .QN(n6585) );
  DFFR_X1 \id_ex/busA_q_reg[18]  ( .D(n6682), .CK(clk), .RN(n3277), .Q(n2807), 
        .QN(n6584) );
  DFFR_X1 \id_ex/busA_q_reg[19]  ( .D(n6681), .CK(clk), .RN(n3279), .Q(n2806), 
        .QN(n6583) );
  DFFR_X1 \id_ex/busA_q_reg[20]  ( .D(n6680), .CK(clk), .RN(n3279), .Q(n2805), 
        .QN(n6582) );
  DFFR_X1 \id_ex/busA_q_reg[21]  ( .D(n6679), .CK(clk), .RN(n3277), .Q(n2804), 
        .QN(n6581) );
  DFFR_X1 \id_ex/busA_q_reg[22]  ( .D(n6678), .CK(clk), .RN(n3279), .Q(n2803), 
        .QN(n6580) );
  DFFR_X1 \id_ex/busA_q_reg[23]  ( .D(n6677), .CK(clk), .RN(n3277), .Q(n2802), 
        .QN(n6579) );
  DFFR_X1 \id_ex/busA_q_reg[24]  ( .D(n6676), .CK(clk), .RN(n3279), .Q(n2801), 
        .QN(n6578) );
  DFFR_X1 \id_ex/busA_q_reg[25]  ( .D(n6675), .CK(clk), .RN(n3277), .Q(n2800), 
        .QN(n6577) );
  DFFR_X1 \id_ex/busA_q_reg[26]  ( .D(n6674), .CK(clk), .RN(n3279), .Q(n2799), 
        .QN(n6576) );
  DFFR_X1 \id_ex/busA_q_reg[27]  ( .D(n6673), .CK(clk), .RN(n3277), .Q(n2676), 
        .QN(n6575) );
  DFFR_X1 \id_ex/busA_q_reg[28]  ( .D(n6672), .CK(clk), .RN(n3279), .Q(n2675), 
        .QN(n6574) );
  DFFR_X1 \id_ex/busA_q_reg[29]  ( .D(n6671), .CK(clk), .RN(n3277), .Q(n2674), 
        .QN(n6573) );
  DFFR_X1 \id_ex/busA_q_reg[30]  ( .D(n6670), .CK(clk), .RN(n3277), .Q(n2640)
         );
  DFFR_X1 \id_ex/busA_q_reg[31]  ( .D(n6669), .CK(clk), .RN(n3272), .Q(n2639)
         );
  DFFR_X1 \id_ex/busB_q_reg[0]  ( .D(n6732), .CK(clk), .RN(n3271), .Q(n2652)
         );
  DFFR_X1 \id_ex/busB_q_reg[1]  ( .D(n6731), .CK(clk), .RN(n3276), .Q(n2660)
         );
  DFFR_X1 \id_ex/busB_q_reg[2]  ( .D(n6730), .CK(clk), .RN(n3270), .Q(n2659)
         );
  DFFR_X1 \id_ex/busB_q_reg[3]  ( .D(n6729), .CK(clk), .RN(n3275), .Q(n2658)
         );
  DFFR_X1 \id_ex/busB_q_reg[4]  ( .D(n6728), .CK(clk), .RN(n3270), .Q(n2657)
         );
  DFFR_X1 \id_ex/busB_q_reg[5]  ( .D(n6727), .CK(clk), .RN(n3275), .Q(n2672), 
        .QN(n6555) );
  DFFR_X1 \id_ex/busB_q_reg[6]  ( .D(n6726), .CK(clk), .RN(n3270), .Q(n2656)
         );
  DFFR_X1 \id_ex/busB_q_reg[7]  ( .D(n6725), .CK(clk), .RN(n3275), .Q(n2655)
         );
  DFFR_X1 \id_ex/busB_q_reg[8]  ( .D(n6724), .CK(clk), .RN(n3270), .Q(n2638)
         );
  DFFR_X1 \id_ex/busB_q_reg[9]  ( .D(n6723), .CK(clk), .RN(n3275), .Q(n2677), 
        .QN(n6554) );
  DFFR_X1 \id_ex/busB_q_reg[10]  ( .D(n6722), .CK(clk), .RN(n3276), .Q(n2634)
         );
  DFFR_X1 \id_ex/busB_q_reg[11]  ( .D(n6721), .CK(clk), .RN(n3271), .QN(n6566)
         );
  DFFR_X1 \id_ex/busB_q_reg[12]  ( .D(n6720), .CK(clk), .RN(n3276), .Q(n2654)
         );
  DFFR_X1 \id_ex/busB_q_reg[13]  ( .D(n6719), .CK(clk), .RN(n3271), .Q(n2637)
         );
  DFFR_X1 \id_ex/busB_q_reg[14]  ( .D(n6718), .CK(clk), .RN(n3276), .QN(n6565)
         );
  DFFR_X1 \id_ex/busB_q_reg[15]  ( .D(n6717), .CK(clk), .RN(n3271), .Q(n2653)
         );
  DFFR_X1 \id_ex/busB_q_reg[16]  ( .D(n6716), .CK(clk), .RN(n3276), .Q(n2813), 
        .QN(n6564) );
  DFFR_X1 \id_ex/busB_q_reg[17]  ( .D(n6715), .CK(clk), .RN(n3271), .Q(n2651)
         );
  DFFR_X1 \id_ex/busB_q_reg[18]  ( .D(n6714), .CK(clk), .RN(n3276), .Q(n2606)
         );
  DFFR_X1 \id_ex/busB_q_reg[19]  ( .D(n6713), .CK(clk), .RN(n3271), .Q(n2820), 
        .QN(n6563) );
  DFFR_X1 \id_ex/busB_q_reg[20]  ( .D(n6712), .CK(clk), .RN(n3271), .Q(n2819), 
        .QN(n6562) );
  DFFR_X1 \id_ex/busB_q_reg[21]  ( .D(n6711), .CK(clk), .RN(n3276), .Q(n2814), 
        .QN(n6561) );
  DFFR_X1 \id_ex/busB_q_reg[22]  ( .D(n6710), .CK(clk), .RN(n3271), .Q(n2818), 
        .QN(n6560) );
  DFFR_X1 \id_ex/busB_q_reg[23]  ( .D(n6709), .CK(clk), .RN(n3276), .Q(n2610)
         );
  DFFR_X1 \id_ex/busB_q_reg[24]  ( .D(n6708), .CK(clk), .RN(n3271), .Q(n2607)
         );
  DFFR_X1 \id_ex/busB_q_reg[25]  ( .D(n6707), .CK(clk), .RN(n3276), .Q(n2817), 
        .QN(n6559) );
  DFFR_X1 \id_ex/busB_q_reg[26]  ( .D(n6706), .CK(clk), .RN(n3271), .Q(n2609)
         );
  DFFR_X1 \id_ex/busB_q_reg[27]  ( .D(n6705), .CK(clk), .RN(n3275), .Q(n2608)
         );
  DFFR_X1 \id_ex/busB_q_reg[28]  ( .D(n6704), .CK(clk), .RN(n3271), .Q(n2816), 
        .QN(n6558) );
  DFFR_X1 \id_ex/busB_q_reg[29]  ( .D(n6703), .CK(clk), .RN(n3275), .Q(n2815), 
        .QN(n6557) );
  DFFR_X1 \id_ex/busB_q_reg[30]  ( .D(n6702), .CK(clk), .RN(n3275), .Q(n2812), 
        .QN(n6556) );
  DFFR_X1 \id_ex/busB_q_reg[31]  ( .D(n6701), .CK(clk), .RN(n3270), .Q(n3021)
         );
  DFFR_X1 \id_ex/aluCtrl_q_reg[0]  ( .D(n2018), .CK(clk), .RN(n3278), .Q(n2787), .QN(n6617) );
  DFFR_X1 \id_ex/aluCtrl_q_reg[2]  ( .D(n2016), .CK(clk), .RN(n3278), .Q(n2663), .QN(n6600) );
  DFFR_X1 \if_id/incPC_q_reg[0]  ( .D(n6753), .CK(clk), .RN(n3268), .Q(n2619)
         );
  DFFR_X1 \id_ex/incPC_q_reg[0]  ( .D(n6764), .CK(clk), .RN(n3273), .Q(n2736), 
        .QN(n6596) );
  DFFR_X1 \if_id/incPC_q_reg[1]  ( .D(n6752), .CK(clk), .RN(n3254), .Q(n2618)
         );
  DFFR_X1 \id_ex/incPC_q_reg[1]  ( .D(n6763), .CK(clk), .RN(n3269), .Q(n2735), 
        .QN(n6595) );
  DFFR_X1 \if_id/incPC_q_reg[2]  ( .D(n1981), .CK(clk), .RN(n3267), .Q(n2930)
         );
  DFFR_X1 \id_ex/incPC_q_reg[2]  ( .D(n1980), .CK(clk), .RN(n3272), .Q(n2734), 
        .QN(n6521) );
  DFFR_X1 \if_id/incPC_q_reg[3]  ( .D(n1977), .CK(clk), .RN(n3254), .Q(n2617)
         );
  DFFR_X1 \id_ex/incPC_q_reg[3]  ( .D(n1976), .CK(clk), .RN(n3269), .Q(n2733), 
        .QN(n6520) );
  DFFR_X1 \if_id/incPC_q_reg[4]  ( .D(n1973), .CK(clk), .RN(n3267), .Q(n2616)
         );
  DFFR_X1 \id_ex/incPC_q_reg[4]  ( .D(n1972), .CK(clk), .RN(n3272), .Q(n2732), 
        .QN(n6519) );
  DFFR_X1 \if_id/incPC_q_reg[6]  ( .D(n1969), .CK(clk), .RN(n3267), .Q(n2615)
         );
  DFFR_X1 \id_ex/incPC_q_reg[6]  ( .D(n1968), .CK(clk), .RN(n3272), .Q(n2731), 
        .QN(n6518) );
  DFFR_X1 \if_id/incPC_q_reg[7]  ( .D(n1966), .CK(clk), .RN(n3254), .Q(n2614)
         );
  DFFR_X1 \id_ex/incPC_q_reg[7]  ( .D(n1965), .CK(clk), .RN(n3268), .Q(n2730), 
        .QN(n6517) );
  DFFR_X1 \if_id/incPC_q_reg[8]  ( .D(n1963), .CK(clk), .RN(n3267), .Q(n2613)
         );
  DFFR_X1 \id_ex/incPC_q_reg[8]  ( .D(n1962), .CK(clk), .RN(n3272), .Q(n2729), 
        .QN(n6516) );
  DFFR_X1 \if_id/incPC_q_reg[9]  ( .D(n1960), .CK(clk), .RN(n3254), .Q(n2612)
         );
  DFFR_X1 \id_ex/incPC_q_reg[9]  ( .D(n1959), .CK(clk), .RN(n3268), .Q(n2728), 
        .QN(n6515) );
  DFFR_X1 \if_id/incPC_q_reg[12]  ( .D(n1957), .CK(clk), .RN(n3255), .Q(n2983), 
        .QN(n6514) );
  DFFR_X1 \id_ex/incPC_q_reg[12]  ( .D(n1956), .CK(clk), .RN(n3269), .Q(n2727), 
        .QN(n6513) );
  DFFR_X1 \if_id/incPC_q_reg[5]  ( .D(n1946), .CK(clk), .RN(n3254), .Q(n2611)
         );
  DFFR_X1 \id_ex/incPC_q_reg[5]  ( .D(n1945), .CK(clk), .RN(n3268), .Q(n2726), 
        .QN(n6512) );
  DFFR_X1 \if_id/incPC_q_reg[31]  ( .D(n1917), .CK(clk), .RN(n3267), .Q(n2929)
         );
  DFFR_X1 \id_ex/incPC_q_reg[31]  ( .D(n1916), .CK(clk), .RN(n3272), .Q(n2725), 
        .QN(n6510) );
  DFFS_X2 \id_ex/instr_q_reg[4]  ( .D(n6774), .CK(clk), .SN(n3280), .Q(
        instr_2[4]) );
  DFFS_X2 \id_ex/instr_q_reg[2]  ( .D(n6776), .CK(clk), .SN(n3280), .Q(
        instr_2[2]) );
  DFFS_X2 \id_ex/not_trap_q_reg  ( .D(n3042), .CK(clk), .SN(n3280), .QN(n6341)
         );
  DFFS_X2 \ex_mem/not_trap_q_reg  ( .D(\ex_mem/N242 ), .CK(clk), .SN(n3280), 
        .Q(not_trap_3) );
  DFFS_X2 \id_ex/instr_q_reg[0]  ( .D(\id_ex/N4 ), .CK(clk), .SN(n3279), .Q(
        instr_2[0]) );
  DFF_X2 \mem_wb/memRdData_q_reg[0]  ( .D(n2267), .CK(clk), .Q(
        \wb/dsize_reg/z2 [0]), .QN(n2695) );
  DFF_X2 \mem_wb/memRdData_q_reg[1]  ( .D(n2266), .CK(clk), .Q(
        \wb/dsize_reg/z2 [1]), .QN(n2828) );
  DFF_X2 \mem_wb/memRdData_q_reg[2]  ( .D(n2265), .CK(clk), .Q(
        \wb/dsize_reg/z2 [2]), .QN(n2830) );
  DFF_X2 \mem_wb/memRdData_q_reg[3]  ( .D(n2264), .CK(clk), .Q(
        \wb/dsize_reg/z2 [3]), .QN(n2992) );
  DFF_X2 \mem_wb/memRdData_q_reg[4]  ( .D(n2263), .CK(clk), .Q(
        \wb/dsize_reg/z2 [4]), .QN(n2705) );
  DFF_X2 \mem_wb/memRdData_q_reg[5]  ( .D(n2262), .CK(clk), .Q(
        \wb/dsize_reg/z2 [5]), .QN(n2694) );
  DFF_X2 \mem_wb/memRdData_q_reg[6]  ( .D(n2261), .CK(clk), .Q(
        \wb/dsize_reg/z2 [6]), .QN(n2693) );
  DFF_X2 \mem_wb/memRdData_q_reg[7]  ( .D(n2260), .CK(clk), .Q(
        \wb/dsize_reg/z2 [7]), .QN(n2704) );
  DFF_X2 \mem_wb/memRdData_q_reg[8]  ( .D(n2259), .CK(clk), .Q(
        \wb/dsize_reg/z2 [8]), .QN(n2702) );
  DFF_X2 \mem_wb/memRdData_q_reg[9]  ( .D(n2258), .CK(clk), .Q(
        \wb/dsize_reg/z2 [9]), .QN(n2898) );
  DFF_X2 \mem_wb/memRdData_q_reg[10]  ( .D(n2257), .CK(clk), .Q(
        \wb/dsize_reg/z2 [10]), .QN(n2959) );
  DFF_X2 \mem_wb/memRdData_q_reg[11]  ( .D(n2256), .CK(clk), .Q(
        \wb/dsize_reg/z2 [11]), .QN(n2827) );
  DFF_X2 \mem_wb/memRdData_q_reg[12]  ( .D(n2255), .CK(clk), .Q(
        \wb/dsize_reg/z2 [12]), .QN(n3086) );
  DFF_X2 \mem_wb/memRdData_q_reg[13]  ( .D(n2254), .CK(clk), .Q(
        \wb/dsize_reg/z2 [13]), .QN(n2829) );
  DFF_X2 \mem_wb/memRdData_q_reg[14]  ( .D(n2253), .CK(clk), .Q(
        \wb/dsize_reg/z2 [14]), .QN(n2892) );
  DFF_X2 \mem_wb/memRdData_q_reg[15]  ( .D(n2252), .CK(clk), .Q(
        \wb/dsize_reg/z2 [15]), .QN(n2893) );
  DFF_X2 \mem_wb/memRdData_q_reg[16]  ( .D(n2251), .CK(clk), .Q(
        \wb/dsize_reg/z2 [16]), .QN(n2668) );
  DFF_X2 \mem_wb/memRdData_q_reg[17]  ( .D(n2250), .CK(clk), .Q(
        \wb/dsize_reg/z2 [17]), .QN(n2670) );
  DFF_X2 \mem_wb/memRdData_q_reg[18]  ( .D(n2249), .CK(clk), .Q(
        \wb/dsize_reg/z2 [18]), .QN(n2701) );
  DFF_X2 \mem_wb/memRdData_q_reg[19]  ( .D(n2248), .CK(clk), .Q(
        \wb/dsize_reg/z2 [19]), .QN(n3124) );
  DFF_X2 \mem_wb/memRdData_q_reg[20]  ( .D(n2247), .CK(clk), .Q(
        \wb/dsize_reg/z2 [20]), .QN(n2699) );
  DFF_X2 \mem_wb/memRdData_q_reg[21]  ( .D(n2246), .CK(clk), .Q(
        \wb/dsize_reg/z2 [21]), .QN(n2719) );
  DFF_X2 \mem_wb/memRdData_q_reg[22]  ( .D(n2245), .CK(clk), .Q(
        \wb/dsize_reg/z2 [22]), .QN(n2687) );
  DFF_X2 \mem_wb/memRdData_q_reg[23]  ( .D(n2244), .CK(clk), .Q(
        \wb/dsize_reg/z2 [23]), .QN(n2707) );
  DFF_X2 \mem_wb/memRdData_q_reg[24]  ( .D(n2243), .CK(clk), .Q(
        \wb/dsize_reg/z2 [24]), .QN(n2667) );
  DFF_X2 \mem_wb/memRdData_q_reg[25]  ( .D(n2242), .CK(clk), .Q(
        \wb/dsize_reg/z2 [25]), .QN(n2703) );
  DFF_X2 \mem_wb/memRdData_q_reg[26]  ( .D(n2241), .CK(clk), .Q(
        \wb/dsize_reg/z2 [26]), .QN(n2665) );
  DFF_X2 \mem_wb/memRdData_q_reg[27]  ( .D(n2240), .CK(clk), .Q(
        \wb/dsize_reg/z2 [27]), .QN(n2666) );
  DFF_X2 \mem_wb/memRdData_q_reg[28]  ( .D(n2239), .CK(clk), .Q(
        \wb/dsize_reg/z2 [28]), .QN(n2686) );
  DFF_X2 \mem_wb/memRdData_q_reg[29]  ( .D(n2238), .CK(clk), .Q(
        \wb/dsize_reg/z2 [29]), .QN(n2673) );
  DFF_X2 \mem_wb/memRdData_q_reg[30]  ( .D(n2237), .CK(clk), .Q(
        \wb/dsize_reg/z2 [30]), .QN(n2783) );
  DFF_X2 \mem_wb/memRdData_q_reg[31]  ( .D(n2236), .CK(clk), .Q(
        \wb/dsize_reg/z2 [31]), .QN(n2845) );
  DFF_X2 \mem_wb/aluRes_q_reg[0]  ( .D(n2235), .CK(clk), .QN(n6340) );
  DFF_X2 \mem_wb/aluRes_q_reg[16]  ( .D(n6662), .CK(clk), .Q(n2850), .QN(n6339) );
  DFF_X2 \mem_wb/aluRes_q_reg[21]  ( .D(n6657), .CK(clk), .QN(n6338) );
  DFF_X2 \mem_wb/aluRes_q_reg[22]  ( .D(n6656), .CK(clk), .QN(n6337) );
  DFF_X2 \mem_wb/aluRes_q_reg[23]  ( .D(n6655), .CK(clk), .QN(n6336) );
  DFF_X2 \mem_wb/aluRes_q_reg[24]  ( .D(n6654), .CK(clk), .QN(n6335) );
  DFF_X2 \mem_wb/aluRes_q_reg[25]  ( .D(n6653), .CK(clk), .QN(n6334) );
  DFF_X2 \mem_wb/aluRes_q_reg[31]  ( .D(n6647), .CK(clk), .Q(n2950), .QN(n6333) );
  DFF_X2 \mem_wb/aluRes_q_reg[4]  ( .D(n2227), .CK(clk), .QN(n6332) );
  DFF_X2 \mem_wb/aluRes_q_reg[9]  ( .D(n6645), .CK(clk), .Q(n3024), .QN(n6331)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[2]  ( .D(n2225), .CK(clk), .QN(n6330) );
  DFF_X2 \mem_wb/aluRes_q_reg[1]  ( .D(n2224), .CK(clk), .QN(n6329) );
  DFF_X2 \mem_wb/aluRes_q_reg[3]  ( .D(n2223), .CK(clk), .QN(n6328) );
  DFF_X2 \mem_wb/aluRes_q_reg[6]  ( .D(n2222), .CK(clk), .QN(n6327) );
  DFF_X2 \mem_wb/aluRes_q_reg[11]  ( .D(n6667), .CK(clk), .Q(n2811), .QN(n6326) );
  DFF_X2 \mem_wb/aluRes_q_reg[7]  ( .D(n2220), .CK(clk), .Q(n3031), .QN(n6325)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[29]  ( .D(n6649), .CK(clk), .QN(n6324) );
  DFF_X2 \mem_wb/aluRes_q_reg[8]  ( .D(n6646), .CK(clk), .Q(n3025), .QN(n6323)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[12]  ( .D(n6666), .CK(clk), .Q(n3026), .QN(n6322) );
  DFF_X2 \mem_wb/aluRes_q_reg[13]  ( .D(n6665), .CK(clk), .Q(n2848), .QN(n6321) );
  DFF_X2 \mem_wb/aluRes_q_reg[10]  ( .D(n6668), .CK(clk), .Q(n2989), .QN(n6320) );
  DFF_X2 \mem_wb/reg31Val_q_reg[30]  ( .D(n2174), .CK(clk), .Q(reg31Val_0[30]), 
        .QN(n2980) );
  DFF_X2 \mem_wb/aluRes_q_reg[30]  ( .D(n6648), .CK(clk), .Q(n2995), .QN(n6319) );
  DFF_X2 \mem_wb/aluRes_q_reg[19]  ( .D(n6659), .CK(clk), .Q(n2991), .QN(n6318) );
  DFFS_X2 \if_id/instr_q_reg[4]  ( .D(n2143), .CK(clk), .SN(n3279), .Q(n2712), 
        .QN(n6317) );
  DFFS_X2 \if_id/instr_q_reg[2]  ( .D(n2141), .CK(clk), .SN(n3279), .Q(n2871), 
        .QN(n6316) );
  DFFS_X2 \if_id/instr_q_reg[0]  ( .D(n2139), .CK(clk), .SN(n3279), .Q(n2837), 
        .QN(n6315) );
  DFF_X2 \mem_wb/fp_q_reg  ( .D(n2128), .CK(clk), .Q(n3084), .QN(n6314) );
  DFF_X2 \ex_mem/dSize_q_reg[0]  ( .D(n2125), .CK(clk), .Q(dSize[0]) );
  DFF_X2 \mem_wb/dSize_q_reg[0]  ( .D(n2124), .CK(clk), .QN(n6313) );
  DFF_X2 \ex_mem/dSize_q_reg[1]  ( .D(n2122), .CK(clk), .Q(dSize[1]) );
  DFF_X2 \mem_wb/dSize_q_reg[1]  ( .D(n2121), .CK(clk), .Q(n2722), .QN(n6312)
         );
  DFF_X2 \mem_wb/rd_q_reg[1]  ( .D(n6642), .CK(clk), .Q(rd[1]) );
  DFF_X2 \mem_wb/rd_q_reg[2]  ( .D(n6641), .CK(clk), .Q(rd[2]) );
  DFFRS_X2 \ifetch/dffa/q_reg[30]  ( .D(n2015), .CK(clk), .RN(n1914), .SN(
        n1913), .Q(n2961) );
  DFFRS_X2 \ifetch/dffa/q_reg[29]  ( .D(n2014), .CK(clk), .RN(n1912), .SN(
        n1911), .Q(n2971) );
  DFFRS_X2 \ifetch/dffa/q_reg[28]  ( .D(n2013), .CK(clk), .RN(n1910), .SN(
        n1909), .Q(n2970) );
  DFFRS_X2 \ifetch/dffa/q_reg[27]  ( .D(n2012), .CK(clk), .RN(n1908), .SN(
        n1907), .Q(n2969) );
  DFFRS_X2 \ifetch/dffa/q_reg[26]  ( .D(n2011), .CK(clk), .RN(n1906), .SN(
        n1905), .Q(n2968) );
  DFFRS_X2 \ifetch/dffa/q_reg[25]  ( .D(n2010), .CK(clk), .RN(n1904), .SN(
        n1903), .Q(n2967) );
  DFFRS_X2 \ifetch/dffa/q_reg[24]  ( .D(n2009), .CK(clk), .RN(n1902), .SN(
        n1901), .Q(n2966) );
  DFFRS_X2 \ifetch/dffa/q_reg[23]  ( .D(n2008), .CK(clk), .RN(n1900), .SN(
        n1899), .Q(n2965) );
  DFFRS_X2 \ifetch/dffa/q_reg[22]  ( .D(n2007), .CK(clk), .RN(n1898), .SN(
        n1897), .Q(n2964) );
  DFFRS_X2 \ifetch/dffa/q_reg[21]  ( .D(n2006), .CK(clk), .RN(n1896), .SN(
        n1895), .Q(n2963) );
  DFFRS_X2 \ifetch/dffa/q_reg[20]  ( .D(n2005), .CK(clk), .RN(n1894), .SN(
        n1893), .Q(n2775) );
  DFFRS_X2 \ifetch/dffa/q_reg[19]  ( .D(n2004), .CK(clk), .RN(n1892), .SN(
        n1891), .Q(n2774) );
  DFFRS_X2 \ifetch/dffa/q_reg[18]  ( .D(n2003), .CK(clk), .RN(n1890), .SN(
        n1889), .Q(n2773) );
  DFFRS_X2 \ifetch/dffa/q_reg[17]  ( .D(n2002), .CK(clk), .RN(n1888), .SN(
        n1887), .Q(n2772) );
  DFFRS_X2 \ifetch/dffa/q_reg[16]  ( .D(n2001), .CK(clk), .RN(n1886), .SN(
        n1885), .Q(n2771) );
  DFFRS_X2 \ifetch/dffa/q_reg[15]  ( .D(n2000), .CK(clk), .RN(n1884), .SN(
        n1883), .Q(n2770) );
  DFFRS_X2 \ifetch/dffa/q_reg[14]  ( .D(n1999), .CK(clk), .RN(n1882), .SN(
        n1881), .Q(n2769) );
  DFFRS_X2 \ifetch/dffa/q_reg[13]  ( .D(n1998), .CK(clk), .RN(n1880), .SN(
        n1879), .Q(n2768) );
  DFFRS_X2 \ifetch/dffa/q_reg[11]  ( .D(n1997), .CK(clk), .RN(n1878), .SN(
        n1877), .Q(n2767) );
  DFFRS_X2 \ifetch/dffa/q_reg[10]  ( .D(n1996), .CK(clk), .RN(n1876), .SN(
        n1875), .Q(n2766) );
  DFF_X2 \mem_wb/rd_q_reg[0]  ( .D(n6643), .CK(clk), .Q(rd[0]) );
  DFF_X2 \mem_wb/rd_q_reg[4]  ( .D(n6639), .CK(clk), .Q(rd[4]) );
  DFF_X2 \mem_wb/rd_q_reg[3]  ( .D(n6640), .CK(clk), .Q(rd[3]) );
  DFF_X2 \mem_wb/link_q_reg  ( .D(n1992), .CK(clk), .Q(n3119), .QN(n6311) );
  DFF_X2 \mem_wb/memRd_q_reg  ( .D(n6644), .CK(clk), .Q(n3118), .QN(n6310) );
  DFFRS_X2 \ifetch/dffa/q_reg[0]  ( .D(n1990), .CK(clk), .RN(n1874), .SN(n1873), .QN(n6523) );
  DFF_X2 \mem_wb/reg31Val_q_reg[0]  ( .D(n6638), .CK(clk), .Q(reg31Val_0[0]), 
        .QN(n3032) );
  DFFRS_X2 \ifetch/dffa/q_reg[1]  ( .D(n1986), .CK(clk), .RN(n1872), .SN(n1871), .QN(n6522) );
  DFF_X2 \mem_wb/reg31Val_q_reg[1]  ( .D(n6637), .CK(clk), .Q(reg31Val_0[1])
         );
  DFFRS_X2 \ifetch/dffa/q_reg[2]  ( .D(n6756), .CK(clk), .RN(n1870), .SN(n1869), .Q(n2765) );
  DFF_X2 \mem_wb/reg31Val_q_reg[2]  ( .D(n1979), .CK(clk), .Q(reg31Val_0[2])
         );
  DFFRS_X2 \ifetch/dffa/q_reg[3]  ( .D(n1978), .CK(clk), .RN(n1868), .SN(n1867), .Q(n3035) );
  DFF_X2 \mem_wb/reg31Val_q_reg[3]  ( .D(n1975), .CK(clk), .Q(reg31Val_0[3]), 
        .QN(n3022) );
  DFFRS_X2 \ifetch/dffa/q_reg[4]  ( .D(n1974), .CK(clk), .RN(n1866), .SN(n1865), .Q(n3034) );
  DFF_X2 \mem_wb/reg31Val_q_reg[4]  ( .D(n1971), .CK(clk), .Q(reg31Val_0[4])
         );
  DFFRS_X2 \ifetch/dffa/q_reg[6]  ( .D(n1970), .CK(clk), .RN(n1864), .SN(n1863), .Q(n3036) );
  DFFRS_X2 \ifetch/dffa/q_reg[7]  ( .D(n1967), .CK(clk), .RN(n1862), .SN(n1861), .Q(n3039) );
  DFFRS_X2 \ifetch/dffa/q_reg[8]  ( .D(n1964), .CK(clk), .RN(n1860), .SN(n1859), .Q(n3038) );
  DFFRS_X2 \ifetch/dffa/q_reg[9]  ( .D(n1961), .CK(clk), .RN(n1858), .SN(n1857), .Q(n3040) );
  DFFRS_X2 \ifetch/dffa/q_reg[12]  ( .D(n1958), .CK(clk), .RN(n1856), .SN(
        n1855), .Q(n2962) );
  DFF_X2 \mem_wb/reg31Val_q_reg[29]  ( .D(n1955), .CK(clk), .Q(reg31Val_0[29]), 
        .QN(n2986) );
  DFF_X2 \mem_wb/reg31Val_q_reg[28]  ( .D(n1954), .CK(clk), .Q(reg31Val_0[28]), 
        .QN(n3023) );
  DFF_X2 \mem_wb/aluRes_q_reg[28]  ( .D(n6650), .CK(clk), .Q(n2996), .QN(n6309) );
  DFF_X2 \mem_wb/reg31Val_q_reg[27]  ( .D(n1952), .CK(clk), .Q(reg31Val_0[27]), 
        .QN(n2977) );
  DFF_X2 \mem_wb/aluRes_q_reg[27]  ( .D(n6651), .CK(clk), .QN(n6308) );
  DFF_X2 \mem_wb/reg31Val_q_reg[26]  ( .D(n1950), .CK(clk), .Q(reg31Val_0[26]), 
        .QN(n2976) );
  DFF_X2 \mem_wb/aluRes_q_reg[26]  ( .D(n6652), .CK(clk), .QN(n6307) );
  DFF_X2 \mem_wb/aluRes_q_reg[5]  ( .D(n1948), .CK(clk), .Q(n3125), .QN(n6306)
         );
  DFFRS_X2 \ifetch/dffa/q_reg[5]  ( .D(n1947), .CK(clk), .RN(n1854), .SN(n1853), .Q(n3037) );
  DFF_X2 \mem_wb/reg31Val_q_reg[6]  ( .D(n1944), .CK(clk), .Q(reg31Val_0[6])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[5]  ( .D(n1943), .CK(clk), .Q(reg31Val_0[5])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[8]  ( .D(n1942), .CK(clk), .Q(reg31Val_0[8])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[7]  ( .D(n1941), .CK(clk), .Q(reg31Val_0[7])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[9]  ( .D(n1940), .CK(clk), .Q(reg31Val_0[9]), 
        .QN(n2889) );
  DFF_X2 \mem_wb/reg31Val_q_reg[11]  ( .D(n1939), .CK(clk), .Q(reg31Val_0[11])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[10]  ( .D(n1938), .CK(clk), .Q(reg31Val_0[10])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[25]  ( .D(n1937), .CK(clk), .Q(reg31Val_0[25]), 
        .QN(n2985) );
  DFF_X2 \mem_wb/reg31Val_q_reg[24]  ( .D(n1936), .CK(clk), .Q(reg31Val_0[24]), 
        .QN(n2979) );
  DFF_X2 \mem_wb/reg31Val_q_reg[23]  ( .D(n1935), .CK(clk), .Q(reg31Val_0[23]), 
        .QN(n2978) );
  DFF_X2 \mem_wb/reg31Val_q_reg[22]  ( .D(n1934), .CK(clk), .Q(reg31Val_0[22]), 
        .QN(n2928) );
  DFF_X2 \mem_wb/reg31Val_q_reg[21]  ( .D(n1933), .CK(clk), .Q(reg31Val_0[21]), 
        .QN(n2987) );
  DFF_X2 \mem_wb/reg31Val_q_reg[20]  ( .D(n1932), .CK(clk), .Q(reg31Val_0[20]), 
        .QN(n2927) );
  DFF_X2 \mem_wb/reg31Val_q_reg[19]  ( .D(n1931), .CK(clk), .Q(reg31Val_0[19]), 
        .QN(n2988) );
  DFF_X2 \mem_wb/reg31Val_q_reg[18]  ( .D(n1930), .CK(clk), .Q(reg31Val_0[18]), 
        .QN(n2922) );
  DFF_X2 \mem_wb/reg31Val_q_reg[17]  ( .D(n1929), .CK(clk), .Q(reg31Val_0[17]), 
        .QN(n2874) );
  DFF_X2 \mem_wb/reg31Val_q_reg[16]  ( .D(n1928), .CK(clk), .Q(reg31Val_0[16])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[15]  ( .D(n1927), .CK(clk), .Q(reg31Val_0[15]), 
        .QN(n2925) );
  DFF_X2 \mem_wb/reg31Val_q_reg[14]  ( .D(n1926), .CK(clk), .Q(reg31Val_0[14]), 
        .QN(n2982) );
  DFF_X2 \mem_wb/aluRes_q_reg[14]  ( .D(n6664), .CK(clk), .QN(n6305) );
  DFF_X2 \mem_wb/aluRes_q_reg[20]  ( .D(n6658), .CK(clk), .QN(n6304) );
  DFF_X2 \mem_wb/aluRes_q_reg[15]  ( .D(n6663), .CK(clk), .Q(n3027), .QN(n6303) );
  DFF_X2 \mem_wb/aluRes_q_reg[18]  ( .D(n6660), .CK(clk), .QN(n6302) );
  DFF_X2 \mem_wb/aluRes_q_reg[17]  ( .D(n6661), .CK(clk), .QN(n6301) );
  DFF_X2 \mem_wb/reg31Val_q_reg[13]  ( .D(n1920), .CK(clk), .Q(reg31Val_0[13]), 
        .QN(n2882) );
  DFF_X2 \mem_wb/reg31Val_q_reg[12]  ( .D(n1919), .CK(clk), .Q(reg31Val_0[12]), 
        .QN(n2924) );
  DFFRS_X2 \ifetch/dffa/q_reg[31]  ( .D(n1918), .CK(clk), .RN(n1852), .SN(
        n1851), .Q(n3029), .QN(n6511) );
  DFFR_X2 \id_ex/busB_sel_q_reg[1]  ( .D(\id_ex/N41 ), .CK(clk), .RN(n3254), 
        .QN(n6232) );
  DFFR_X2 \id_ex/busB_sel_q_reg[0]  ( .D(\id_ex/N40 ), .CK(clk), .RN(n3255), 
        .Q(n3122), .QN(n6237) );
  DFFR_X2 \ex_mem/imm32_q_reg[10]  ( .D(\ex_mem/N141 ), .CK(clk), .RN(n3262), 
        .QN(n6202) );
  DFFR_X2 \ex_mem/incPC_q_reg[10]  ( .D(\ex_mem/N45 ), .CK(clk), .RN(n3250), 
        .Q(n2856), .QN(n6279) );
  DFFR_X2 \ex_mem/incPC_q_reg[4]  ( .D(\ex_mem/N39 ), .CK(clk), .RN(n3260), 
        .Q(n2852), .QN(n6188) );
  DFFR_X2 \ex_mem/incPC_q_reg[3]  ( .D(\ex_mem/N38 ), .CK(clk), .RN(n3260), 
        .Q(n2710), .QN(n6189) );
  DFFR_X2 \if_id/instr_q_reg[27]  ( .D(n2166), .CK(clk), .RN(n3253), .Q(n2594), 
        .QN(n6589) );
  DFFR_X2 \id_ex/aluCtrl_q_reg[1]  ( .D(n2017), .CK(clk), .RN(n3278), .Q(n2602), .QN(n6603) );
  DFFR_X2 \ex_mem/incPC_q_reg[2]  ( .D(\ex_mem/N37 ), .CK(clk), .RN(n3261), 
        .QN(n6190) );
  DFFR_X2 \ex_mem/incPC_q_reg[11]  ( .D(\ex_mem/N46 ), .CK(clk), .RN(n3250), 
        .Q(n2631), .QN(n6278) );
  DFFR_X2 \ex_mem/imm32_q_reg[11]  ( .D(\ex_mem/N142 ), .CK(clk), .RN(n3262), 
        .Q(n2896), .QN(n6203) );
  DFFR_X2 \mem_wb/regWr_q_reg  ( .D(\mem_wb/N36 ), .CK(clk), .RN(n3265), .Q(
        regWr), .QN(n3139) );
  DFFR_X2 \ex_mem/incPC_q_reg[0]  ( .D(\ex_mem/N35 ), .CK(clk), .RN(n3261), 
        .Q(reg31Val_3[0]) );
  DFFR_X2 \ex_mem/incPC_q_reg[1]  ( .D(\ex_mem/N36 ), .CK(clk), .RN(n3261), 
        .Q(reg31Val_3[1]) );
  DFFR_X2 \ex_mem/incPC_q_reg[6]  ( .D(\ex_mem/N41 ), .CK(clk), .RN(n3260), 
        .Q(n2671), .QN(n6187) );
  DFFR_X2 \ex_mem/incPC_q_reg[5]  ( .D(\ex_mem/N40 ), .CK(clk), .RN(n3259), 
        .Q(n2669), .QN(n6177) );
  DFFR_X2 \ex_mem/incPC_q_reg[16]  ( .D(\ex_mem/N51 ), .CK(clk), .RN(n3250), 
        .QN(n6274) );
  DFFR_X2 \ex_mem/incPC_q_reg[17]  ( .D(\ex_mem/N52 ), .CK(clk), .RN(n3250), 
        .Q(n2700), .QN(n6273) );
  DFFR_X2 \ex_mem/imm32_q_reg[17]  ( .D(\ex_mem/N148 ), .CK(clk), .RN(n3262), 
        .Q(n2998), .QN(n6209) );
  DFFR_X2 \ex_mem/imm32_q_reg[16]  ( .D(\ex_mem/N147 ), .CK(clk), .RN(n3262), 
        .QN(n6208) );
  DFFR_X2 \ex_mem/aluRes_q_reg[14]  ( .D(\ex_mem/N210 ), .CK(clk), .RN(n3258), 
        .Q(memAddr[14]), .QN(n6176) );
  DFFR_X2 \id_ex/aluSrc_q_reg  ( .D(n2136), .CK(clk), .RN(n3278), .Q(n3097), 
        .QN(n6615) );
  DFFR_X2 \ex_mem/incPC_q_reg[7]  ( .D(\ex_mem/N42 ), .CK(clk), .RN(n3260), 
        .Q(n2683), .QN(n6186) );
  DFF_X1 \mem_wb/reg31Val_q_reg[31]  ( .D(n1915), .CK(clk), .Q(reg31Val_0[31])
         );
  INV_X8 U2578 ( .A(n2576), .ZN(n2577) );
  NAND3_X2 U2579 ( .A1(n3142), .A2(n3652), .A3(n3648), .ZN(n3650) );
  NAND2_X1 U2580 ( .A1(n3463), .A2(n3462), .ZN(n3468) );
  NAND3_X2 U2581 ( .A1(\wb/dsize_reg/z2 [28]), .A2(n3177), .A3(n4440), .ZN(
        n4219) );
  INV_X4 U2582 ( .A(n4073), .ZN(n4440) );
  NAND2_X2 U2583 ( .A1(n4406), .A2(n4405), .ZN(n4077) );
  XNOR2_X1 U2584 ( .A(n5638), .B(n5421), .ZN(n5986) );
  NAND3_X4 U2585 ( .A1(\wb/dsize_reg/z2 [11]), .A2(n4355), .A3(n4354), .ZN(
        n4366) );
  NAND4_X2 U2586 ( .A1(n3243), .A2(n3172), .A3(n4262), .A4(n4263), .ZN(n4271)
         );
  NAND2_X4 U2587 ( .A1(n3645), .A2(n3644), .ZN(n3652) );
  INV_X1 U2588 ( .A(n3645), .ZN(n3647) );
  XNOR2_X1 U2589 ( .A(n3752), .B(n3755), .ZN(n3754) );
  INV_X8 U2590 ( .A(n2680), .ZN(n3184) );
  OAI221_X4 U2591 ( .B1(n6567), .B2(n3155), .C1(n3185), .C2(n4466), .A(n4465), 
        .ZN(n5444) );
  NAND2_X1 U2592 ( .A1(n3789), .A2(n3784), .ZN(n3792) );
  AOI22_X1 U2593 ( .A1(n3225), .A2(n5189), .B1(n5947), .B2(n5678), .ZN(n4991)
         );
  NAND2_X4 U2594 ( .A1(n3700), .A2(n2826), .ZN(n3702) );
  INV_X8 U2595 ( .A(n3622), .ZN(n3337) );
  AOI21_X1 U2596 ( .B1(n3624), .B2(n3623), .A(n3622), .ZN(n3626) );
  NAND4_X4 U2597 ( .A1(n3681), .A2(n3680), .A3(iAddr[29]), .A4(n3813), .ZN(
        n3682) );
  INV_X16 U2598 ( .A(n3800), .ZN(n3813) );
  INV_X2 U2599 ( .A(n5172), .ZN(n4826) );
  NAND2_X4 U2600 ( .A1(n3397), .A2(n3631), .ZN(n3586) );
  INV_X4 U2601 ( .A(n4916), .ZN(n2576) );
  AOI22_X1 U2602 ( .A1(n3225), .A2(n5679), .B1(n6029), .B2(n5678), .ZN(n5683)
         );
  INV_X1 U2603 ( .A(n5679), .ZN(n5136) );
  OAI211_X4 U2604 ( .C1(n3612), .C2(n2857), .A(n3611), .B(n3610), .ZN(n3613)
         );
  NAND4_X4 U2605 ( .A1(n4437), .A2(n4436), .A3(n4435), .A4(n4460), .ZN(n3062)
         );
  INV_X2 U2606 ( .A(n5226), .ZN(n4072) );
  XNOR2_X1 U2607 ( .A(n5669), .B(n5668), .ZN(n5975) );
  NAND3_X1 U2608 ( .A1(n5333), .A2(n5330), .A3(n5668), .ZN(n4913) );
  OAI221_X1 U2609 ( .B1(n6575), .B2(n3155), .C1(n4507), .C2(n3184), .A(n4506), 
        .ZN(n5173) );
  OAI221_X1 U2610 ( .B1(n6577), .B2(n3155), .C1(n4484), .C2(n3184), .A(n4483), 
        .ZN(n5199) );
  OAI221_X1 U2611 ( .B1(n6579), .B2(n3155), .C1(n4464), .C2(n3184), .A(n4463), 
        .ZN(n5865) );
  OAI221_X1 U2612 ( .B1(n6578), .B2(n3155), .C1(n4692), .C2(n3184), .A(n4691), 
        .ZN(n5825) );
  OAI221_X1 U2613 ( .B1(n6582), .B2(n3155), .C1(n4722), .C2(n3184), .A(n4721), 
        .ZN(n5172) );
  OAI221_X1 U2614 ( .B1(n6583), .B2(n3155), .C1(n4071), .C2(n3184), .A(n4070), 
        .ZN(n5226) );
  NAND3_X1 U2615 ( .A1(n5150), .A2(n5151), .A3(n3184), .ZN(n4446) );
  NAND3_X1 U2616 ( .A1(n5143), .A2(n5142), .A3(n3184), .ZN(n4617) );
  AND3_X2 U2617 ( .A1(n4877), .A2(n4878), .A3(n3184), .ZN(n2926) );
  NAND2_X4 U2618 ( .A1(n3721), .A2(n2690), .ZN(n3717) );
  INV_X8 U2619 ( .A(n3308), .ZN(n3721) );
  NAND2_X4 U2620 ( .A1(n3708), .A2(n2689), .ZN(n3710) );
  NAND2_X1 U2621 ( .A1(n2683), .A2(n2919), .ZN(n3456) );
  NAND2_X4 U2622 ( .A1(n3307), .A2(n2683), .ZN(n3308) );
  NAND2_X2 U2623 ( .A1(op0_1), .A2(n6385), .ZN(n6492) );
  XNOR2_X1 U2624 ( .A(n3714), .B(n2631), .ZN(n3715) );
  NAND2_X4 U2625 ( .A1(n3712), .A2(n2856), .ZN(n3714) );
  INV_X2 U2626 ( .A(n6408), .ZN(n2578) );
  INV_X4 U2627 ( .A(n2578), .ZN(n2579) );
  NAND3_X4 U2628 ( .A1(n6137), .A2(n2780), .A3(n6588), .ZN(n6421) );
  INV_X4 U2629 ( .A(n3142), .ZN(n2580) );
  AOI21_X2 U2630 ( .B1(n6430), .B2(n6431), .A(n6432), .ZN(n6429) );
  NAND3_X4 U2631 ( .A1(n3306), .A2(n3305), .A3(n3304), .ZN(n3719) );
  NOR2_X4 U2632 ( .A1(n6188), .A2(n6189), .ZN(n3306) );
  NAND2_X4 U2633 ( .A1(n5198), .A2(n4445), .ZN(n5555) );
  OAI221_X2 U2634 ( .B1(n6569), .B2(n3155), .C1(n4482), .C2(n3184), .A(n4481), 
        .ZN(n5198) );
  NOR2_X4 U2635 ( .A1(n3687), .A2(n6277), .ZN(n2585) );
  NAND2_X4 U2636 ( .A1(n3685), .A2(n2698), .ZN(n3687) );
  NOR2_X4 U2637 ( .A1(n3729), .A2(n6263), .ZN(n2586) );
  NAND2_X4 U2638 ( .A1(n3727), .A2(n2696), .ZN(n3729) );
  INV_X4 U2639 ( .A(n6190), .ZN(n2581) );
  INV_X4 U2640 ( .A(n2581), .ZN(n2582) );
  INV_X1 U2641 ( .A(n2581), .ZN(n2583) );
  INV_X16 U2642 ( .A(n3150), .ZN(n4129) );
  INV_X4 U2643 ( .A(n3220), .ZN(n3222) );
  INV_X8 U2644 ( .A(n3220), .ZN(n3221) );
  NAND2_X2 U2645 ( .A1(n5261), .A2(n4975), .ZN(n6018) );
  INV_X8 U2646 ( .A(n3072), .ZN(n3073) );
  INV_X4 U2647 ( .A(n4152), .ZN(n3072) );
  INV_X4 U2648 ( .A(n3175), .ZN(n3179) );
  NOR2_X2 U2649 ( .A1(n6213), .A2(n6269), .ZN(n3338) );
  OAI21_X2 U2650 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n5490) );
  AOI21_X2 U2651 ( .B1(n4257), .B2(n4256), .A(n4255), .ZN(n4258) );
  NAND3_X2 U2652 ( .A1(n4252), .A2(n4251), .A3(n3925), .ZN(n4259) );
  NOR3_X2 U2653 ( .A1(n5268), .A2(n3156), .A3(n5267), .ZN(n5296) );
  NOR3_X2 U2654 ( .A1(n5293), .A2(n5292), .A3(n5291), .ZN(n5294) );
  INV_X16 U2655 ( .A(n3145), .ZN(n4355) );
  INV_X8 U2656 ( .A(n3235), .ZN(n3233) );
  INV_X4 U2657 ( .A(n4525), .ZN(n3170) );
  NAND2_X2 U2658 ( .A1(n5045), .A2(n2588), .ZN(n5749) );
  NOR3_X2 U2659 ( .A1(n5841), .A2(n5043), .A3(n5840), .ZN(n5045) );
  NAND2_X2 U2660 ( .A1(n5836), .A2(n5889), .ZN(n5043) );
  INV_X8 U2661 ( .A(n5705), .ZN(n4966) );
  NAND2_X2 U2662 ( .A1(n4792), .A2(n5397), .ZN(n4658) );
  NAND3_X2 U2663 ( .A1(n5151), .A2(n4438), .A3(n5150), .ZN(n4448) );
  NAND3_X2 U2664 ( .A1(n4444), .A2(n5148), .A3(n5149), .ZN(n4447) );
  NAND2_X2 U2665 ( .A1(iAddr[17]), .A2(iAddr[21]), .ZN(n3678) );
  NOR2_X2 U2666 ( .A1(n4591), .A2(n3137), .ZN(n4593) );
  INV_X4 U2667 ( .A(n5346), .ZN(n4592) );
  NAND2_X2 U2668 ( .A1(n6018), .A2(n4975), .ZN(n6022) );
  NAND4_X2 U2669 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .ZN(n6015)
         );
  NAND3_X2 U2670 ( .A1(n4530), .A2(n4537), .A3(n4529), .ZN(n4542) );
  AOI21_X2 U2671 ( .B1(n4538), .B2(n4537), .A(n4536), .ZN(n4541) );
  NOR2_X2 U2672 ( .A1(n4523), .A2(n4544), .ZN(n4730) );
  NOR2_X2 U2673 ( .A1(n3368), .A2(n3476), .ZN(n3369) );
  NOR2_X2 U2674 ( .A1(n3341), .A2(n3340), .ZN(n3437) );
  NOR2_X2 U2675 ( .A1(n6214), .A2(n6268), .ZN(n3340) );
  NOR2_X2 U2676 ( .A1(n3580), .A2(n3574), .ZN(n3341) );
  OAI22_X2 U2677 ( .A1(n6215), .A2(n6267), .B1(n3403), .B2(n3437), .ZN(n3411)
         );
  NAND3_X2 U2678 ( .A1(n3671), .A2(iAddr[8]), .A3(iAddr[7]), .ZN(n3739) );
  INV_X4 U2679 ( .A(n3743), .ZN(n3671) );
  INV_X4 U2680 ( .A(n4679), .ZN(n4763) );
  NOR2_X2 U2681 ( .A1(n3075), .A2(n4384), .ZN(n4385) );
  NAND2_X2 U2682 ( .A1(n5586), .A2(n4445), .ZN(n5581) );
  NAND2_X2 U2683 ( .A1(n4279), .A2(n4278), .ZN(n4281) );
  NAND3_X2 U2684 ( .A1(n4276), .A2(n4275), .A3(n4274), .ZN(n4282) );
  AOI21_X2 U2685 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n4226) );
  NAND3_X2 U2686 ( .A1(n4311), .A2(n4310), .A3(n4309), .ZN(n6091) );
  OAI21_X2 U2687 ( .B1(n5768), .B2(n5767), .A(n5766), .ZN(n5770) );
  NOR2_X2 U2688 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  NOR3_X2 U2689 ( .A1(n5241), .A2(n5247), .A3(n5469), .ZN(n5250) );
  NAND3_X1 U2690 ( .A1(n4440), .A2(\wb/dsize_reg/z2 [31]), .A3(n3167), .ZN(
        n3924) );
  INV_X4 U2691 ( .A(n3234), .ZN(n3232) );
  INV_X4 U2692 ( .A(n3236), .ZN(n3234) );
  OAI21_X2 U2693 ( .B1(n3576), .B2(n3575), .A(n3574), .ZN(n3578) );
  NOR2_X2 U2694 ( .A1(n3572), .A2(n3625), .ZN(n3573) );
  OAI21_X2 U2695 ( .B1(n3417), .B2(n3416), .A(n3142), .ZN(n3420) );
  INV_X4 U2696 ( .A(n3657), .ZN(n3142) );
  NAND2_X2 U2697 ( .A1(n6229), .A2(n3202), .ZN(n3657) );
  INV_X4 U2698 ( .A(n3142), .ZN(n3143) );
  AOI21_X2 U2699 ( .B1(n4056), .B2(n3177), .A(n4055), .ZN(n4057) );
  NOR2_X2 U2700 ( .A1(n4062), .A2(n4061), .ZN(n4066) );
  NAND3_X2 U2701 ( .A1(reg31Val_0[19]), .A2(n3170), .A3(n3153), .ZN(n4065) );
  NAND4_X2 U2702 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4228)
         );
  NOR2_X2 U2703 ( .A1(n4138), .A2(n4137), .ZN(n4143) );
  NAND3_X2 U2704 ( .A1(n4964), .A2(n4963), .A3(n4962), .ZN(n5681) );
  NOR3_X2 U2705 ( .A1(n5057), .A2(n5747), .A3(n5063), .ZN(n5065) );
  NOR2_X2 U2706 ( .A1(n5063), .A2(n5062), .ZN(n5064) );
  NAND3_X2 U2707 ( .A1(n3088), .A2(n4560), .A3(n4561), .ZN(n5386) );
  NAND3_X2 U2708 ( .A1(n4698), .A2(n4697), .A3(n4696), .ZN(n5262) );
  NAND3_X2 U2709 ( .A1(n4590), .A2(n4589), .A3(n4588), .ZN(n5322) );
  NAND3_X2 U2710 ( .A1(n4202), .A2(n4201), .A3(n4200), .ZN(n5704) );
  NOR3_X2 U2711 ( .A1(n4615), .A2(n4614), .A3(n4613), .ZN(n4620) );
  INV_X4 U2712 ( .A(n2626), .ZN(n5948) );
  NOR2_X2 U2713 ( .A1(n3245), .A2(n3233), .ZN(n4171) );
  NOR2_X2 U2714 ( .A1(n2994), .A2(n3108), .ZN(n5037) );
  NAND2_X2 U2715 ( .A1(n4598), .A2(n5339), .ZN(n5326) );
  AOI21_X2 U2716 ( .B1(n4563), .B2(n4616), .A(n4562), .ZN(n4564) );
  NAND2_X2 U2717 ( .A1(n2680), .A2(regWrData[13]), .ZN(n4559) );
  NAND3_X2 U2718 ( .A1(n4642), .A2(n4641), .A3(n4640), .ZN(n5574) );
  NAND3_X1 U2719 ( .A1(n4639), .A2(n4638), .A3(n4637), .ZN(n4640) );
  NAND2_X2 U2720 ( .A1(n2605), .A2(n5305), .ZN(n5307) );
  NAND2_X2 U2721 ( .A1(n5458), .A2(n5233), .ZN(n5725) );
  OAI21_X2 U2722 ( .B1(n3057), .B2(n5237), .A(n5727), .ZN(n5470) );
  NOR2_X2 U2723 ( .A1(n6010), .A2(n5709), .ZN(n5710) );
  INV_X4 U2724 ( .A(n3138), .ZN(n3175) );
  NOR2_X2 U2725 ( .A1(n3547), .A2(n3463), .ZN(n3361) );
  NOR2_X2 U2726 ( .A1(n2670), .A2(n3172), .ZN(n4396) );
  NOR3_X2 U2727 ( .A1(n4390), .A2(n6301), .A3(n3173), .ZN(n4393) );
  NOR3_X2 U2728 ( .A1(n4391), .A2(n3173), .A3(n2874), .ZN(n4392) );
  INV_X4 U2729 ( .A(n4774), .ZN(n4837) );
  NOR3_X2 U2730 ( .A1(n4794), .A2(n4793), .A3(n5338), .ZN(n4795) );
  NOR2_X2 U2731 ( .A1(n4736), .A2(n5271), .ZN(n4737) );
  NAND2_X2 U2732 ( .A1(n5740), .A2(n5102), .ZN(n5244) );
  NAND2_X2 U2733 ( .A1(n4324), .A2(n4323), .ZN(n4326) );
  NOR2_X2 U2734 ( .A1(n4292), .A2(n3245), .ZN(n4294) );
  NOR2_X2 U2735 ( .A1(n4291), .A2(n4290), .ZN(n4296) );
  NAND2_X2 U2736 ( .A1(n5921), .A2(n5922), .ZN(n5840) );
  INV_X4 U2737 ( .A(n5470), .ZN(n5467) );
  NAND3_X2 U2738 ( .A1(n5244), .A2(n3056), .A3(n5243), .ZN(n5466) );
  NAND2_X2 U2739 ( .A1(n5903), .A2(n5022), .ZN(n5889) );
  INV_X4 U2740 ( .A(n5216), .ZN(n4838) );
  NAND2_X2 U2741 ( .A1(n5040), .A2(n5015), .ZN(n5919) );
  NAND4_X2 U2742 ( .A1(n4674), .A2(n4672), .A3(n5398), .A4(n4673), .ZN(n5941)
         );
  NOR3_X2 U2743 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(n4674) );
  INV_X4 U2744 ( .A(n4227), .ZN(n4981) );
  AOI211_X2 U2745 ( .C1(n6015), .C2(n6014), .A(n6013), .B(n6012), .ZN(n6035)
         );
  NOR2_X2 U2746 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  NAND3_X2 U2747 ( .A1(n6022), .A2(n6021), .A3(n6020), .ZN(n6034) );
  NAND3_X2 U2748 ( .A1(n6019), .A2(n6018), .A3(n4867), .ZN(n6020) );
  NAND2_X1 U2749 ( .A1(n4357), .A2(n2950), .ZN(n4300) );
  OAI21_X2 U2750 ( .B1(n3515), .B2(n3516), .A(n3350), .ZN(n3351) );
  OAI21_X2 U2751 ( .B1(n3449), .B2(n3353), .A(n3454), .ZN(n3474) );
  NAND2_X2 U2752 ( .A1(n3602), .A2(n3601), .ZN(n3619) );
  NOR2_X2 U2753 ( .A1(n3620), .A2(n3342), .ZN(n3377) );
  NAND3_X2 U2754 ( .A1(n3440), .A2(n3606), .A3(n3414), .ZN(n3342) );
  OAI21_X2 U2755 ( .B1(n4473), .B2(n4330), .A(n4331), .ZN(n4337) );
  NAND2_X2 U2756 ( .A1(reg31Val_3[0]), .A2(n2840), .ZN(n3755) );
  NAND2_X2 U2757 ( .A1(n6486), .A2(n6478), .ZN(n6448) );
  NAND3_X2 U2758 ( .A1(n3670), .A2(iAddr[6]), .A3(iAddr[5]), .ZN(n3743) );
  INV_X4 U2759 ( .A(iAddr[19]), .ZN(n3675) );
  NAND2_X2 U2760 ( .A1(n3773), .A2(iAddr[18]), .ZN(n3777) );
  INV_X4 U2761 ( .A(n3775), .ZN(n3773) );
  NOR2_X2 U2762 ( .A1(n3669), .A2(n3668), .ZN(n3673) );
  NOR3_X2 U2763 ( .A1(n3944), .A2(n3943), .A3(n3942), .ZN(n3948) );
  NOR3_X2 U2764 ( .A1(n4390), .A2(n6337), .A3(n3173), .ZN(n3944) );
  NAND3_X2 U2765 ( .A1(n3990), .A2(n4153), .A3(n3167), .ZN(n4276) );
  NOR2_X2 U2766 ( .A1(n3172), .A2(n2898), .ZN(n3989) );
  NAND3_X2 U2767 ( .A1(n3986), .A2(n3232), .A3(n3176), .ZN(n4278) );
  NOR2_X2 U2768 ( .A1(n3172), .A2(n2889), .ZN(n3986) );
  NAND2_X2 U2769 ( .A1(n4524), .A2(memAddr[8]), .ZN(n4283) );
  NAND2_X2 U2770 ( .A1(n5188), .A2(n3041), .ZN(n4774) );
  INV_X4 U2771 ( .A(n3058), .ZN(n3059) );
  NAND3_X2 U2772 ( .A1(n4402), .A2(n4401), .A3(n4400), .ZN(n4410) );
  NAND3_X2 U2773 ( .A1(n4407), .A2(n4405), .A3(n4406), .ZN(n4409) );
  INV_X4 U2774 ( .A(n5678), .ZN(n5091) );
  INV_X1 U2775 ( .A(n3186), .ZN(n3200) );
  NAND3_X2 U2776 ( .A1(n4421), .A2(n4420), .A3(n4419), .ZN(n5185) );
  INV_X4 U2777 ( .A(n3203), .ZN(n3202) );
  NOR2_X2 U2778 ( .A1(n4753), .A2(n6036), .ZN(n4756) );
  OAI21_X1 U2779 ( .B1(n5650), .B2(n5399), .A(n5917), .ZN(n5401) );
  NAND3_X2 U2780 ( .A1(n4516), .A2(n4515), .A3(n4445), .ZN(n5404) );
  NAND2_X2 U2781 ( .A1(n3099), .A2(n3100), .ZN(n4602) );
  NAND2_X2 U2782 ( .A1(n5492), .A2(n3098), .ZN(n3100) );
  NOR2_X2 U2783 ( .A1(n2777), .A2(n4924), .ZN(n4830) );
  INV_X4 U2784 ( .A(n2680), .ZN(n3185) );
  INV_X4 U2785 ( .A(n2723), .ZN(n3155) );
  NAND3_X2 U2786 ( .A1(n6076), .A2(n6075), .A3(n6603), .ZN(n6077) );
  NOR2_X2 U2787 ( .A1(setInv_2), .A2(n2787), .ZN(n6089) );
  OAI21_X2 U2788 ( .B1(n2622), .B2(n6094), .A(n2602), .ZN(n6095) );
  NOR2_X2 U2789 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NOR2_X2 U2790 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NOR2_X2 U2791 ( .A1(n6088), .A2(n6087), .ZN(n6093) );
  NAND2_X2 U2792 ( .A1(n6046), .A2(n6045), .ZN(n6101) );
  NAND3_X1 U2793 ( .A1(\wb/dsize_reg/z2 [1]), .A2(n4001), .A3(n3176), .ZN(
        n4612) );
  NAND3_X1 U2794 ( .A1(reg31Val_0[1]), .A2(n3232), .A3(n3176), .ZN(n4611) );
  NOR2_X2 U2795 ( .A1(n4442), .A2(n3124), .ZN(n3123) );
  NAND3_X1 U2796 ( .A1(reg31Val_0[4]), .A2(n3232), .A3(n3176), .ZN(n4213) );
  NAND2_X2 U2797 ( .A1(n4153), .A2(n3167), .ZN(n4442) );
  NAND3_X2 U2798 ( .A1(\wb/dsize_reg/z2 [6]), .A2(n4010), .A3(n3167), .ZN(
        n4381) );
  NAND3_X1 U2799 ( .A1(reg31Val_0[6]), .A2(n3232), .A3(n3176), .ZN(n4380) );
  AOI21_X2 U2800 ( .B1(n4012), .B2(n3177), .A(n4011), .ZN(n4386) );
  NOR2_X1 U2801 ( .A1(n2687), .A2(n3073), .ZN(n4012) );
  NOR2_X2 U2802 ( .A1(n2783), .A2(n4528), .ZN(n4011) );
  INV_X8 U2803 ( .A(n3073), .ZN(n4153) );
  NAND2_X2 U2804 ( .A1(n4045), .A2(n3105), .ZN(n4264) );
  NOR2_X1 U2805 ( .A1(n2665), .A2(n3073), .ZN(n4045) );
  NAND2_X2 U2806 ( .A1(n4015), .A2(n3167), .ZN(n4577) );
  NAND3_X1 U2807 ( .A1(n3177), .A2(n2811), .A3(n4357), .ZN(n4576) );
  NAND3_X2 U2808 ( .A1(n4355), .A2(n3177), .A3(\wb/dsize_reg/z2 [11]), .ZN(
        n4579) );
  NAND3_X2 U2809 ( .A1(n3177), .A2(n3232), .A3(reg31Val_0[11]), .ZN(n4578) );
  NOR2_X1 U2810 ( .A1(n2686), .A2(n3073), .ZN(n4035) );
  NOR2_X1 U2811 ( .A1(n2673), .A2(n3073), .ZN(n4039) );
  INV_X4 U2812 ( .A(n4104), .ZN(n4170) );
  AOI21_X2 U2813 ( .B1(n3516), .B2(n3523), .A(n3515), .ZN(n3518) );
  AOI21_X2 U2814 ( .B1(n3605), .B2(n3606), .A(n3143), .ZN(n3604) );
  NAND2_X2 U2815 ( .A1(n3590), .A2(n3589), .ZN(n3592) );
  NOR2_X2 U2816 ( .A1(n3614), .A2(n3621), .ZN(n3587) );
  OAI21_X2 U2817 ( .B1(n3580), .B2(n3579), .A(n3142), .ZN(n3583) );
  OAI21_X2 U2818 ( .B1(n3413), .B2(n3610), .A(n3412), .ZN(n3415) );
  NOR2_X2 U2819 ( .A1(n3580), .A2(n3403), .ZN(n3404) );
  NOR2_X2 U2820 ( .A1(n3424), .A2(n3143), .ZN(n3432) );
  AOI21_X1 U2821 ( .B1(n3423), .B2(n2692), .A(n3422), .ZN(n3424) );
  NAND2_X2 U2822 ( .A1(n3201), .A2(n2596), .ZN(n3757) );
  OAI21_X2 U2823 ( .B1(n6222), .B2(n6260), .A(n3807), .ZN(n3387) );
  NOR2_X2 U2824 ( .A1(n6511), .A2(n3204), .ZN(n3390) );
  INV_X4 U2825 ( .A(n3285), .ZN(n3281) );
  NOR2_X1 U2826 ( .A1(n3197), .A2(n2837), .ZN(n6133) );
  INV_X4 U2827 ( .A(n3202), .ZN(n3215) );
  NOR2_X2 U2828 ( .A1(n3664), .A2(n3663), .ZN(n3681) );
  NOR2_X2 U2829 ( .A1(n3667), .A2(n3666), .ZN(n3680) );
  AOI21_X2 U2830 ( .B1(n3750), .B2(n3749), .A(n3748), .ZN(n3828) );
  NOR2_X2 U2831 ( .A1(n3197), .A2(n3302), .ZN(n6132) );
  NOR2_X2 U2832 ( .A1(n3196), .A2(n6369), .ZN(n3889) );
  OAI21_X2 U2833 ( .B1(n3793), .B2(n3792), .A(n3791), .ZN(n3794) );
  AOI21_X2 U2834 ( .B1(n3764), .B2(n3763), .A(n3766), .ZN(n3922) );
  NAND3_X2 U2835 ( .A1(reg31Val_0[25]), .A2(n3170), .A3(n3969), .ZN(n3970) );
  NOR3_X2 U2836 ( .A1(n3968), .A2(n3967), .A3(n3966), .ZN(n3972) );
  NAND3_X2 U2837 ( .A1(n3170), .A2(\wb/dsize_reg/z2 [25]), .A3(n4114), .ZN(
        n3971) );
  NAND2_X2 U2838 ( .A1(n4524), .A2(memAddr[2]), .ZN(n4164) );
  NAND3_X2 U2839 ( .A1(n4023), .A2(n4022), .A3(n4021), .ZN(n4375) );
  NAND3_X2 U2840 ( .A1(reg31Val_0[29]), .A2(n3170), .A3(n3945), .ZN(n4021) );
  NOR3_X2 U2841 ( .A1(n4020), .A2(n4019), .A3(n4018), .ZN(n4023) );
  NAND3_X2 U2842 ( .A1(n3171), .A2(\wb/dsize_reg/z2 [29]), .A3(n4114), .ZN(
        n4022) );
  NAND2_X2 U2843 ( .A1(n4283), .A2(n4284), .ZN(n4290) );
  NAND2_X2 U2844 ( .A1(n4129), .A2(n2634), .ZN(n4263) );
  NOR2_X2 U2845 ( .A1(n3122), .A2(n6555), .ZN(n3121) );
  NAND2_X2 U2846 ( .A1(n4524), .A2(memAddr[15]), .ZN(n4233) );
  NAND3_X2 U2847 ( .A1(n3171), .A2(n3177), .A3(n4103), .ZN(n4107) );
  NAND3_X2 U2848 ( .A1(n4117), .A2(n4116), .A3(n4115), .ZN(n4413) );
  NAND3_X2 U2849 ( .A1(reg31Val_0[20]), .A2(n3170), .A3(n3969), .ZN(n4115) );
  NOR3_X2 U2850 ( .A1(n4113), .A2(n4112), .A3(n4111), .ZN(n4117) );
  NAND3_X2 U2851 ( .A1(n3170), .A2(\wb/dsize_reg/z2 [20]), .A3(n4114), .ZN(
        n4116) );
  NAND3_X2 U2852 ( .A1(n4355), .A2(n3177), .A3(n4119), .ZN(n4122) );
  NOR2_X2 U2853 ( .A1(n4548), .A2(n4735), .ZN(n4549) );
  AOI21_X2 U2854 ( .B1(n4546), .B2(n3226), .A(n4763), .ZN(n4550) );
  NOR2_X2 U2855 ( .A1(n4742), .A2(n2592), .ZN(n4743) );
  NOR2_X2 U2856 ( .A1(n2627), .A2(n4900), .ZN(n4744) );
  OAI21_X2 U2857 ( .B1(n3228), .B2(n4809), .A(n4816), .ZN(n4810) );
  NOR2_X2 U2858 ( .A1(n5179), .A2(n2592), .ZN(n4823) );
  OAI21_X2 U2859 ( .B1(n2842), .B2(n4820), .A(n4819), .ZN(n4821) );
  NOR2_X2 U2860 ( .A1(n5938), .A2(n6029), .ZN(n4820) );
  OAI21_X2 U2861 ( .B1(n4816), .B2(n3230), .A(n3227), .ZN(n4817) );
  NOR2_X2 U2862 ( .A1(n5972), .A2(n2718), .ZN(n4919) );
  INV_X4 U2863 ( .A(n5068), .ZN(n5071) );
  NOR2_X2 U2864 ( .A1(n3228), .A2(n5067), .ZN(n5072) );
  OAI21_X2 U2865 ( .B1(n5120), .B2(n2627), .A(n5090), .ZN(n5095) );
  NOR2_X2 U2866 ( .A1(n5091), .A2(n2626), .ZN(n5094) );
  NOR2_X2 U2867 ( .A1(n5092), .A2(n2592), .ZN(n5093) );
  NOR2_X2 U2868 ( .A1(n5075), .A2(n2778), .ZN(n5076) );
  INV_X4 U2869 ( .A(n5111), .ZN(n5114) );
  OAI21_X2 U2870 ( .B1(n5111), .B2(n3230), .A(n3227), .ZN(n5112) );
  NOR2_X2 U2871 ( .A1(n3228), .A2(n5110), .ZN(n5115) );
  BUF_X4 U2872 ( .A(n6048), .Z(n3129) );
  NOR2_X2 U2873 ( .A1(n5482), .A2(n2778), .ZN(n5117) );
  INV_X8 U2874 ( .A(n3173), .ZN(n3171) );
  INV_X4 U2875 ( .A(n3195), .ZN(n3194) );
  INV_X4 U2876 ( .A(n3200), .ZN(n3196) );
  NOR2_X2 U2877 ( .A1(n5184), .A2(n5183), .ZN(n5194) );
  NOR3_X2 U2878 ( .A1(n5186), .A2(n3209), .A3(n5185), .ZN(n5193) );
  NOR3_X2 U2879 ( .A1(n5173), .A2(n5545), .A3(n5172), .ZN(n5177) );
  NOR2_X2 U2880 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NOR2_X2 U2881 ( .A1(n5897), .A2(n5656), .ZN(n5201) );
  NOR2_X2 U2882 ( .A1(n5195), .A2(n5262), .ZN(n5203) );
  NOR2_X1 U2883 ( .A1(n5209), .A2(n2778), .ZN(n5214) );
  NOR2_X2 U2884 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  OAI21_X2 U2885 ( .B1(n5216), .B2(n3230), .A(n3227), .ZN(n5210) );
  OAI21_X2 U2886 ( .B1(n5720), .B2(n3230), .A(n3227), .ZN(n5254) );
  NOR2_X2 U2887 ( .A1(n3228), .A2(n5253), .ZN(n5256) );
  NOR2_X1 U2888 ( .A1(n5301), .A2(n2626), .ZN(n5317) );
  NOR2_X2 U2889 ( .A1(n5315), .A2(n2627), .ZN(n5316) );
  OAI21_X2 U2890 ( .B1(n5602), .B2(n2778), .A(n5263), .ZN(n5318) );
  NOR2_X2 U2891 ( .A1(n5601), .A2(n2779), .ZN(n5258) );
  NOR2_X2 U2892 ( .A1(n2718), .A2(n5345), .ZN(n5350) );
  AOI21_X2 U2893 ( .B1(n3226), .B2(n5348), .A(n5347), .ZN(n5349) );
  NAND3_X2 U2894 ( .A1(n4729), .A2(n4728), .A3(n4727), .ZN(n5387) );
  NOR2_X2 U2895 ( .A1(n2718), .A2(n5376), .ZN(n5382) );
  NOR2_X2 U2896 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  OAI21_X2 U2897 ( .B1(n5377), .B2(n3229), .A(n3227), .ZN(n5378) );
  NOR2_X2 U2898 ( .A1(n5986), .A2(n2718), .ZN(n5426) );
  OAI21_X2 U2899 ( .B1(n5492), .B2(n3229), .A(n6008), .ZN(n5493) );
  NOR2_X2 U2900 ( .A1(n5502), .A2(n5501), .ZN(n5507) );
  NOR2_X2 U2901 ( .A1(n5976), .A2(n2718), .ZN(n5558) );
  AOI21_X2 U2902 ( .B1(n3226), .B2(n5556), .A(n5555), .ZN(n5557) );
  NOR2_X2 U2903 ( .A1(n5561), .A2(n2592), .ZN(n5562) );
  OAI21_X2 U2904 ( .B1(n3156), .B2(n3229), .A(n3226), .ZN(n5580) );
  NOR2_X2 U2905 ( .A1(n5973), .A2(n2718), .ZN(n5584) );
  NOR2_X2 U2906 ( .A1(n5602), .A2(n2626), .ZN(n5605) );
  NOR2_X2 U2907 ( .A1(n5603), .A2(n2592), .ZN(n5604) );
  OAI21_X2 U2908 ( .B1(n5595), .B2(n3228), .A(n6040), .ZN(n5596) );
  NOR2_X2 U2909 ( .A1(n5600), .A2(n3229), .ZN(n5595) );
  NOR2_X2 U2910 ( .A1(n2718), .A2(n5594), .ZN(n5598) );
  NOR2_X2 U2911 ( .A1(n5877), .A2(n2626), .ZN(n5654) );
  NOR2_X1 U2912 ( .A1(n5982), .A2(n2718), .ZN(n5655) );
  AOI21_X2 U2913 ( .B1(n3226), .B2(n5635), .A(n5634), .ZN(n5636) );
  NOR2_X2 U2914 ( .A1(n5975), .A2(n2718), .ZN(n5675) );
  NOR2_X2 U2915 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  OAI21_X2 U2916 ( .B1(n5670), .B2(n3229), .A(n6008), .ZN(n5671) );
  NOR2_X2 U2917 ( .A1(n5602), .A2(n2779), .ZN(n5776) );
  NOR2_X2 U2918 ( .A1(n6091), .A2(n3226), .ZN(n5774) );
  NAND3_X2 U2919 ( .A1(n4927), .A2(n4926), .A3(n4925), .ZN(n5802) );
  AOI21_X2 U2920 ( .B1(n5447), .B2(n5127), .A(n2905), .ZN(n4925) );
  NOR2_X2 U2921 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  OAI21_X2 U2922 ( .B1(n5816), .B2(n3229), .A(n6008), .ZN(n5810) );
  NOR2_X2 U2923 ( .A1(n5877), .A2(n2778), .ZN(n5882) );
  NOR2_X2 U2924 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  OAI21_X2 U2925 ( .B1(n5884), .B2(n3229), .A(n6008), .ZN(n5878) );
  NOR2_X2 U2926 ( .A1(n5359), .A2(n5358), .ZN(n5362) );
  NOR2_X2 U2927 ( .A1(n5906), .A2(n2778), .ZN(n5911) );
  NOR2_X2 U2928 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  OAI21_X2 U2929 ( .B1(n5913), .B2(n3229), .A(n6008), .ZN(n5907) );
  OAI21_X2 U2930 ( .B1(n2842), .B2(n5952), .A(n5951), .ZN(n5953) );
  NOR2_X2 U2931 ( .A1(n5948), .A2(n5947), .ZN(n5952) );
  OAI21_X2 U2932 ( .B1(n5946), .B2(n2718), .A(n5945), .ZN(n5954) );
  INV_X4 U2933 ( .A(n2627), .ZN(n5938) );
  OAI21_X2 U2934 ( .B1(n4609), .B2(n3184), .A(n4608), .ZN(n5940) );
  INV_X4 U2935 ( .A(n6057), .ZN(n6052) );
  NAND3_X1 U2936 ( .A1(n3998), .A2(n4624), .A3(n4623), .ZN(regWrData[2]) );
  NAND2_X2 U2937 ( .A1(n3102), .A2(n3925), .ZN(regWrData[7]) );
  AOI22_X2 U2938 ( .A1(n4291), .A2(n3178), .B1(n4292), .B2(n3178), .ZN(n4031)
         );
  NAND4_X2 U2939 ( .A1(n4042), .A2(n4041), .A3(n4339), .A4(n4040), .ZN(
        regWrData[13]) );
  NAND3_X2 U2940 ( .A1(n3232), .A2(reg31Val_0[13]), .A3(n3167), .ZN(n4042) );
  NAND3_X1 U2941 ( .A1(n2848), .A2(n4357), .A3(n3167), .ZN(n4041) );
  NAND2_X2 U2942 ( .A1(\wb/dsize_reg/z2 [13]), .A2(n3151), .ZN(n4040) );
  OAI21_X2 U2943 ( .B1(n6372), .B2(n3895), .A(n3894), .ZN(n2129) );
  NOR2_X2 U2944 ( .A1(n3109), .A2(n5538), .ZN(n3108) );
  NOR2_X2 U2945 ( .A1(n4632), .A2(n4631), .ZN(n4633) );
  NOR2_X2 U2946 ( .A1(n4636), .A2(n4639), .ZN(n4632) );
  NOR2_X2 U2947 ( .A1(n4630), .A2(n4629), .ZN(n4631) );
  NOR3_X2 U2948 ( .A1(n4427), .A2(n4450), .A3(n4426), .ZN(n4437) );
  NOR2_X2 U2949 ( .A1(n4427), .A2(n4816), .ZN(n4371) );
  NOR2_X2 U2950 ( .A1(n5720), .A2(n4273), .ZN(n4370) );
  NOR2_X2 U2951 ( .A1(n4377), .A2(n4431), .ZN(n4418) );
  NAND3_X2 U2952 ( .A1(n4838), .A2(n5005), .A3(n5860), .ZN(n4377) );
  NOR2_X2 U2953 ( .A1(n4416), .A2(n4415), .ZN(n4417) );
  NAND3_X2 U2954 ( .A1(n4453), .A2(n4846), .A3(n5071), .ZN(n4415) );
  INV_X4 U2955 ( .A(n3108), .ZN(n5032) );
  NOR3_X2 U2956 ( .A1(n5738), .A2(n3057), .A3(n5736), .ZN(n5743) );
  INV_X4 U2957 ( .A(n5734), .ZN(n5738) );
  NOR2_X2 U2958 ( .A1(n4330), .A2(n3174), .ZN(n3103) );
  NAND2_X2 U2959 ( .A1(n4657), .A2(n5395), .ZN(n4792) );
  NOR2_X2 U2960 ( .A1(zeroExt_2), .A2(n4590), .ZN(n4591) );
  AOI21_X2 U2961 ( .B1(n3085), .B2(n4321), .A(n3245), .ZN(n4324) );
  NAND2_X2 U2962 ( .A1(n5639), .A2(n4603), .ZN(n5528) );
  NAND3_X2 U2963 ( .A1(reg31Val_0[1]), .A2(n3243), .A3(n3232), .ZN(n4173) );
  NAND2_X2 U2964 ( .A1(n5572), .A2(n5575), .ZN(n4644) );
  NOR2_X2 U2965 ( .A1(n5785), .A2(n4975), .ZN(n4974) );
  NOR2_X2 U2966 ( .A1(n5555), .A2(n4975), .ZN(n4976) );
  NAND2_X2 U2967 ( .A1(n4966), .A2(n4885), .ZN(n5277) );
  NOR2_X2 U2968 ( .A1(n4671), .A2(n4670), .ZN(n4672) );
  NOR2_X2 U2969 ( .A1(n3245), .A2(n2668), .ZN(n4533) );
  NOR2_X2 U2970 ( .A1(n3243), .A2(n6616), .ZN(n4536) );
  NAND3_X2 U2971 ( .A1(n4531), .A2(n3173), .A3(n4532), .ZN(n4537) );
  NOR2_X2 U2972 ( .A1(n3245), .A2(n2667), .ZN(n4529) );
  NOR2_X2 U2973 ( .A1(n5724), .A2(n5723), .ZN(n5728) );
  NOR3_X2 U2974 ( .A1(n5971), .A2(n5970), .A3(n6004), .ZN(n5974) );
  OAI21_X2 U2975 ( .B1(n6015), .B2(n2776), .A(n6008), .ZN(n6009) );
  NAND2_X2 U2976 ( .A1(n4329), .A2(n4328), .ZN(n4330) );
  NAND2_X2 U2977 ( .A1(n5942), .A2(n5041), .ZN(n4770) );
  OAI21_X2 U2978 ( .B1(n4244), .B2(n4245), .A(n4243), .ZN(n4553) );
  NAND2_X2 U2979 ( .A1(n5662), .A2(n4652), .ZN(n5334) );
  INV_X4 U2980 ( .A(n4408), .ZN(n4407) );
  INV_X8 U2981 ( .A(n3187), .ZN(n3186) );
  INV_X4 U2982 ( .A(n5171), .ZN(n3187) );
  NAND2_X2 U2983 ( .A1(n6495), .A2(n3215), .ZN(n5171) );
  NAND4_X2 U2984 ( .A1(n6252), .A2(n6251), .A3(n6448), .A4(n2841), .ZN(n6495)
         );
  INV_X4 U2985 ( .A(n5321), .ZN(n3203) );
  OAI21_X2 U2986 ( .B1(n6228), .B2(n3301), .A(n6227), .ZN(n5321) );
  AOI211_X2 U2987 ( .C1(n4267), .C2(n3177), .A(n4266), .B(n4265), .ZN(n4268)
         );
  NOR2_X2 U2988 ( .A1(n3181), .A2(n3145), .ZN(n4347) );
  NOR2_X2 U2989 ( .A1(n3154), .A2(n2882), .ZN(n4344) );
  NAND2_X2 U2990 ( .A1(n3131), .A2(n3132), .ZN(n4565) );
  NOR3_X2 U2991 ( .A1(n3085), .A2(n4513), .A3(n4512), .ZN(n4514) );
  NOR2_X2 U2992 ( .A1(n4289), .A2(n4288), .ZN(n4298) );
  NOR3_X2 U2993 ( .A1(n3177), .A2(n3244), .A3(n4290), .ZN(n4289) );
  NAND2_X2 U2994 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  NOR2_X2 U2995 ( .A1(n4253), .A2(n3245), .ZN(n4257) );
  NOR2_X2 U2996 ( .A1(n3075), .A2(n4254), .ZN(n4256) );
  NOR2_X2 U2997 ( .A1(n3243), .A2(n2839), .ZN(n4255) );
  INV_X4 U2998 ( .A(n5535), .ZN(n5397) );
  NAND3_X2 U2999 ( .A1(n4700), .A2(n3217), .A3(n4699), .ZN(n5274) );
  OAI21_X2 U3000 ( .B1(n4960), .B2(n4928), .A(n6022), .ZN(n4860) );
  NAND2_X2 U3001 ( .A1(n5396), .A2(n5395), .ZN(n5553) );
  NOR2_X2 U3002 ( .A1(n4384), .A2(n4383), .ZN(n4387) );
  NAND2_X2 U3003 ( .A1(n5611), .A2(n4643), .ZN(n5575) );
  INV_X4 U3004 ( .A(n5574), .ZN(n4643) );
  NOR2_X2 U3005 ( .A1(n3245), .A2(n4183), .ZN(n4185) );
  NAND2_X2 U3006 ( .A1(n4648), .A2(n4647), .ZN(n5592) );
  NOR2_X2 U3007 ( .A1(n2701), .A2(n3073), .ZN(n3995) );
  NAND3_X2 U3008 ( .A1(\wb/dsize_reg/z2 [26]), .A2(n3176), .A3(n4440), .ZN(
        n4626) );
  NOR2_X2 U3009 ( .A1(n4277), .A2(n3245), .ZN(n4279) );
  NOR2_X2 U3010 ( .A1(n4207), .A2(n4206), .ZN(n4212) );
  NOR2_X2 U3011 ( .A1(n4209), .A2(n4208), .ZN(n4211) );
  NOR2_X2 U3012 ( .A1(\wb/dsize_reg/z2 [20]), .A2(n3245), .ZN(n4210) );
  NOR2_X2 U3013 ( .A1(n4217), .A2(n4216), .ZN(n4223) );
  NOR2_X2 U3014 ( .A1(n3245), .A2(n4221), .ZN(n4222) );
  NAND3_X2 U3015 ( .A1(n4220), .A2(n4219), .A3(n4218), .ZN(n4221) );
  NOR2_X2 U3016 ( .A1(n4209), .A2(n3245), .ZN(n4205) );
  NOR2_X2 U3017 ( .A1(n3170), .A2(n4208), .ZN(n4204) );
  NOR2_X2 U3018 ( .A1(n3243), .A2(n2838), .ZN(n4203) );
  NOR2_X2 U3019 ( .A1(n5289), .A2(n5288), .ZN(n5292) );
  NOR3_X2 U3020 ( .A1(n5748), .A2(n5747), .A3(n5853), .ZN(n5753) );
  NOR2_X2 U3021 ( .A1(n3245), .A2(n4302), .ZN(n4308) );
  NOR3_X2 U3022 ( .A1(n4306), .A2(n4305), .A3(n3244), .ZN(n4307) );
  NOR2_X2 U3023 ( .A1(n2887), .A2(n4302), .ZN(n4301) );
  NOR2_X2 U3024 ( .A1(n2891), .A2(n3245), .ZN(n4299) );
  NAND2_X2 U3025 ( .A1(n5514), .A2(n5509), .ZN(n6027) );
  AOI22_X2 U3026 ( .A1(n2605), .A2(n4943), .B1(n2685), .B2(n6017), .ZN(n4956)
         );
  NAND2_X2 U3027 ( .A1(n4851), .A2(n4850), .ZN(n5123) );
  AOI21_X2 U3028 ( .B1(n4929), .B2(n5017), .A(n3218), .ZN(n4851) );
  INV_X4 U3029 ( .A(n5838), .ZN(n5917) );
  NAND2_X2 U3030 ( .A1(n4733), .A2(n4734), .ZN(n4811) );
  NAND3_X2 U3031 ( .A1(n4518), .A2(n3216), .A3(n4517), .ZN(n5121) );
  NAND3_X2 U3032 ( .A1(n4480), .A2(n3216), .A3(n4479), .ZN(n5305) );
  INV_X4 U3033 ( .A(n4975), .ZN(n5082) );
  INV_X4 U3034 ( .A(n3056), .ZN(n3057) );
  NOR2_X2 U3035 ( .A1(n5245), .A2(n5466), .ZN(n5246) );
  NOR2_X2 U3036 ( .A1(n5703), .A2(n5702), .ZN(n5715) );
  NAND3_X2 U3037 ( .A1(\wb/dsize_reg/z2 [25]), .A2(n3176), .A3(n4440), .ZN(
        n4183) );
  NAND3_X2 U3038 ( .A1(reg31Val_0[2]), .A2(n3232), .A3(n3176), .ZN(n4492) );
  NAND2_X2 U3039 ( .A1(n3136), .A2(n4153), .ZN(n4405) );
  NAND3_X2 U3040 ( .A1(reg31Val_0[5]), .A2(n3232), .A3(n3168), .ZN(n4400) );
  NAND2_X2 U3041 ( .A1(n4075), .A2(n3167), .ZN(n4402) );
  NOR2_X2 U3042 ( .A1(n3154), .A2(n2924), .ZN(n4316) );
  INV_X8 U3043 ( .A(n3169), .ZN(n3168) );
  NOR2_X2 U3044 ( .A1(n6202), .A2(n6279), .ZN(n3505) );
  NOR3_X2 U3045 ( .A1(n3372), .A2(n3553), .A3(n3499), .ZN(n3374) );
  NAND2_X2 U3046 ( .A1(n3371), .A2(n3365), .ZN(n3366) );
  NAND3_X2 U3047 ( .A1(n3334), .A2(n3333), .A3(n3436), .ZN(n3335) );
  INV_X4 U3048 ( .A(n3378), .ZN(n3423) );
  NOR2_X2 U3049 ( .A1(n3382), .A2(n3645), .ZN(n3385) );
  NAND3_X2 U3050 ( .A1(n5334), .A2(n5395), .A3(n4913), .ZN(n4890) );
  NOR2_X2 U3051 ( .A1(zeroExt_2), .A2(n2926), .ZN(n4478) );
  OAI21_X2 U3052 ( .B1(n3142), .B2(n3665), .A(iAddr[27]), .ZN(n3663) );
  NOR2_X2 U3053 ( .A1(n3665), .A2(n3806), .ZN(n3664) );
  INV_X4 U3054 ( .A(n3074), .ZN(n3927) );
  NAND3_X2 U3055 ( .A1(n4357), .A2(n2850), .A3(n3075), .ZN(n3074) );
  NOR2_X2 U3056 ( .A1(n4147), .A2(n3172), .ZN(n3930) );
  NOR2_X2 U3057 ( .A1(n2668), .A2(n3145), .ZN(n3928) );
  NOR2_X2 U3058 ( .A1(n2707), .A2(n3172), .ZN(n3951) );
  NOR2_X2 U3059 ( .A1(n2667), .A2(n3172), .ZN(n3959) );
  NOR3_X2 U3060 ( .A1(n4390), .A2(n6334), .A3(n3173), .ZN(n3968) );
  NOR3_X2 U3061 ( .A1(n4390), .A2(n6324), .A3(n3173), .ZN(n4020) );
  NOR2_X2 U3062 ( .A1(n3172), .A2(n4054), .ZN(n4056) );
  NOR2_X2 U3063 ( .A1(n2783), .A2(n3145), .ZN(n4053) );
  NOR2_X2 U3064 ( .A1(n6302), .A2(n3064), .ZN(n4102) );
  NOR3_X2 U3065 ( .A1(n4390), .A2(n6304), .A3(n3173), .ZN(n4113) );
  NOR2_X2 U3066 ( .A1(n6307), .A2(n3172), .ZN(n4120) );
  NOR2_X2 U3067 ( .A1(n2665), .A2(n3172), .ZN(n4119) );
  NOR2_X2 U3068 ( .A1(n2666), .A2(n3172), .ZN(n4126) );
  NOR2_X2 U3069 ( .A1(n4393), .A2(n4392), .ZN(n4398) );
  AOI21_X2 U3070 ( .B1(n4114), .B2(n4396), .A(n4395), .ZN(n4397) );
  OAI21_X2 U3071 ( .B1(n4570), .B2(n4886), .A(n4804), .ZN(n4806) );
  AOI21_X2 U3072 ( .B1(n5221), .B2(n5918), .A(n5832), .ZN(n4843) );
  OAI21_X2 U3073 ( .B1(n4961), .B2(n6019), .A(n6018), .ZN(n5260) );
  NOR2_X2 U3074 ( .A1(n5747), .A2(n5031), .ZN(n5047) );
  NOR2_X2 U3075 ( .A1(n5061), .A2(n5791), .ZN(n5062) );
  INV_X4 U3076 ( .A(n3186), .ZN(n3199) );
  NAND2_X2 U3077 ( .A1(n2680), .A2(regWrData[10]), .ZN(n4590) );
  OAI21_X2 U3078 ( .B1(n5342), .B2(n5498), .A(n5341), .ZN(n5344) );
  AOI21_X2 U3079 ( .B1(n5025), .B2(n5846), .A(n5844), .ZN(n5026) );
  AOI21_X2 U3080 ( .B1(n5018), .B2(n5919), .A(n5840), .ZN(n5028) );
  NOR2_X2 U3081 ( .A1(n5500), .A2(n2777), .ZN(n5501) );
  NOR2_X2 U3082 ( .A1(n3123), .A2(n4194), .ZN(n4195) );
  NOR3_X2 U3083 ( .A1(n4192), .A2(n4191), .A3(n3244), .ZN(n4196) );
  NAND3_X2 U3084 ( .A1(n5143), .A2(n5142), .A3(n4611), .ZN(n4615) );
  NAND2_X2 U3085 ( .A1(n4985), .A2(n5511), .ZN(n3082) );
  INV_X4 U3086 ( .A(n5618), .ZN(n5611) );
  OAI21_X2 U3087 ( .B1(n4961), .B2(n4695), .A(n6018), .ZN(n5448) );
  NAND2_X2 U3088 ( .A1(n5852), .A2(n5851), .ZN(n5854) );
  OAI21_X2 U3089 ( .B1(n4969), .B2(n4968), .A(n3157), .ZN(n4971) );
  NAND2_X2 U3090 ( .A1(n5886), .A2(n5887), .ZN(n5888) );
  NAND2_X2 U3091 ( .A1(n5207), .A2(n3090), .ZN(n5922) );
  INV_X4 U3092 ( .A(n2777), .ZN(n5514) );
  NAND2_X2 U3093 ( .A1(n5962), .A2(n5961), .ZN(n5966) );
  NAND3_X2 U3094 ( .A1(\wb/dsize_reg/z2 [0]), .A2(n4001), .A3(n3176), .ZN(
        n5148) );
  INV_X4 U3095 ( .A(n4027), .ZN(n4291) );
  INV_X4 U3096 ( .A(n4030), .ZN(n4292) );
  NOR2_X2 U3097 ( .A1(n3086), .A2(n3152), .ZN(n3085) );
  NOR2_X2 U3098 ( .A1(n3152), .A2(n2892), .ZN(n4471) );
  NAND3_X2 U3099 ( .A1(n3105), .A2(\wb/dsize_reg/z2 [30]), .A3(n4153), .ZN(
        n3104) );
  NOR2_X2 U3100 ( .A1(n3154), .A2(n2925), .ZN(n4235) );
  NOR2_X2 U3101 ( .A1(n2845), .A2(n3073), .ZN(n4085) );
  NOR2_X2 U3102 ( .A1(n3152), .A2(n2893), .ZN(n4086) );
  NOR2_X2 U3103 ( .A1(n2670), .A2(n3145), .ZN(n4093) );
  NAND2_X2 U3104 ( .A1(n3504), .A2(n3568), .ZN(n3560) );
  AOI21_X2 U3105 ( .B1(n3560), .B2(n2847), .A(n3505), .ZN(n3507) );
  AOI21_X2 U3106 ( .B1(n3498), .B2(n2894), .A(n3497), .ZN(n3500) );
  NOR2_X2 U3107 ( .A1(n3477), .A2(n3476), .ZN(n3479) );
  NOR2_X2 U3108 ( .A1(n3621), .A2(n3620), .ZN(n3623) );
  NAND3_X2 U3109 ( .A1(n2851), .A2(n3593), .A3(n2711), .ZN(n3438) );
  AOI21_X2 U3110 ( .B1(n4881), .B2(n3226), .A(n4880), .ZN(n4882) );
  INV_X4 U3111 ( .A(n3312), .ZN(n3685) );
  NAND2_X2 U3112 ( .A1(n3311), .A2(n2631), .ZN(n3312) );
  NAND2_X2 U3113 ( .A1(n3313), .A2(n2682), .ZN(n3314) );
  NAND2_X2 U3114 ( .A1(n3692), .A2(n3331), .ZN(n3694) );
  INV_X4 U3115 ( .A(n3318), .ZN(n3700) );
  NAND2_X2 U3116 ( .A1(n3317), .A2(n2824), .ZN(n3318) );
  NAND2_X2 U3117 ( .A1(n3321), .A2(n2810), .ZN(n3322) );
  NAND2_X2 U3118 ( .A1(n3309), .A2(n3716), .ZN(n3310) );
  NOR2_X2 U3119 ( .A1(n6177), .A2(n6187), .ZN(n3304) );
  INV_X4 U3120 ( .A(n3719), .ZN(n3307) );
  AOI21_X2 U3121 ( .B1(n3142), .B2(n3754), .A(n3753), .ZN(n3830) );
  NOR2_X2 U3122 ( .A1(n6191), .A2(n3757), .ZN(n3753) );
  NOR2_X2 U3123 ( .A1(n3213), .A2(n3759), .ZN(n3760) );
  OAI21_X2 U3124 ( .B1(n6192), .B2(n3757), .A(n3756), .ZN(n3758) );
  NAND3_X2 U3125 ( .A1(n3142), .A2(n3755), .A3(n2890), .ZN(n3756) );
  INV_X4 U3126 ( .A(n3284), .ZN(n3283) );
  NAND2_X2 U3127 ( .A1(n3325), .A2(n2822), .ZN(n3817) );
  INV_X4 U3128 ( .A(n3284), .ZN(n3282) );
  INV_X4 U3129 ( .A(\mem_wb/N41 ), .ZN(n3295) );
  INV_X4 U3130 ( .A(\mem_wb/N41 ), .ZN(n3298) );
  INV_X4 U3131 ( .A(\mem_wb/N41 ), .ZN(n3297) );
  INV_X4 U3132 ( .A(\mem_wb/N41 ), .ZN(n3296) );
  NOR2_X2 U3133 ( .A1(n2846), .A2(n2797), .ZN(n3684) );
  NOR2_X2 U3134 ( .A1(n6236), .A2(n3211), .ZN(n3683) );
  INV_X4 U3135 ( .A(\mem_wb/N41 ), .ZN(n3285) );
  NOR2_X2 U3136 ( .A1(n6402), .A2(n6400), .ZN(n6401) );
  INV_X4 U3137 ( .A(\mem_wb/N41 ), .ZN(n3286) );
  NOR2_X2 U3138 ( .A1(n2975), .A2(n6396), .ZN(n6381) );
  OAI21_X2 U3139 ( .B1(n6412), .B2(n6588), .A(n3835), .ZN(n3903) );
  NOR2_X2 U3140 ( .A1(n3197), .A2(n2788), .ZN(n3835) );
  INV_X4 U3141 ( .A(n3198), .ZN(n3190) );
  NOR2_X2 U3142 ( .A1(n3812), .A2(n3811), .ZN(n3814) );
  OAI21_X2 U3143 ( .B1(n3803), .B2(iAddr[28]), .A(n3805), .ZN(n3804) );
  AOI21_X2 U3144 ( .B1(n3799), .B2(n3798), .A(n3813), .ZN(n3908) );
  AOI21_X2 U3145 ( .B1(n3677), .B2(n3786), .A(n3785), .ZN(n3911) );
  OAI21_X2 U3146 ( .B1(n3778), .B2(n3777), .A(n3776), .ZN(n3780) );
  AOI21_X2 U3147 ( .B1(n3775), .B2(n3774), .A(n3779), .ZN(n3914) );
  OAI21_X2 U3148 ( .B1(iAddr[14]), .B2(n2876), .A(n3770), .ZN(n3769) );
  INV_X4 U3149 ( .A(n3198), .ZN(n3189) );
  INV_X4 U3150 ( .A(\mem_wb/N41 ), .ZN(n3287) );
  NAND3_X2 U3151 ( .A1(reg31Val_0[22]), .A2(n3170), .A3(n3945), .ZN(n3946) );
  NAND3_X2 U3152 ( .A1(n3170), .A2(\wb/dsize_reg/z2 [22]), .A3(n4114), .ZN(
        n3947) );
  NOR2_X2 U3153 ( .A1(n4759), .A2(n4774), .ZN(n4760) );
  AOI21_X2 U3154 ( .B1(n4996), .B2(n3226), .A(n4995), .ZN(n4997) );
  OAI21_X2 U3155 ( .B1(n5003), .B2(n2776), .A(n3227), .ZN(n4998) );
  INV_X4 U3156 ( .A(\mem_wb/N41 ), .ZN(n3290) );
  INV_X4 U3157 ( .A(\mem_wb/N41 ), .ZN(n3289) );
  NOR2_X2 U3158 ( .A1(n5411), .A2(n2779), .ZN(n5414) );
  NOR2_X2 U3159 ( .A1(n5405), .A2(n5404), .ZN(n5406) );
  NOR2_X2 U3160 ( .A1(n5991), .A2(n2718), .ZN(n5407) );
  AOI21_X2 U3161 ( .B1(n5460), .B2(n3226), .A(n5459), .ZN(n5461) );
  OAI21_X2 U3162 ( .B1(n5463), .B2(n3230), .A(n6008), .ZN(n5464) );
  OAI22_X2 U3163 ( .A1(n5481), .A2(n2626), .B1(n5480), .B2(n2592), .ZN(n5484)
         );
  NOR2_X2 U3164 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND3_X2 U3165 ( .A1(n4833), .A2(n4832), .A3(n4831), .ZN(n5544) );
  NOR2_X2 U3166 ( .A1(n4830), .A2(n4829), .ZN(n4831) );
  NOR2_X2 U3167 ( .A1(n2718), .A2(n5615), .ZN(n5621) );
  NOR2_X2 U3168 ( .A1(n5809), .A2(n2779), .ZN(n5788) );
  NOR2_X2 U3169 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  NOR2_X2 U3170 ( .A1(n5799), .A2(n2592), .ZN(n5800) );
  OAI21_X2 U3171 ( .B1(n5856), .B2(n3229), .A(n6008), .ZN(n5857) );
  NOR2_X2 U3172 ( .A1(n3228), .A2(n5855), .ZN(n5861) );
  OAI21_X2 U3173 ( .B1(n5867), .B2(n2627), .A(n5866), .ZN(n5872) );
  OAI21_X2 U3174 ( .B1(n5870), .B2(n2626), .A(n5869), .ZN(n5871) );
  INV_X4 U3175 ( .A(n6065), .ZN(n5995) );
  NOR2_X2 U3176 ( .A1(n5877), .A2(n2779), .ZN(n5862) );
  NAND3_X2 U3177 ( .A1(setInv_2), .A2(n6075), .A3(n6088), .ZN(n6001) );
  NOR2_X2 U3178 ( .A1(n2602), .A2(n2787), .ZN(n6080) );
  NOR2_X2 U3179 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  NAND3_X2 U3180 ( .A1(n6100), .A2(n2663), .A3(n2595), .ZN(n6102) );
  NAND3_X2 U3181 ( .A1(n5149), .A2(n5148), .A3(n5147), .ZN(regWrData[0]) );
  NOR2_X2 U3182 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  NAND3_X2 U3183 ( .A1(n4007), .A2(n4006), .A3(n4193), .ZN(regWrData[3]) );
  NOR2_X2 U3184 ( .A1(n4190), .A2(n4191), .ZN(n4006) );
  NAND3_X2 U3185 ( .A1(n3982), .A2(n4215), .A3(n3981), .ZN(regWrData[4]) );
  NOR2_X2 U3186 ( .A1(n4206), .A2(n3979), .ZN(n3982) );
  NAND3_X2 U3187 ( .A1(reg31Val_0[9]), .A2(n3232), .A3(n3167), .ZN(n4155) );
  NAND3_X2 U3188 ( .A1(n4151), .A2(n4150), .A3(n4149), .ZN(regWrData[16]) );
  NAND3_X2 U3189 ( .A1(n3977), .A2(n3976), .A3(n3975), .ZN(regWrData[31]) );
  OAI21_X2 U3190 ( .B1(n6523), .B2(n3209), .A(n3831), .ZN(iAddr[0]) );
  OAI21_X2 U3191 ( .B1(n6522), .B2(n3205), .A(n3830), .ZN(iAddr[1]) );
  NAND2_X2 U3192 ( .A1(n3659), .A2(n2903), .ZN(n3531) );
  OAI211_X2 U3193 ( .C1(n3528), .C2(n3657), .A(n3527), .B(n3526), .ZN(iAddr[3]) );
  OAI211_X2 U3194 ( .C1(n3521), .C2(n3657), .A(n3520), .B(n3519), .ZN(iAddr[4]) );
  NAND2_X2 U3195 ( .A1(n3659), .A2(n2901), .ZN(n3520) );
  NAND3_X2 U3196 ( .A1(n3545), .A2(n3544), .A3(n3543), .ZN(iAddr[5]) );
  NAND3_X2 U3197 ( .A1(n3559), .A2(n3558), .A3(n3557), .ZN(iAddr[7]) );
  NAND3_X2 U3198 ( .A1(n3571), .A2(n3570), .A3(n3569), .ZN(iAddr[9]) );
  NAND3_X2 U3199 ( .A1(n3471), .A2(n3470), .A3(n2879), .ZN(iAddr[12]) );
  NAND3_X2 U3200 ( .A1(n3609), .A2(n3608), .A3(n3607), .ZN(iAddr[18]) );
  NAND2_X2 U3201 ( .A1(n3615), .A2(n3142), .ZN(n3617) );
  NAND3_X2 U3202 ( .A1(n3596), .A2(n3595), .A3(n3594), .ZN(iAddr[20]) );
  NOR2_X2 U3203 ( .A1(n3577), .A2(n3578), .ZN(n3584) );
  NOR2_X2 U3204 ( .A1(n3414), .A2(n3415), .ZN(n3421) );
  AOI21_X2 U3205 ( .B1(n3432), .B2(n3431), .A(n3430), .ZN(n3434) );
  NOR2_X2 U3206 ( .A1(n6179), .A2(n3757), .ZN(n3430) );
  NOR2_X2 U3207 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NOR2_X2 U3208 ( .A1(n6224), .A2(n3757), .ZN(n3389) );
  NOR2_X2 U3209 ( .A1(n6517), .A2(n3208), .ZN(\ex_mem/N42 ) );
  NOR2_X2 U3210 ( .A1(n6628), .A2(n3207), .ZN(\ex_mem/N147 ) );
  NOR2_X2 U3211 ( .A1(n6627), .A2(n3207), .ZN(\ex_mem/N148 ) );
  NOR2_X2 U3212 ( .A1(n6542), .A2(n3208), .ZN(\ex_mem/N52 ) );
  NOR2_X2 U3213 ( .A1(n6543), .A2(n3208), .ZN(\ex_mem/N51 ) );
  NOR2_X2 U3214 ( .A1(n6512), .A2(n3209), .ZN(\ex_mem/N40 ) );
  NOR2_X2 U3215 ( .A1(n6518), .A2(n3208), .ZN(\ex_mem/N41 ) );
  NOR2_X2 U3216 ( .A1(n6595), .A2(n3208), .ZN(\ex_mem/N36 ) );
  NOR2_X2 U3217 ( .A1(n6596), .A2(n3208), .ZN(\ex_mem/N35 ) );
  NOR2_X2 U3218 ( .A1(n6606), .A2(n3207), .ZN(\ex_mem/N142 ) );
  NOR2_X2 U3219 ( .A1(n6547), .A2(n3208), .ZN(\ex_mem/N46 ) );
  NOR2_X2 U3220 ( .A1(n6521), .A2(n3208), .ZN(\ex_mem/N37 ) );
  NOR2_X2 U3221 ( .A1(n6520), .A2(n3208), .ZN(\ex_mem/N38 ) );
  NOR2_X2 U3222 ( .A1(n6519), .A2(n3208), .ZN(\ex_mem/N39 ) );
  NOR2_X2 U3223 ( .A1(n6548), .A2(n3207), .ZN(\ex_mem/N45 ) );
  NOR2_X2 U3224 ( .A1(n6629), .A2(n3207), .ZN(\ex_mem/N141 ) );
  BUF_X4 U3225 ( .A(n3727), .Z(n3076) );
  INV_X4 U3226 ( .A(n3285), .ZN(n3280) );
  INV_X4 U3227 ( .A(n3288), .ZN(n3271) );
  INV_X4 U3228 ( .A(n3286), .ZN(n3277) );
  OAI21_X2 U3229 ( .B1(n6609), .B2(n3188), .A(n3872), .ZN(n2105) );
  OAI21_X2 U3230 ( .B1(n6629), .B2(n3188), .A(n3876), .ZN(n6770) );
  OAI21_X2 U3231 ( .B1(n6630), .B2(n3188), .A(n3877), .ZN(n6769) );
  OAI21_X2 U3232 ( .B1(n6631), .B2(n3188), .A(n3878), .ZN(n6768) );
  INV_X4 U3233 ( .A(n3286), .ZN(n3276) );
  OAI21_X2 U3234 ( .B1(n6633), .B2(n3188), .A(n3881), .ZN(n6766) );
  OAI21_X2 U3235 ( .B1(n6634), .B2(n3188), .A(n3882), .ZN(n6773) );
  OAI21_X2 U3236 ( .B1(n6635), .B2(n3188), .A(n3885), .ZN(n6777) );
  INV_X4 U3237 ( .A(n3287), .ZN(n3274) );
  OAI21_X2 U3238 ( .B1(n6636), .B2(n3188), .A(n3888), .ZN(n6775) );
  OAI21_X2 U3239 ( .B1(n6616), .B2(n3188), .A(n3890), .ZN(n2120) );
  INV_X4 U3240 ( .A(n3287), .ZN(n3275) );
  INV_X4 U3241 ( .A(n3292), .ZN(n3272) );
  OAI21_X2 U3242 ( .B1(n6598), .B2(n3188), .A(n5169), .ZN(n6772) );
  AOI21_X2 U3243 ( .B1(setInv_2), .B2(n3196), .A(n6391), .ZN(n6390) );
  INV_X4 U3244 ( .A(n3286), .ZN(n3278) );
  INV_X4 U3245 ( .A(n3288), .ZN(n3269) );
  INV_X4 U3246 ( .A(n3287), .ZN(n3273) );
  INV_X4 U3247 ( .A(n3288), .ZN(n3268) );
  NOR2_X2 U3248 ( .A1(n3926), .A2(n3211), .ZN(\ex_mem/N106 ) );
  NOR2_X2 U3249 ( .A1(n3934), .A2(n3208), .ZN(\ex_mem/N115 ) );
  NOR2_X2 U3250 ( .A1(n3941), .A2(n3209), .ZN(\ex_mem/N120 ) );
  NOR2_X2 U3251 ( .A1(n3949), .A2(n3210), .ZN(\ex_mem/N121 ) );
  NOR2_X2 U3252 ( .A1(n3957), .A2(n3211), .ZN(\ex_mem/N122 ) );
  NOR2_X2 U3253 ( .A1(n3965), .A2(n3208), .ZN(\ex_mem/N123 ) );
  NOR2_X2 U3254 ( .A1(n3973), .A2(n3211), .ZN(\ex_mem/N124 ) );
  NOR2_X2 U3255 ( .A1(n3978), .A2(n3208), .ZN(\ex_mem/N130 ) );
  AOI21_X2 U3256 ( .B1(n3171), .B2(regWrData[31]), .A(n4302), .ZN(n3978) );
  NOR2_X2 U3257 ( .A1(n3983), .A2(n3211), .ZN(\ex_mem/N103 ) );
  AOI211_X2 U3258 ( .C1(n3171), .C2(regWrData[4]), .A(n4208), .B(n4209), .ZN(
        n3983) );
  NOR2_X2 U3259 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  AOI21_X2 U3260 ( .B1(n3170), .B2(regWrData[2]), .A(n3999), .ZN(n4000) );
  AOI21_X2 U3261 ( .B1(n4005), .B2(n4176), .A(n3209), .ZN(\ex_mem/N100 ) );
  AOI21_X2 U3262 ( .B1(n3171), .B2(regWrData[1]), .A(n4004), .ZN(n4005) );
  NOR2_X2 U3263 ( .A1(n4008), .A2(n3211), .ZN(\ex_mem/N102 ) );
  AOI211_X2 U3264 ( .C1(n3171), .C2(regWrData[3]), .A(n4188), .B(n4192), .ZN(
        n4008) );
  AOI21_X2 U3265 ( .B1(n4014), .B2(n4379), .A(n3208), .ZN(\ex_mem/N105 ) );
  AOI21_X2 U3266 ( .B1(n3171), .B2(regWrData[6]), .A(n4013), .ZN(n4014) );
  NOR2_X2 U3267 ( .A1(n4017), .A2(n3211), .ZN(\ex_mem/N110 ) );
  NOR2_X2 U3268 ( .A1(n4024), .A2(n3211), .ZN(\ex_mem/N128 ) );
  NOR2_X2 U3269 ( .A1(n4034), .A2(n3211), .ZN(\ex_mem/N107 ) );
  AOI21_X2 U3270 ( .B1(n4038), .B2(n4314), .A(n3208), .ZN(\ex_mem/N111 ) );
  AOI21_X2 U3271 ( .B1(n3171), .B2(regWrData[12]), .A(n4037), .ZN(n4038) );
  AOI21_X2 U3272 ( .B1(n4044), .B2(n3093), .A(n3206), .ZN(\ex_mem/N112 ) );
  AOI21_X2 U3273 ( .B1(n3171), .B2(regWrData[13]), .A(n4043), .ZN(n4044) );
  NOR2_X2 U3274 ( .A1(n4051), .A2(n3211), .ZN(\ex_mem/N109 ) );
  NOR2_X2 U3275 ( .A1(n6510), .A2(n3211), .ZN(\ex_mem/N66 ) );
  NOR2_X2 U3276 ( .A1(n4060), .A2(n3211), .ZN(\ex_mem/N129 ) );
  NOR2_X2 U3277 ( .A1(n4067), .A2(n3211), .ZN(\ex_mem/N118 ) );
  NOR2_X2 U3278 ( .A1(n4072), .A2(n3210), .ZN(n2552) );
  NOR2_X2 U3279 ( .A1(n4079), .A2(n3211), .ZN(\ex_mem/N104 ) );
  AOI211_X2 U3280 ( .C1(n3171), .C2(regWrData[5]), .A(n3113), .B(n4078), .ZN(
        n4079) );
  AOI21_X2 U3281 ( .B1(n3171), .B2(regWrData[14]), .A(n4082), .ZN(n4084) );
  AOI21_X2 U3282 ( .B1(n4091), .B2(n4233), .A(n3208), .ZN(\ex_mem/N114 ) );
  AOI21_X2 U3283 ( .B1(n3170), .B2(regWrData[15]), .A(n4090), .ZN(n4091) );
  NOR2_X2 U3284 ( .A1(n4101), .A2(n3210), .ZN(\ex_mem/N116 ) );
  AOI21_X2 U3285 ( .B1(n3171), .B2(regWrData[17]), .A(n4395), .ZN(n4101) );
  NOR2_X2 U3286 ( .A1(n4110), .A2(n3210), .ZN(\ex_mem/N117 ) );
  NOR2_X2 U3287 ( .A1(n4118), .A2(n3210), .ZN(\ex_mem/N119 ) );
  NOR2_X2 U3288 ( .A1(n4125), .A2(n3210), .ZN(\ex_mem/N125 ) );
  NOR2_X2 U3289 ( .A1(n4134), .A2(n3210), .ZN(\ex_mem/N126 ) );
  NOR2_X2 U3290 ( .A1(n4144), .A2(n3210), .ZN(\ex_mem/N127 ) );
  NOR2_X2 U3291 ( .A1(n4742), .A2(n3210), .ZN(n2537) );
  NOR2_X2 U3292 ( .A1(n4550), .A2(n4549), .ZN(n4748) );
  NOR2_X2 U3293 ( .A1(n4750), .A2(n3210), .ZN(n2532) );
  NOR2_X2 U3294 ( .A1(n5179), .A2(n3210), .ZN(n2547) );
  NOR2_X2 U3295 ( .A1(n4822), .A2(n4821), .ZN(n4825) );
  NOR2_X2 U3296 ( .A1(n4826), .A2(n3210), .ZN(n2555) );
  NOR2_X2 U3297 ( .A1(n4897), .A2(n3210), .ZN(n2538) );
  NOR2_X2 U3298 ( .A1(n5178), .A2(n3210), .ZN(n2548) );
  NOR2_X2 U3299 ( .A1(n4907), .A2(n3209), .ZN(n2528) );
  NOR2_X2 U3300 ( .A1(n4908), .A2(n3209), .ZN(n2540) );
  NOR2_X2 U3301 ( .A1(n4909), .A2(n3209), .ZN(n2545) );
  NOR2_X2 U3302 ( .A1(n5181), .A2(n3209), .ZN(n2550) );
  NOR2_X2 U3303 ( .A1(n5799), .A2(n3209), .ZN(n2541) );
  NOR2_X2 U3304 ( .A1(n4910), .A2(n3209), .ZN(n2536) );
  AOI211_X2 U3305 ( .C1(n4921), .C2(n4920), .A(n4919), .B(n4918), .ZN(n4993)
         );
  NOR2_X2 U3306 ( .A1(n4994), .A2(n3209), .ZN(n2535) );
  NOR2_X2 U3307 ( .A1(n5092), .A2(n3209), .ZN(n2556) );
  NOR3_X2 U3308 ( .A1(n5095), .A2(n5094), .A3(n5093), .ZN(n5096) );
  OAI21_X2 U3309 ( .B1(n5072), .B2(n5071), .A(n5070), .ZN(n5077) );
  INV_X4 U3310 ( .A(n3291), .ZN(n3259) );
  NOR2_X2 U3311 ( .A1(n5098), .A2(n3209), .ZN(n2559) );
  NAND2_X2 U3312 ( .A1(n5135), .A2(n5134), .ZN(\ex_mem/N224 ) );
  AOI211_X2 U3313 ( .C1(n3129), .C2(n6005), .A(n5118), .B(n5117), .ZN(n5135)
         );
  NOR2_X2 U3314 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  NOR2_X2 U3315 ( .A1(n6513), .A2(n3209), .ZN(\ex_mem/N47 ) );
  NOR2_X2 U3316 ( .A1(n6515), .A2(n3209), .ZN(\ex_mem/N44 ) );
  NOR2_X2 U3317 ( .A1(n6516), .A2(n3209), .ZN(\ex_mem/N43 ) );
  NOR2_X2 U3318 ( .A1(n5136), .A2(n3208), .ZN(n2557) );
  NOR2_X2 U3319 ( .A1(n5137), .A2(n3208), .ZN(n2558) );
  INV_X4 U3320 ( .A(n3291), .ZN(n3260) );
  NOR2_X2 U3321 ( .A1(n5141), .A2(n3208), .ZN(n2534) );
  NOR2_X2 U3322 ( .A1(n5603), .A2(n3208), .ZN(n6734) );
  NOR2_X2 U3323 ( .A1(n6007), .A2(n3208), .ZN(n6733) );
  NOR2_X2 U3324 ( .A1(n6616), .A2(n3208), .ZN(\ex_mem/N131 ) );
  NOR2_X2 U3325 ( .A1(n6636), .A2(n3207), .ZN(\ex_mem/N132 ) );
  NOR2_X2 U3326 ( .A1(n6601), .A2(n3210), .ZN(\ex_mem/N133 ) );
  NOR2_X2 U3327 ( .A1(n6635), .A2(n3207), .ZN(\ex_mem/N134 ) );
  NOR2_X2 U3328 ( .A1(n6602), .A2(n3206), .ZN(\ex_mem/N135 ) );
  NOR2_X2 U3329 ( .A1(n6634), .A2(n3206), .ZN(\ex_mem/N136 ) );
  INV_X4 U3330 ( .A(n3291), .ZN(n3261) );
  NOR2_X2 U3331 ( .A1(n6633), .A2(n3206), .ZN(\ex_mem/N137 ) );
  NOR2_X2 U3332 ( .A1(n6632), .A2(n3207), .ZN(\ex_mem/N138 ) );
  NOR2_X2 U3333 ( .A1(n6631), .A2(n3207), .ZN(\ex_mem/N139 ) );
  NOR2_X2 U3334 ( .A1(n6630), .A2(n3210), .ZN(\ex_mem/N140 ) );
  NOR2_X2 U3335 ( .A1(n6607), .A2(n3208), .ZN(\ex_mem/N143 ) );
  NOR2_X2 U3336 ( .A1(n6604), .A2(n3207), .ZN(\ex_mem/N144 ) );
  NOR2_X2 U3337 ( .A1(n6608), .A2(n3207), .ZN(\ex_mem/N145 ) );
  NOR2_X2 U3338 ( .A1(n6609), .A2(n3207), .ZN(\ex_mem/N146 ) );
  INV_X4 U3339 ( .A(n3290), .ZN(n3262) );
  NOR2_X2 U3340 ( .A1(n6626), .A2(n3207), .ZN(\ex_mem/N149 ) );
  NOR2_X2 U3341 ( .A1(n6625), .A2(n3207), .ZN(\ex_mem/N150 ) );
  NOR2_X2 U3342 ( .A1(n6624), .A2(n3207), .ZN(\ex_mem/N151 ) );
  NOR2_X2 U3343 ( .A1(n6623), .A2(n3207), .ZN(\ex_mem/N152 ) );
  NOR2_X2 U3344 ( .A1(n6622), .A2(n3207), .ZN(\ex_mem/N153 ) );
  NOR2_X2 U3345 ( .A1(n6621), .A2(n3207), .ZN(\ex_mem/N154 ) );
  NOR2_X2 U3346 ( .A1(n6620), .A2(n3207), .ZN(\ex_mem/N155 ) );
  NOR2_X2 U3347 ( .A1(n6619), .A2(n3207), .ZN(\ex_mem/N156 ) );
  NOR2_X2 U3348 ( .A1(n6611), .A2(n3206), .ZN(\ex_mem/N157 ) );
  NOR2_X2 U3349 ( .A1(n6610), .A2(n3206), .ZN(\ex_mem/N158 ) );
  NOR2_X2 U3350 ( .A1(n6613), .A2(n3206), .ZN(\ex_mem/N159 ) );
  NOR2_X2 U3351 ( .A1(n6614), .A2(n3206), .ZN(\ex_mem/N160 ) );
  NOR2_X2 U3352 ( .A1(n6612), .A2(n3206), .ZN(\ex_mem/N161 ) );
  NOR2_X2 U3353 ( .A1(n6605), .A2(n3206), .ZN(\ex_mem/N162 ) );
  NOR2_X2 U3354 ( .A1(n5561), .A2(n3206), .ZN(n2542) );
  NOR2_X2 U3355 ( .A1(n5182), .A2(n3206), .ZN(n2551) );
  NOR2_X2 U3356 ( .A1(n5180), .A2(n3206), .ZN(n2546) );
  NOR2_X2 U3357 ( .A1(n5153), .A2(n3206), .ZN(n2539) );
  NOR2_X2 U3358 ( .A1(n5157), .A2(n3206), .ZN(n2554) );
  NOR2_X2 U3359 ( .A1(n5161), .A2(n3206), .ZN(n2553) );
  NOR2_X2 U3360 ( .A1(n5162), .A2(n3206), .ZN(n2531) );
  NOR2_X2 U3361 ( .A1(n5480), .A2(n3205), .ZN(n2533) );
  NOR2_X2 U3362 ( .A1(n5163), .A2(n3205), .ZN(n2544) );
  NOR2_X2 U3363 ( .A1(n5773), .A2(n3205), .ZN(n2530) );
  NOR2_X2 U3364 ( .A1(n6226), .A2(n3205), .ZN(\ex_mem/N240 ) );
  NOR2_X2 U3365 ( .A1(n5164), .A2(n3196), .ZN(n6765) );
  NOR2_X2 U3366 ( .A1(n6368), .A2(n2635), .ZN(n5164) );
  NOR2_X2 U3367 ( .A1(n6598), .A2(n3205), .ZN(\ex_mem/N229 ) );
  NOR2_X2 U3368 ( .A1(n6253), .A2(n3205), .ZN(\ex_mem/N230 ) );
  NOR2_X2 U3369 ( .A1(n6235), .A2(n3205), .ZN(\ex_mem/N231 ) );
  NOR2_X2 U3370 ( .A1(n6525), .A2(n3205), .ZN(\ex_mem/N233 ) );
  NOR2_X2 U3371 ( .A1(n6526), .A2(n3205), .ZN(\ex_mem/N234 ) );
  NOR2_X2 U3372 ( .A1(n6597), .A2(n3205), .ZN(\ex_mem/N235 ) );
  NOR2_X2 U3373 ( .A1(n6524), .A2(n3205), .ZN(\ex_mem/N236 ) );
  NOR2_X2 U3374 ( .A1(n3208), .A2(n2878), .ZN(\ex_mem/N237 ) );
  INV_X4 U3375 ( .A(n3289), .ZN(n3265) );
  NOR2_X2 U3376 ( .A1(n6233), .A2(n3205), .ZN(\ex_mem/N239 ) );
  NOR2_X2 U3377 ( .A1(n6368), .A2(n3196), .ZN(\id_ex/N42 ) );
  NOR2_X2 U3378 ( .A1(n2786), .A2(n3205), .ZN(\ex_mem/N241 ) );
  INV_X4 U3379 ( .A(n3290), .ZN(n3263) );
  NOR2_X2 U3380 ( .A1(n2593), .A2(n3204), .ZN(\ex_mem/N246 ) );
  INV_X4 U3381 ( .A(n3292), .ZN(n3257) );
  NOR2_X2 U3382 ( .A1(n2782), .A2(n3204), .ZN(\ex_mem/N247 ) );
  NOR2_X2 U3383 ( .A1(n5166), .A2(n3204), .ZN(\ex_mem/N99 ) );
  AOI21_X2 U3384 ( .B1(n3171), .B2(regWrData[0]), .A(n5165), .ZN(n5166) );
  INV_X4 U3385 ( .A(n3290), .ZN(n3264) );
  NAND2_X2 U3386 ( .A1(n6490), .A2(n6386), .ZN(n5167) );
  INV_X4 U3387 ( .A(n3292), .ZN(n3256) );
  NOR2_X2 U3388 ( .A1(n2781), .A2(n3204), .ZN(\ex_mem/N243 ) );
  INV_X4 U3389 ( .A(n3289), .ZN(n3266) );
  INV_X4 U3390 ( .A(n3289), .ZN(n3267) );
  NOR2_X2 U3391 ( .A1(1'b0), .A2(n3196), .ZN(\id_ex/N44 ) );
  NOR2_X2 U3392 ( .A1(n3196), .A2(n6552), .ZN(n6112) );
  NOR2_X2 U3393 ( .A1(n3197), .A2(n6551), .ZN(n6113) );
  NOR2_X2 U3394 ( .A1(n3196), .A2(n6550), .ZN(n6114) );
  NOR2_X2 U3395 ( .A1(n3196), .A2(n6549), .ZN(n6115) );
  NOR2_X2 U3396 ( .A1(n3197), .A2(n6527), .ZN(n6116) );
  NOR2_X2 U3397 ( .A1(n3197), .A2(n6553), .ZN(n6134) );
  NOR2_X2 U3398 ( .A1(n3197), .A2(n2832), .ZN(n6118) );
  NOR2_X2 U3399 ( .A1(n3197), .A2(n2835), .ZN(n6119) );
  NOR2_X2 U3400 ( .A1(n3197), .A2(n2834), .ZN(n6120) );
  NOR2_X2 U3401 ( .A1(n3197), .A2(n2709), .ZN(n6127) );
  NOR2_X2 U3402 ( .A1(n3197), .A2(n2831), .ZN(n6121) );
  NOR2_X2 U3403 ( .A1(n6589), .A2(n3196), .ZN(\id_ex/N31 ) );
  NOR2_X2 U3404 ( .A1(n3197), .A2(n6587), .ZN(n6128) );
  NOR2_X2 U3405 ( .A1(n6590), .A2(n3196), .ZN(\id_ex/N33 ) );
  NOR2_X2 U3406 ( .A1(n6486), .A2(n3196), .ZN(\id_ex/N38 ) );
  INV_X4 U3407 ( .A(n3849), .ZN(n6131) );
  NOR2_X2 U3408 ( .A1(n3197), .A2(n6592), .ZN(n6125) );
  NOR2_X2 U3409 ( .A1(n3197), .A2(n6593), .ZN(n6126) );
  NOR2_X2 U3410 ( .A1(n2629), .A2(n3204), .ZN(\ex_mem/N245 ) );
  NOR2_X2 U3411 ( .A1(n2628), .A2(n3204), .ZN(\ex_mem/N244 ) );
  NOR3_X2 U3412 ( .A1(n5206), .A2(n5205), .A3(n5204), .ZN(\ex_mem/N232 ) );
  INV_X4 U3413 ( .A(n3299), .ZN(n3248) );
  AOI211_X2 U3414 ( .C1(n5216), .C2(n5215), .A(n5214), .B(n5213), .ZN(n5232)
         );
  NOR3_X2 U3415 ( .A1(n5318), .A2(n5317), .A3(n5316), .ZN(n5319) );
  OAI21_X2 U3416 ( .B1(n5256), .B2(n3063), .A(n5255), .ZN(n5259) );
  NOR2_X2 U3417 ( .A1(n6529), .A2(n3204), .ZN(\ex_mem/N65 ) );
  NOR2_X2 U3418 ( .A1(n6530), .A2(n3204), .ZN(\ex_mem/N64 ) );
  NOR2_X2 U3419 ( .A1(n6531), .A2(n3204), .ZN(\ex_mem/N63 ) );
  NOR2_X2 U3420 ( .A1(n6532), .A2(n3204), .ZN(\ex_mem/N62 ) );
  NOR2_X2 U3421 ( .A1(n6533), .A2(n3204), .ZN(\ex_mem/N61 ) );
  NOR2_X2 U3422 ( .A1(n6534), .A2(n3204), .ZN(\ex_mem/N60 ) );
  NOR2_X2 U3423 ( .A1(n6535), .A2(n3208), .ZN(\ex_mem/N59 ) );
  NOR2_X2 U3424 ( .A1(n6536), .A2(n3208), .ZN(\ex_mem/N58 ) );
  NOR2_X2 U3425 ( .A1(n6537), .A2(n3208), .ZN(\ex_mem/N57 ) );
  NOR2_X2 U3426 ( .A1(n6538), .A2(n3208), .ZN(\ex_mem/N56 ) );
  NOR2_X2 U3427 ( .A1(n6539), .A2(n3208), .ZN(\ex_mem/N55 ) );
  NOR2_X2 U3428 ( .A1(n6540), .A2(n3204), .ZN(\ex_mem/N54 ) );
  NOR2_X2 U3429 ( .A1(n6541), .A2(n3208), .ZN(\ex_mem/N53 ) );
  NOR2_X2 U3430 ( .A1(n6544), .A2(n3208), .ZN(\ex_mem/N50 ) );
  NOR2_X2 U3431 ( .A1(n6545), .A2(n3208), .ZN(\ex_mem/N49 ) );
  NOR2_X2 U3432 ( .A1(n6546), .A2(n3208), .ZN(\ex_mem/N48 ) );
  INV_X4 U3433 ( .A(n3293), .ZN(n3250) );
  AOI211_X2 U3434 ( .C1(n5352), .C2(n5351), .A(n5350), .B(n5349), .ZN(n5367)
         );
  AOI211_X2 U3435 ( .C1(n5377), .C2(n5383), .A(n5382), .B(n5381), .ZN(n5391)
         );
  AOI211_X2 U3436 ( .C1(n5428), .C2(n5427), .A(n5426), .B(n5425), .ZN(n5457)
         );
  NOR2_X2 U3437 ( .A1(n5497), .A2(n5496), .ZN(n5522) );
  AOI211_X2 U3438 ( .C1(n5560), .C2(n5559), .A(n5558), .B(n5557), .ZN(n5568)
         );
  AOI211_X2 U3439 ( .C1(n3156), .C2(n5585), .A(n5584), .B(n5583), .ZN(n5590)
         );
  AOI211_X2 U3440 ( .C1(n5600), .C2(n5599), .A(n5598), .B(n5597), .ZN(n5609)
         );
  NOR2_X2 U3441 ( .A1(n5605), .A2(n5604), .ZN(n5607) );
  NOR2_X2 U3442 ( .A1(n5637), .A2(n5636), .ZN(n5660) );
  NOR2_X2 U3443 ( .A1(n5655), .A2(n5654), .ZN(n5659) );
  INV_X4 U3444 ( .A(n3293), .ZN(n3251) );
  AOI211_X2 U3445 ( .C1(n5670), .C2(n5676), .A(n5675), .B(n5674), .ZN(n5685)
         );
  NOR3_X2 U3446 ( .A1(n5776), .A2(n5775), .A3(n5774), .ZN(n5777) );
  AOI211_X2 U3447 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5813), .ZN(n5830)
         );
  NAND2_X2 U3448 ( .A1(n5873), .A2(n5874), .ZN(\ex_mem/N219 ) );
  AOI211_X2 U3449 ( .C1(n6005), .C2(n5995), .A(n5863), .B(n5862), .ZN(n5874)
         );
  NOR2_X2 U3450 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  OAI21_X2 U3451 ( .B1(n5861), .B2(n5860), .A(n5859), .ZN(n5863) );
  AOI211_X2 U3452 ( .C1(n5884), .C2(n5883), .A(n5882), .B(n5881), .ZN(n5902)
         );
  AOI211_X2 U3453 ( .C1(n5913), .C2(n5912), .A(n5911), .B(n5910), .ZN(n5936)
         );
  NOR2_X2 U3454 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  INV_X4 U3455 ( .A(n3293), .ZN(n3252) );
  AOI211_X2 U3456 ( .C1(n5616), .C2(n5622), .A(n5621), .B(n5620), .ZN(n5630)
         );
  NOR2_X2 U3457 ( .A1(n2843), .A2(n2625), .ZN(n5359) );
  OAI21_X2 U3458 ( .B1(n5616), .B2(n3229), .A(n6008), .ZN(n5617) );
  NOR2_X2 U3459 ( .A1(n2625), .A2(n5499), .ZN(n5502) );
  NOR2_X2 U3460 ( .A1(n5354), .A2(n2625), .ZN(n4829) );
  NAND4_X2 U3461 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n2584)
         );
  NAND4_X2 U3462 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6096)
         );
  OAI222_X2 U3463 ( .A1(n6318), .A2(n4162), .B1(n3124), .B2(n3152), .C1(n3154), 
        .C2(n2988), .ZN(regWrData[19]) );
  NAND2_X2 U3464 ( .A1(n5368), .A2(n3130), .ZN(n3132) );
  XNOR2_X1 U3465 ( .A(n5021), .B(n5908), .ZN(n5914) );
  OAI211_X4 U3466 ( .C1(n4978), .C2(n3157), .A(n5266), .B(n4977), .ZN(n5087)
         );
  NAND2_X4 U3467 ( .A1(n5651), .A2(n5638), .ZN(n4599) );
  NAND2_X2 U3468 ( .A1(n5011), .A2(n5885), .ZN(n5920) );
  OAI21_X2 U3469 ( .B1(n4841), .B2(n5011), .A(n5885), .ZN(n5221) );
  INV_X2 U3470 ( .A(n4790), .ZN(n5179) );
  INV_X2 U3471 ( .A(n5864), .ZN(n5867) );
  AOI22_X1 U3472 ( .A1(n3225), .A2(n5825), .B1(n5948), .B2(n5864), .ZN(n5828)
         );
  OAI21_X4 U3473 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(n6032) );
  NAND2_X1 U3474 ( .A1(n5080), .A2(n6002), .ZN(n4462) );
  NOR4_X2 U3475 ( .A1(n4449), .A2(n5492), .A3(n6603), .A4(n3061), .ZN(n4435)
         );
  XNOR2_X2 U3476 ( .A(n4883), .B(n4566), .ZN(n2587) );
  INV_X4 U3477 ( .A(n2587), .ZN(n4895) );
  OAI211_X2 U3478 ( .C1(n4570), .C2(n4803), .A(n3059), .B(n4673), .ZN(n2588)
         );
  INV_X4 U3479 ( .A(n4883), .ZN(n4880) );
  OAI211_X2 U3480 ( .C1(n4570), .C2(n4803), .A(n3059), .B(n4673), .ZN(n5044)
         );
  INV_X2 U3481 ( .A(n5044), .ZN(n5845) );
  NAND2_X4 U3482 ( .A1(n5196), .A2(n3041), .ZN(n4735) );
  INV_X4 U3483 ( .A(n4935), .ZN(n4911) );
  AOI21_X1 U3484 ( .B1(n4917), .B2(n3226), .A(n4935), .ZN(n4918) );
  INV_X4 U3485 ( .A(n5616), .ZN(n2589) );
  OAI211_X2 U3486 ( .C1(n4169), .C2(n4168), .A(n4167), .B(n4166), .ZN(n5610)
         );
  NOR2_X2 U3487 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  XNOR2_X1 U3488 ( .A(n3706), .B(n2810), .ZN(n3707) );
  NAND3_X2 U3489 ( .A1(n4089), .A2(n4238), .A3(n4088), .ZN(regWrData[15]) );
  NOR2_X2 U3490 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  OAI221_X1 U3491 ( .B1(n6586), .B2(n3155), .C1(n4552), .C2(n3184), .A(n4551), 
        .ZN(n4790) );
  NAND3_X2 U3492 ( .A1(n4687), .A2(n4686), .A3(n4685), .ZN(n5451) );
  XOR2_X2 U3493 ( .A(n4773), .B(n3221), .Z(n2724) );
  OAI21_X1 U3494 ( .B1(n2589), .B2(n5277), .A(n5276), .ZN(n5278) );
  AND2_X2 U3495 ( .A1(n3156), .A2(n2589), .ZN(n2908) );
  INV_X1 U3496 ( .A(n5610), .ZN(n5616) );
  NAND2_X2 U3497 ( .A1(n5707), .A2(n4575), .ZN(n5647) );
  INV_X4 U3498 ( .A(n5958), .ZN(n5959) );
  NAND2_X2 U3499 ( .A1(n5959), .A2(n5960), .ZN(n5967) );
  NAND2_X1 U3500 ( .A1(n5960), .A2(n5959), .ZN(n3128) );
  INV_X1 U3501 ( .A(n5397), .ZN(n2591) );
  NAND2_X4 U3502 ( .A1(n4661), .A2(n5531), .ZN(n5398) );
  NAND3_X4 U3503 ( .A1(n4226), .A2(n4225), .A3(n4224), .ZN(n5661) );
  INV_X8 U3504 ( .A(n3060), .ZN(n3061) );
  NAND2_X2 U3505 ( .A1(n3214), .A2(n2872), .ZN(n2592) );
  INV_X4 U3506 ( .A(n2625), .ZN(n5695) );
  INV_X4 U3507 ( .A(n3214), .ZN(n3209) );
  INV_X4 U3508 ( .A(n3214), .ZN(n3208) );
  NAND3_X2 U3509 ( .A1(n6448), .A2(n3684), .A3(n3683), .ZN(n3816) );
  INV_X4 U3510 ( .A(n3200), .ZN(n3195) );
  INV_X4 U3511 ( .A(\mem_wb/N41 ), .ZN(n3291) );
  INV_X4 U3512 ( .A(n2779), .ZN(n5947) );
  INV_X8 U3513 ( .A(n4525), .ZN(n3174) );
  INV_X16 U3514 ( .A(n3199), .ZN(n3197) );
  INV_X4 U3515 ( .A(n2778), .ZN(n6029) );
  INV_X4 U3516 ( .A(n2776), .ZN(n3231) );
  INV_X8 U3517 ( .A(n3174), .ZN(n3172) );
  INV_X8 U3518 ( .A(n3173), .ZN(n3075) );
  INV_X1 U3519 ( .A(n3201), .ZN(n3212) );
  INV_X4 U3520 ( .A(n3214), .ZN(n3204) );
  INV_X4 U3521 ( .A(n3214), .ZN(n3205) );
  INV_X8 U3522 ( .A(n3195), .ZN(n3193) );
  INV_X4 U3523 ( .A(\mem_wb/N41 ), .ZN(n3288) );
  INV_X4 U3524 ( .A(n3292), .ZN(n3253) );
  INV_X4 U3525 ( .A(n3288), .ZN(n3258) );
  INV_X4 U3526 ( .A(n3291), .ZN(n3270) );
  OR2_X4 U3527 ( .A1(n6587), .A2(op0_1), .ZN(n2603) );
  AND2_X4 U3528 ( .A1(n5670), .A2(n3157), .ZN(n2605) );
  INV_X4 U3529 ( .A(n6008), .ZN(n3228) );
  AND2_X4 U3530 ( .A1(n5940), .A2(n4445), .ZN(n2620) );
  AND2_X4 U3531 ( .A1(n6231), .A2(n6254), .ZN(n2723) );
  INV_X4 U3532 ( .A(n2844), .ZN(n3224) );
  AND2_X4 U3533 ( .A1(n2708), .A2(n6618), .ZN(n2621) );
  INV_X4 U3534 ( .A(n2789), .ZN(n3240) );
  INV_X4 U3535 ( .A(n2789), .ZN(n3239) );
  XNOR2_X2 U3536 ( .A(n5718), .B(n6088), .ZN(n2622) );
  NAND2_X1 U3537 ( .A1(n6037), .A2(n5610), .ZN(n6036) );
  AND2_X4 U3538 ( .A1(n3213), .A2(n3282), .ZN(n2623) );
  INV_X8 U3539 ( .A(n3144), .ZN(n3145) );
  INV_X2 U3540 ( .A(n3203), .ZN(n3201) );
  INV_X4 U3541 ( .A(n3202), .ZN(n3214) );
  INV_X4 U3542 ( .A(n3156), .ZN(n3157) );
  INV_X8 U3543 ( .A(n5704), .ZN(n3156) );
  INV_X4 U3544 ( .A(n3757), .ZN(n3659) );
  INV_X4 U3545 ( .A(n3816), .ZN(n3164) );
  NAND2_X2 U3546 ( .A1(n5616), .A2(n6037), .ZN(n2625) );
  NAND2_X2 U3547 ( .A1(n2621), .A2(n6015), .ZN(n2626) );
  NAND2_X2 U3548 ( .A1(n2621), .A2(n5969), .ZN(n2627) );
  INV_X4 U3549 ( .A(\mem_wb/N41 ), .ZN(n3294) );
  INV_X4 U3550 ( .A(n3292), .ZN(n3254) );
  INV_X4 U3551 ( .A(n3292), .ZN(n3255) );
  INV_X4 U3552 ( .A(n3293), .ZN(n3249) );
  NAND2_X1 U3553 ( .A1(n4083), .A2(n3159), .ZN(n4329) );
  AND2_X4 U3554 ( .A1(n6254), .A2(n2888), .ZN(n2680) );
  AND2_X2 U3555 ( .A1(n3156), .A2(n5670), .ZN(n2685) );
  INV_X4 U3556 ( .A(n4162), .ZN(n4139) );
  AND2_X4 U3557 ( .A1(n3428), .A2(n3426), .ZN(n2692) );
  AND2_X2 U3558 ( .A1(n6600), .A2(n6603), .ZN(n2706) );
  INV_X16 U3559 ( .A(n3179), .ZN(n3177) );
  INV_X16 U3560 ( .A(n3179), .ZN(n3178) );
  AND3_X4 U3561 ( .A1(n6100), .A2(n6600), .A3(n2602), .ZN(n2708) );
  AND2_X4 U3562 ( .A1(n3577), .A2(n3405), .ZN(n2711) );
  INV_X4 U3563 ( .A(n3213), .ZN(n3207) );
  INV_X4 U3564 ( .A(n3201), .ZN(n3213) );
  INV_X4 U3565 ( .A(n3213), .ZN(n3210) );
  INV_X4 U3566 ( .A(n3213), .ZN(n3206) );
  AND2_X4 U3567 ( .A1(n5858), .A2(n5009), .ZN(n2714) );
  INV_X4 U3568 ( .A(n3220), .ZN(n3219) );
  INV_X4 U3569 ( .A(n5719), .ZN(n3220) );
  AND2_X4 U3570 ( .A1(n6225), .A2(n2664), .ZN(n2715) );
  AND2_X4 U3571 ( .A1(n2664), .A2(n2601), .ZN(n2717) );
  NAND3_X2 U3572 ( .A1(n6100), .A2(n6618), .A3(n2663), .ZN(n2718) );
  AND2_X4 U3573 ( .A1(n5885), .A2(n5922), .ZN(n2720) );
  XOR2_X2 U3574 ( .A(iAddr[3]), .B(iAddr[2]), .Z(n2721) );
  NAND3_X2 U3575 ( .A1(n2706), .A2(n6100), .A3(n4545), .ZN(n6008) );
  INV_X4 U3576 ( .A(n3054), .ZN(n3055) );
  INV_X1 U3577 ( .A(n3145), .ZN(n4001) );
  INV_X4 U3578 ( .A(n3199), .ZN(n3198) );
  AND2_X4 U3579 ( .A1(n3795), .A2(n3794), .ZN(n2760) );
  AND2_X4 U3580 ( .A1(n3214), .A2(n5322), .ZN(n2761) );
  AND2_X4 U3581 ( .A1(n3194), .A2(n2974), .ZN(n2762) );
  AND2_X4 U3582 ( .A1(n3194), .A2(n2973), .ZN(n2763) );
  AND2_X4 U3583 ( .A1(n3194), .A2(n2972), .ZN(n2764) );
  INV_X4 U3584 ( .A(n3816), .ZN(n3166) );
  INV_X4 U3585 ( .A(n3816), .ZN(n3165) );
  NAND3_X2 U3586 ( .A1(n2708), .A2(n6617), .A3(n2595), .ZN(n2776) );
  NAND2_X2 U3587 ( .A1(n5616), .A2(n6040), .ZN(n2777) );
  INV_X4 U3588 ( .A(n3757), .ZN(n3161) );
  NAND2_X2 U3589 ( .A1(n4730), .A2(n6015), .ZN(n2778) );
  NAND2_X2 U3590 ( .A1(n4730), .A2(n5969), .ZN(n2779) );
  INV_X4 U3591 ( .A(\mem_wb/N41 ), .ZN(n3299) );
  INV_X4 U3592 ( .A(\mem_wb/N41 ), .ZN(n3293) );
  INV_X4 U3593 ( .A(\mem_wb/N41 ), .ZN(n3292) );
  INV_X4 U3594 ( .A(n4136), .ZN(n3149) );
  INV_X8 U3595 ( .A(n3149), .ZN(n3150) );
  NAND3_X2 U3596 ( .A1(n3216), .A2(n4462), .A3(n4461), .ZN(n6017) );
  INV_X4 U3597 ( .A(n6017), .ZN(n6019) );
  AND2_X4 U3598 ( .A1(n6386), .A2(n6413), .ZN(n2788) );
  AND2_X4 U3599 ( .A1(n6230), .A2(n2601), .ZN(n2789) );
  OR3_X4 U3600 ( .A1(n3087), .A2(n6329), .A3(n3244), .ZN(n2790) );
  INV_X4 U3601 ( .A(n5661), .ZN(n5670) );
  AND2_X4 U3602 ( .A1(n5670), .A2(n5261), .ZN(n2836) );
  INV_X4 U3603 ( .A(n5490), .ZN(n5492) );
  AND4_X4 U3604 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n2842)
         );
  AND3_X4 U3605 ( .A1(n4740), .A2(n4984), .A3(n4739), .ZN(n2843) );
  INV_X4 U3606 ( .A(n3117), .ZN(n3112) );
  AND3_X4 U3607 ( .A1(n6100), .A2(n2595), .A3(n2706), .ZN(n2844) );
  INV_X4 U3608 ( .A(n5914), .ZN(n5928) );
  XOR2_X2 U3609 ( .A(n6202), .B(n6279), .Z(n2847) );
  AND2_X4 U3610 ( .A1(n5036), .A2(n3106), .ZN(n2849) );
  AND2_X4 U3611 ( .A1(n3436), .A2(n3606), .ZN(n2851) );
  AND2_X4 U3612 ( .A1(n3156), .A2(n3110), .ZN(n2853) );
  INV_X4 U3613 ( .A(n5651), .ZN(n4598) );
  AND2_X4 U3614 ( .A1(n3598), .A2(n3597), .ZN(n2857) );
  XOR2_X2 U3615 ( .A(n6221), .B(n6261), .Z(n2870) );
  OR2_X4 U3616 ( .A1(n5354), .A2(n5510), .ZN(n2875) );
  AND2_X4 U3617 ( .A1(n3768), .A2(iAddr[13]), .ZN(n2876) );
  OR2_X4 U3618 ( .A1(n3243), .A2(n6636), .ZN(n2877) );
  INV_X4 U3619 ( .A(n2717), .ZN(n3242) );
  INV_X4 U3620 ( .A(n2717), .ZN(n3241) );
  OR2_X4 U3621 ( .A1(n6223), .A2(n3757), .ZN(n2879) );
  OR2_X4 U3622 ( .A1(n6162), .A2(n3757), .ZN(n2880) );
  AND3_X4 U3623 ( .A1(n3427), .A2(n3426), .A3(n3425), .ZN(n2881) );
  INV_X4 U3624 ( .A(n3195), .ZN(n3191) );
  INV_X4 U3625 ( .A(n3195), .ZN(n3192) );
  INV_X4 U3626 ( .A(n3198), .ZN(n3188) );
  AND2_X4 U3627 ( .A1(n4355), .A2(\wb/dsize_reg/z2 [31]), .ZN(n2887) );
  OR2_X4 U3628 ( .A1(reg31Val_3[0]), .A2(n2840), .ZN(n2890) );
  AND2_X4 U3629 ( .A1(reg31Val_0[31]), .A2(n3233), .ZN(n2891) );
  NAND2_X2 U3630 ( .A1(n4164), .A2(n4163), .ZN(n4622) );
  INV_X4 U3631 ( .A(n4622), .ZN(n4165) );
  INV_X16 U3632 ( .A(n3153), .ZN(n3154) );
  INV_X8 U3633 ( .A(n4343), .ZN(n3153) );
  AND2_X4 U3634 ( .A1(n3465), .A2(n3464), .ZN(n2894) );
  AND2_X4 U3635 ( .A1(n5886), .A2(n4769), .ZN(n2895) );
  AND2_X4 U3636 ( .A1(n3512), .A2(n3511), .ZN(n2897) );
  INV_X4 U3637 ( .A(n5941), .ZN(n3068) );
  NAND2_X2 U3638 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  OR2_X4 U3639 ( .A1(n4934), .A2(n2625), .ZN(n2900) );
  INV_X4 U3640 ( .A(n3762), .ZN(n3766) );
  INV_X4 U3641 ( .A(n3064), .ZN(n3065) );
  OR2_X4 U3642 ( .A1(n6196), .A2(n6188), .ZN(n2904) );
  AND2_X4 U3643 ( .A1(n5514), .A2(n5261), .ZN(n2905) );
  AND2_X4 U3644 ( .A1(n3740), .A2(n3739), .ZN(n2906) );
  AND2_X4 U3645 ( .A1(n3744), .A2(n3743), .ZN(n2907) );
  AND2_X4 U3646 ( .A1(n5327), .A2(n5326), .ZN(n2923) );
  INV_X4 U3647 ( .A(n3228), .ZN(n3227) );
  INV_X4 U3648 ( .A(n3228), .ZN(n3226) );
  OR2_X4 U3649 ( .A1(n6221), .A2(n6261), .ZN(n2954) );
  AND2_X4 U3650 ( .A1(n3194), .A2(n2661), .ZN(n2960) );
  NAND2_X2 U3651 ( .A1(n6493), .A2(n6370), .ZN(n6400) );
  NAND3_X2 U3652 ( .A1(n5130), .A2(n5129), .A3(n5128), .ZN(n5623) );
  OAI211_X2 U3653 ( .C1(n6044), .C2(n6040), .A(n5300), .B(n5299), .ZN(n5625)
         );
  AND2_X4 U3654 ( .A1(n3194), .A2(n2975), .ZN(n2981) );
  INV_X4 U3655 ( .A(n3759), .ZN(n3163) );
  INV_X4 U3656 ( .A(n3759), .ZN(n3162) );
  INV_X4 U3657 ( .A(n2715), .ZN(n3238) );
  INV_X4 U3658 ( .A(n2715), .ZN(n3237) );
  AND2_X4 U3659 ( .A1(n3780), .A2(n3781), .ZN(n2984) );
  AND2_X4 U3660 ( .A1(n5726), .A2(n5725), .ZN(n2990) );
  NAND2_X2 U3661 ( .A1(n5244), .A2(n5469), .ZN(n5058) );
  OR2_X4 U3662 ( .A1(n4285), .A2(n3245), .ZN(n2993) );
  AND2_X4 U3663 ( .A1(n4596), .A2(n5397), .ZN(n2994) );
  AND2_X4 U3664 ( .A1(n4036), .A2(n4320), .ZN(n2997) );
  INV_X4 U3665 ( .A(n6615), .ZN(n3245) );
  NAND3_X2 U3666 ( .A1(n6450), .A2(n6492), .A3(n6493), .ZN(n3028) );
  AND2_X4 U3667 ( .A1(n4589), .A2(n4588), .ZN(n3030) );
  INV_X4 U3668 ( .A(n2592), .ZN(n3225) );
  AND2_X4 U3669 ( .A1(n5417), .A2(n5418), .ZN(n3033) );
  INV_X4 U3670 ( .A(n3104), .ZN(n4473) );
  INV_X4 U3671 ( .A(n4069), .ZN(n3183) );
  INV_X4 U3672 ( .A(n4069), .ZN(n3182) );
  INV_X4 U3673 ( .A(n2718), .ZN(n6005) );
  INV_X4 U3674 ( .A(n5368), .ZN(n5377) );
  OAI21_X2 U3675 ( .B1(n4353), .B2(n4352), .A(n4351), .ZN(n5368) );
  INV_X4 U3676 ( .A(n3212), .ZN(n3211) );
  INV_X4 U3677 ( .A(n3231), .ZN(n3230) );
  INV_X4 U3678 ( .A(n3231), .ZN(n3229) );
  OR3_X4 U3679 ( .A1(n3196), .A2(n3821), .A3(n3820), .ZN(n3042) );
  INV_X8 U3680 ( .A(n3158), .ZN(n3159) );
  OR2_X4 U3681 ( .A1(n3197), .A2(rs1[3]), .ZN(n3043) );
  AND2_X4 U3682 ( .A1(n3197), .A2(n2866), .ZN(n3044) );
  AND2_X4 U3683 ( .A1(n3197), .A2(n2860), .ZN(n3045) );
  AND2_X4 U3684 ( .A1(n3197), .A2(n2862), .ZN(n3046) );
  AND2_X4 U3685 ( .A1(n3197), .A2(n2868), .ZN(n3047) );
  AND2_X4 U3686 ( .A1(n3197), .A2(n2873), .ZN(n3048) );
  AND2_X4 U3687 ( .A1(n3197), .A2(n2716), .ZN(n3049) );
  AND2_X4 U3688 ( .A1(n3197), .A2(n2863), .ZN(n3050) );
  AND2_X4 U3689 ( .A1(n3197), .A2(n2865), .ZN(n3051) );
  OR2_X4 U3690 ( .A1(n3197), .A2(n6487), .ZN(n3052) );
  AND2_X4 U3691 ( .A1(n3198), .A2(n2867), .ZN(n3053) );
  INV_X4 U3692 ( .A(\mem_wb/N41 ), .ZN(n3284) );
  INV_X4 U3693 ( .A(n3294), .ZN(n3246) );
  INV_X4 U3694 ( .A(n3292), .ZN(n3247) );
  INV_X4 U3695 ( .A(n3285), .ZN(n3279) );
  NOR2_X2 U3696 ( .A1(n4752), .A2(n5510), .ZN(n4757) );
  NOR2_X2 U3697 ( .A1(n2843), .A2(n5510), .ZN(n4868) );
  NOR2_X2 U3698 ( .A1(n5437), .A2(n5510), .ZN(n5441) );
  OAI221_X2 U3699 ( .B1(n5357), .B2(n5510), .C1(n2843), .C2(n6036), .A(n4741), 
        .ZN(n5385) );
  INV_X4 U3700 ( .A(n5510), .ZN(n5505) );
  NAND2_X2 U3702 ( .A1(n4333), .A2(n4332), .ZN(n4334) );
  NOR2_X2 U3703 ( .A1(n6305), .A2(n3091), .ZN(n4332) );
  INV_X2 U3704 ( .A(n5571), .ZN(n5579) );
  INV_X2 U3705 ( .A(n5988), .ZN(n5376) );
  NAND3_X2 U3706 ( .A1(reg31Val_0[7]), .A2(n3167), .A3(n3232), .ZN(n4249) );
  INV_X4 U3707 ( .A(n6615), .ZN(n3244) );
  OAI222_X2 U3708 ( .A1(n6304), .A2(n4162), .B1(n2699), .B2(n3152), .C1(n3154), 
        .C2(n2927), .ZN(regWrData[20]) );
  INV_X16 U3709 ( .A(n3151), .ZN(n3152) );
  INV_X4 U3710 ( .A(n6312), .ZN(n3054) );
  OAI222_X2 U3711 ( .A1(n6307), .A2(n4162), .B1(n2665), .B2(n3152), .C1(n3154), 
        .C2(n2976), .ZN(regWrData[26]) );
  NOR2_X2 U3712 ( .A1(n5410), .A2(n5226), .ZN(n5176) );
  AOI21_X2 U3713 ( .B1(n4308), .B2(n3180), .A(n4307), .ZN(n4309) );
  INV_X4 U3714 ( .A(n3180), .ZN(n3105) );
  NOR3_X2 U3715 ( .A1(n3180), .A2(n3145), .A3(n2992), .ZN(n4190) );
  INV_X16 U3716 ( .A(n3180), .ZN(n3176) );
  INV_X2 U3717 ( .A(regWrData[26]), .ZN(n4708) );
  INV_X2 U3718 ( .A(regWrData[19]), .ZN(n4071) );
  NAND2_X4 U3719 ( .A1(n3067), .A2(n3158), .ZN(n4525) );
  NAND4_X1 U3720 ( .A1(n3243), .A2(n4249), .A3(n4248), .A4(n4247), .ZN(n4260)
         );
  AOI21_X2 U3721 ( .B1(n4845), .B2(n4844), .A(n4843), .ZN(n4848) );
  INV_X4 U3722 ( .A(regWrData[7]), .ZN(n4586) );
  OAI222_X2 U3723 ( .A1(n6302), .A2(n4162), .B1(n2701), .B2(n3152), .C1(n3154), 
        .C2(n2922), .ZN(regWrData[18]) );
  INV_X1 U3724 ( .A(n5465), .ZN(n5477) );
  INV_X1 U3725 ( .A(n5444), .ZN(n5180) );
  AOI22_X1 U3726 ( .A1(n3225), .A2(n5444), .B1(n5947), .B2(n5864), .ZN(n5455)
         );
  INV_X1 U3727 ( .A(n5963), .ZN(n4776) );
  INV_X4 U3728 ( .A(n5737), .ZN(n3056) );
  INV_X4 U3729 ( .A(n5033), .ZN(n3058) );
  INV_X1 U3730 ( .A(n5990), .ZN(n5896) );
  INV_X1 U3731 ( .A(n5964), .ZN(n5225) );
  INV_X1 U3732 ( .A(n5508), .ZN(n5182) );
  AOI22_X1 U3733 ( .A1(n3225), .A2(n5508), .B1(n6029), .B2(n5864), .ZN(n5520)
         );
  NAND3_X2 U3734 ( .A1(n4215), .A2(n4214), .A3(n4442), .ZN(n4216) );
  NAND3_X2 U3735 ( .A1(\wb/dsize_reg/z2 [4]), .A2(n4355), .A3(n3176), .ZN(
        n4214) );
  NOR3_X2 U3736 ( .A1(n4190), .A2(n4189), .A3(n4188), .ZN(n4197) );
  NOR2_X2 U3737 ( .A1(n4194), .A2(n4189), .ZN(n4007) );
  NOR2_X1 U3738 ( .A1(n5197), .A2(n5196), .ZN(n5202) );
  INV_X1 U3739 ( .A(n5196), .ZN(n4742) );
  AOI211_X2 U3740 ( .C1(n4773), .C2(n4762), .A(n4761), .B(n4760), .ZN(n4789)
         );
  OAI21_X1 U3741 ( .B1(n4773), .B2(n3230), .A(n3227), .ZN(n4758) );
  AOI21_X2 U3742 ( .B1(n5794), .B2(n5820), .A(n5793), .ZN(n5795) );
  OAI222_X1 U3743 ( .A1(n6308), .A2(n4162), .B1(n2666), .B2(n3152), .C1(n3154), 
        .C2(n2977), .ZN(regWrData[27]) );
  OAI222_X1 U3744 ( .A1(n6309), .A2(n4162), .B1(n2686), .B2(n3152), .C1(n3154), 
        .C2(n3023), .ZN(regWrData[28]) );
  OAI222_X1 U3745 ( .A1(n6334), .A2(n4162), .B1(n2703), .B2(n3152), .C1(n3154), 
        .C2(n2985), .ZN(regWrData[25]) );
  OAI222_X1 U3746 ( .A1(n6336), .A2(n4162), .B1(n2707), .B2(n3152), .C1(n3154), 
        .C2(n2978), .ZN(regWrData[23]) );
  OAI222_X1 U3747 ( .A1(n6324), .A2(n4162), .B1(n2673), .B2(n3152), .C1(n3154), 
        .C2(n2986), .ZN(regWrData[29]) );
  OAI222_X1 U3748 ( .A1(n6335), .A2(n4162), .B1(n2667), .B2(n3152), .C1(n3154), 
        .C2(n2979), .ZN(regWrData[24]) );
  OAI222_X1 U3749 ( .A1(n6338), .A2(n4162), .B1(n2719), .B2(n3152), .C1(n3154), 
        .C2(n2987), .ZN(regWrData[21]) );
  OAI22_X2 U3750 ( .A1(n3154), .A2(n2982), .B1(n6305), .B2(n4162), .ZN(n4474)
         );
  AOI21_X2 U3751 ( .B1(n4929), .B2(n4837), .A(n3218), .ZN(n4778) );
  INV_X4 U3752 ( .A(n5543), .ZN(n3060) );
  INV_X4 U3753 ( .A(n5720), .ZN(n3063) );
  AOI21_X2 U3754 ( .B1(n5818), .B2(n5817), .A(n2714), .ZN(n5819) );
  AOI21_X2 U3755 ( .B1(n5792), .B2(n5817), .A(n5791), .ZN(n5793) );
  OAI21_X1 U3756 ( .B1(n2668), .B2(n4442), .A(n4441), .ZN(n4443) );
  OAI21_X1 U3757 ( .B1(n2670), .B2(n4442), .A(n4183), .ZN(n4002) );
  NOR2_X2 U3758 ( .A1(n2699), .A2(n4442), .ZN(n3979) );
  NAND3_X4 U3759 ( .A1(n4569), .A2(n4568), .A3(n4801), .ZN(n4673) );
  INV_X4 U3760 ( .A(n6310), .ZN(n3064) );
  INV_X1 U3761 ( .A(n5885), .ZN(n5217) );
  NAND2_X2 U3762 ( .A1(n5885), .A2(n5013), .ZN(n5014) );
  NAND2_X4 U3763 ( .A1(n5222), .A2(n5221), .ZN(n5224) );
  OAI211_X2 U3764 ( .C1(n5917), .C2(n5916), .A(n3069), .B(n5220), .ZN(n5222)
         );
  INV_X4 U3765 ( .A(n6237), .ZN(n3066) );
  INV_X8 U3766 ( .A(n3066), .ZN(n3067) );
  AOI21_X4 U3767 ( .B1(n3930), .B2(n3178), .A(n3929), .ZN(n3931) );
  OAI22_X2 U3768 ( .A1(n6299), .A2(n3148), .B1(n6564), .B2(n3150), .ZN(n3929)
         );
  INV_X8 U3769 ( .A(n3068), .ZN(n3069) );
  AND3_X4 U3770 ( .A1(n4098), .A2(memAddr[11]), .A3(n3159), .ZN(n3070) );
  INV_X8 U3771 ( .A(n3070), .ZN(n4359) );
  XNOR2_X2 U3772 ( .A(n5071), .B(n3221), .ZN(n3071) );
  INV_X4 U3773 ( .A(n3071), .ZN(n5100) );
  NOR2_X2 U3774 ( .A1(n6618), .A2(n6617), .ZN(n4545) );
  NAND3_X2 U3775 ( .A1(n6618), .A2(n6603), .A3(n6600), .ZN(n4523) );
  NAND4_X2 U3776 ( .A1(n3055), .A2(n3064), .A3(n3235), .A4(n4029), .ZN(n4152)
         );
  XNOR2_X1 U3777 ( .A(n6279), .B(n3712), .ZN(n3713) );
  AOI22_X2 U3778 ( .A1(n5932), .A2(n6029), .B1(n5546), .B2(n5948), .ZN(n4873)
         );
  INV_X4 U3779 ( .A(n3077), .ZN(n4876) );
  OAI211_X1 U3780 ( .C1(n4846), .C2(n3078), .A(n3079), .B(n3080), .ZN(n3077)
         );
  INV_X2 U3781 ( .A(n4999), .ZN(n5798) );
  INV_X8 U3782 ( .A(n4357), .ZN(n3091) );
  XNOR2_X1 U3783 ( .A(n6264), .B(n3076), .ZN(n3728) );
  INV_X4 U3784 ( .A(n3324), .ZN(n3727) );
  NAND3_X2 U3785 ( .A1(n5415), .A2(n5416), .A3(n3033), .ZN(\ex_mem/N208 ) );
  NAND2_X1 U3786 ( .A1(n4989), .A2(n5544), .ZN(n5417) );
  NOR2_X2 U3787 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  XNOR2_X1 U3788 ( .A(n6183), .B(n3685), .ZN(n3686) );
  AOI22_X1 U3789 ( .A1(n5695), .A2(n4855), .B1(n5514), .B2(n4782), .ZN(n4783)
         );
  INV_X2 U3790 ( .A(n4782), .ZN(n4753) );
  AOI22_X1 U3791 ( .A1(n5695), .A2(n4858), .B1(n5505), .B2(n4782), .ZN(n4521)
         );
  OAI21_X2 U3792 ( .B1(n5481), .B2(n2627), .A(n5131), .ZN(n5132) );
  OAI21_X2 U3793 ( .B1(n5120), .B2(n2626), .A(n5119), .ZN(n5133) );
  NOR2_X1 U3794 ( .A1(n5798), .A2(n2627), .ZN(n5801) );
  NOR2_X1 U3795 ( .A1(n5798), .A2(n2779), .ZN(n5563) );
  NOR2_X2 U3796 ( .A1(n5801), .A2(n5800), .ZN(n5804) );
  NOR2_X2 U3797 ( .A1(n5563), .A2(n5562), .ZN(n5566) );
  NAND2_X2 U3798 ( .A1(n3814), .A2(n3813), .ZN(n3815) );
  NAND2_X1 U3799 ( .A1(n2711), .A2(n3586), .ZN(n3344) );
  NAND2_X1 U3800 ( .A1(n3586), .A2(n3606), .ZN(n3621) );
  NAND2_X4 U3801 ( .A1(n3586), .A2(n3633), .ZN(n3409) );
  AOI22_X1 U3802 ( .A1(n5695), .A2(n5438), .B1(n5505), .B2(n5087), .ZN(n5088)
         );
  NAND3_X2 U3803 ( .A1(n4984), .A2(n4983), .A3(n4982), .ZN(n5438) );
  NOR3_X2 U3804 ( .A1(n3344), .A2(n3478), .A3(n3343), .ZN(n3376) );
  NAND2_X1 U3805 ( .A1(n5504), .A2(n5695), .ZN(n5434) );
  AOI21_X1 U3806 ( .B1(n4867), .B2(n5504), .A(n2905), .ZN(n4964) );
  AOI22_X1 U3807 ( .A1(n5514), .A2(n5504), .B1(n5503), .B2(n5695), .ZN(n4861)
         );
  OAI21_X2 U3808 ( .B1(n4961), .B2(n4859), .A(n6018), .ZN(n5504) );
  NAND2_X4 U3809 ( .A1(n3546), .A2(n3457), .ZN(n3494) );
  NAND2_X4 U3810 ( .A1(n5435), .A2(n4985), .ZN(n4986) );
  XNOR2_X1 U3811 ( .A(n3766), .B(n3765), .ZN(n3920) );
  NOR2_X2 U3812 ( .A1(n5412), .A2(n2778), .ZN(n4761) );
  NOR2_X2 U3813 ( .A1(n5412), .A2(n2779), .ZN(n5227) );
  INV_X2 U3814 ( .A(n5412), .ZN(n5384) );
  NOR2_X1 U3815 ( .A1(n5412), .A2(n2627), .ZN(n5413) );
  AOI22_X4 U3816 ( .A1(n5695), .A2(n4864), .B1(n5514), .B2(n4828), .ZN(n4741)
         );
  NAND2_X4 U3817 ( .A1(n4726), .A2(n4725), .ZN(n4828) );
  XNOR2_X1 U3818 ( .A(n6272), .B(n3696), .ZN(n3697) );
  AND2_X4 U3819 ( .A1(n4827), .A2(n3226), .ZN(n3078) );
  OR2_X2 U3820 ( .A1(n5209), .A2(n2779), .ZN(n3079) );
  OR2_X4 U3821 ( .A1(n4835), .A2(n4847), .ZN(n3080) );
  NAND2_X1 U3822 ( .A1(n5127), .A2(n4811), .ZN(n4813) );
  NOR2_X1 U3823 ( .A1(n5357), .A2(n2777), .ZN(n5358) );
  NOR2_X2 U3824 ( .A1(n5357), .A2(n2625), .ZN(n4869) );
  OAI21_X2 U3825 ( .B1(n2580), .B2(n3392), .A(n3391), .ZN(iAddr[31]) );
  NAND3_X1 U3826 ( .A1(n3142), .A2(n3807), .A3(n3806), .ZN(n3810) );
  NOR2_X1 U3827 ( .A1(n3665), .A2(n3807), .ZN(n3667) );
  XNOR2_X1 U3828 ( .A(n6270), .B(n3700), .ZN(n3701) );
  NAND2_X1 U3829 ( .A1(n3484), .A2(n3483), .ZN(n3486) );
  NAND3_X1 U3830 ( .A1(n3357), .A2(n3459), .A3(n3356), .ZN(n3358) );
  NAND2_X4 U3831 ( .A1(n3356), .A2(n3357), .ZN(n3461) );
  XNOR2_X1 U3832 ( .A(n3719), .B(n2683), .ZN(n3720) );
  XNOR2_X1 U3833 ( .A(n6268), .B(n3704), .ZN(n3705) );
  AOI22_X2 U3834 ( .A1(n3225), .A2(n5586), .B1(n6029), .B2(n5680), .ZN(n5588)
         );
  NOR3_X2 U3835 ( .A1(n4745), .A2(n4744), .A3(n4743), .ZN(n4746) );
  AOI22_X1 U3836 ( .A1(n6029), .A2(n5939), .B1(n5938), .B2(n5937), .ZN(n5957)
         );
  INV_X2 U3837 ( .A(n5937), .ZN(n4898) );
  INV_X1 U3838 ( .A(n3371), .ZN(n3372) );
  NOR2_X2 U3839 ( .A1(n6561), .A2(n3150), .ZN(n3936) );
  OAI22_X2 U3840 ( .A1(n6291), .A2(n3148), .B1(n6554), .B2(n3150), .ZN(n4277)
         );
  NAND2_X1 U3841 ( .A1(n5505), .A2(n5511), .ZN(n5517) );
  OAI211_X1 U3842 ( .C1(n6037), .C2(n6044), .A(n6042), .B(n6043), .ZN(n5716)
         );
  OAI211_X4 U3843 ( .C1(n3510), .C2(n3143), .A(n3509), .B(n3508), .ZN(
        iAddr[11]) );
  INV_X2 U3844 ( .A(n3494), .ZN(n3498) );
  OAI22_X4 U3845 ( .A1(n5000), .A2(n2778), .B1(n5798), .B2(n2626), .ZN(n5001)
         );
  NAND2_X4 U3846 ( .A1(n5298), .A2(n5505), .ZN(n5300) );
  NOR3_X2 U3847 ( .A1(n5280), .A2(n5279), .A3(n5278), .ZN(n5295) );
  NOR3_X2 U3848 ( .A1(n5661), .A2(n5275), .A3(n2589), .ZN(n5279) );
  INV_X1 U3849 ( .A(iAddr[10]), .ZN(n3763) );
  NAND2_X1 U3850 ( .A1(n5509), .A2(n5695), .ZN(n3081) );
  AND2_X4 U3851 ( .A1(n3081), .A2(n3082), .ZN(n5128) );
  NAND3_X4 U3852 ( .A1(n4933), .A2(n4984), .A3(n4932), .ZN(n5511) );
  NAND2_X2 U3853 ( .A1(n3451), .A2(n3538), .ZN(n3542) );
  NAND2_X4 U3854 ( .A1(n3345), .A2(n3752), .ZN(n3512) );
  AOI21_X4 U3855 ( .B1(n3592), .B2(n3593), .A(n3143), .ZN(n3591) );
  NAND2_X4 U3856 ( .A1(n3364), .A2(n3496), .ZN(n3371) );
  NAND3_X2 U3857 ( .A1(n3611), .A2(n3598), .A3(n3597), .ZN(n3334) );
  NAND3_X2 U3858 ( .A1(n4802), .A2(n5837), .A3(n5038), .ZN(n4769) );
  NAND2_X2 U3859 ( .A1(n5039), .A2(n5038), .ZN(n5750) );
  AOI22_X4 U3860 ( .A1(n4129), .A2(n2606), .B1(n4524), .B2(memAddr[18]), .ZN(
        n4109) );
  INV_X4 U3861 ( .A(n4474), .ZN(n4080) );
  INV_X2 U3862 ( .A(n4232), .ZN(n4090) );
  NAND3_X2 U3863 ( .A1(n4231), .A2(n4233), .A3(n4232), .ZN(n4234) );
  AOI21_X1 U3864 ( .B1(n3994), .B2(n3993), .A(n3211), .ZN(\ex_mem/N108 ) );
  INV_X8 U3865 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U3866 ( .A1(n5080), .A2(n5631), .ZN(n4703) );
  NAND2_X1 U3867 ( .A1(n4974), .A2(n5080), .ZN(n5265) );
  NAND2_X1 U3868 ( .A1(n5080), .A2(n5662), .ZN(n4509) );
  NAND2_X1 U3869 ( .A1(n5080), .A2(n4818), .ZN(n4732) );
  NAND2_X1 U3870 ( .A1(n5080), .A2(n4911), .ZN(n4709) );
  NAND2_X1 U3871 ( .A1(n5080), .A2(n5707), .ZN(n4467) );
  INV_X16 U3872 ( .A(n4357), .ZN(n3087) );
  NOR4_X1 U3873 ( .A1(n5322), .A2(n5930), .A3(n5190), .A4(n5189), .ZN(n5191)
         );
  INV_X1 U3874 ( .A(n5189), .ZN(n4910) );
  XNOR2_X1 U3875 ( .A(n4880), .B(n3222), .ZN(n4554) );
  AOI21_X1 U3876 ( .B1(n3171), .B2(regWrData[8]), .A(n4290), .ZN(n4034) );
  INV_X4 U3877 ( .A(regWrData[8]), .ZN(n4466) );
  NAND3_X2 U3878 ( .A1(n4033), .A2(n4032), .A3(n4031), .ZN(regWrData[8]) );
  INV_X2 U3879 ( .A(n3085), .ZN(n4319) );
  INV_X2 U3880 ( .A(n4163), .ZN(n3999) );
  NAND3_X1 U3881 ( .A1(n5525), .A2(n5639), .A3(n5533), .ZN(n5420) );
  NAND2_X1 U3882 ( .A1(n4129), .A2(n2657), .ZN(n4220) );
  NAND2_X2 U3883 ( .A1(n4129), .A2(n2638), .ZN(n4284) );
  INV_X2 U3884 ( .A(n4604), .ZN(n4606) );
  INV_X1 U3885 ( .A(n5526), .ZN(n5527) );
  NAND3_X4 U3886 ( .A1(n3171), .A2(\wb/dsize_reg/z2 [28]), .A3(n3151), .ZN(
        n4140) );
  NOR2_X2 U3887 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  INV_X2 U3888 ( .A(n5586), .ZN(n5137) );
  NOR2_X1 U3889 ( .A1(n5174), .A2(n5586), .ZN(n5175) );
  NOR2_X1 U3890 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  INV_X2 U3891 ( .A(n3123), .ZN(n4193) );
  NAND3_X1 U3892 ( .A1(n4153), .A2(\wb/dsize_reg/z2 [25]), .A3(n3167), .ZN(
        n4158) );
  NAND2_X2 U3893 ( .A1(n2680), .A2(regWrData[13]), .ZN(n3088) );
  NAND2_X2 U3894 ( .A1(n5490), .A2(n5494), .ZN(n3099) );
  NAND2_X1 U3895 ( .A1(n5467), .A2(n5466), .ZN(n3089) );
  NAND3_X2 U3896 ( .A1(n4509), .A2(n3216), .A3(n4508), .ZN(n5122) );
  OAI21_X2 U3897 ( .B1(n5290), .B2(n5616), .A(n5306), .ZN(n5291) );
  NAND3_X1 U3898 ( .A1(n4724), .A2(n3217), .A3(n4723), .ZN(n5079) );
  NAND3_X1 U3899 ( .A1(n4944), .A2(n3217), .A3(n4946), .ZN(n4683) );
  NAND3_X2 U3900 ( .A1(n4497), .A2(n3217), .A3(n4496), .ZN(n4959) );
  NAND3_X2 U3901 ( .A1(n4501), .A2(n3217), .A3(n4500), .ZN(n4939) );
  NAND2_X1 U3902 ( .A1(n5123), .A2(n3157), .ZN(n4854) );
  NAND2_X1 U3903 ( .A1(n4938), .A2(n3157), .ZN(n4781) );
  NAND2_X1 U3904 ( .A1(n4981), .A2(n5305), .ZN(n4932) );
  AOI21_X1 U3905 ( .B1(n5082), .B2(n5305), .A(n2836), .ZN(n4488) );
  AOI21_X1 U3906 ( .B1(n4981), .B2(n5706), .A(n2836), .ZN(n4734) );
  AOI221_X2 U3907 ( .B1(n5708), .B2(n5707), .C1(n2685), .C2(n5706), .A(n2853), 
        .ZN(n5714) );
  INV_X1 U3908 ( .A(n5122), .ZN(n4859) );
  NAND2_X1 U3909 ( .A1(n2605), .A2(n5122), .ZN(n4852) );
  AOI21_X2 U3910 ( .B1(n4981), .B2(n5122), .A(n2836), .ZN(n4520) );
  NAND2_X1 U3911 ( .A1(n4981), .A2(n5121), .ZN(n4853) );
  NAND2_X1 U3912 ( .A1(n5082), .A2(n5121), .ZN(n4519) );
  NAND2_X1 U3913 ( .A1(n2605), .A2(n6017), .ZN(n4687) );
  AOI21_X1 U3914 ( .B1(n4981), .B2(n6017), .A(n2836), .ZN(n4470) );
  OAI21_X2 U3915 ( .B1(n4965), .B2(n4960), .A(n6022), .ZN(n4924) );
  OAI21_X2 U3916 ( .B1(n4980), .B2(n4979), .A(n3157), .ZN(n4983) );
  INV_X2 U3917 ( .A(n5282), .ZN(n4967) );
  NAND2_X1 U3918 ( .A1(n5082), .A2(n5712), .ZN(n4733) );
  NAND3_X1 U3919 ( .A1(n5281), .A2(n2589), .A3(n2605), .ZN(n5287) );
  NOR2_X2 U3920 ( .A1(n5084), .A2(n5083), .ZN(n5085) );
  AOI21_X2 U3921 ( .B1(n4947), .B2(n3156), .A(n5711), .ZN(n4954) );
  NOR3_X2 U3922 ( .A1(n4937), .A2(n5711), .A3(n4936), .ZN(n4942) );
  NOR2_X1 U3923 ( .A1(n3156), .A2(n5711), .ZN(n5690) );
  NOR3_X1 U3924 ( .A1(n5270), .A2(n5711), .A3(n5269), .ZN(n4977) );
  OAI221_X2 U3925 ( .B1(n5313), .B2(n5312), .C1(n5311), .C2(n5310), .A(n5127), 
        .ZN(n6028) );
  NAND2_X1 U3926 ( .A1(n4981), .A2(n5079), .ZN(n4865) );
  NAND2_X1 U3927 ( .A1(n5082), .A2(n5079), .ZN(n4725) );
  INV_X2 U3928 ( .A(n5274), .ZN(n5275) );
  OAI21_X2 U3929 ( .B1(n4960), .B2(n4959), .A(n6022), .ZN(n5499) );
  NAND2_X1 U3930 ( .A1(n2605), .A2(n4959), .ZN(n4779) );
  AOI21_X1 U3931 ( .B1(n4981), .B2(n4959), .A(n2836), .ZN(n4503) );
  AOI22_X2 U3932 ( .A1(n4939), .A2(n2605), .B1(n4959), .B2(n2685), .ZN(n4940)
         );
  NAND4_X2 U3933 ( .A1(n5889), .A2(n5921), .A3(n2720), .A4(n5915), .ZN(n5893)
         );
  XOR2_X2 U3934 ( .A(n3223), .B(n4838), .Z(n3090) );
  INV_X16 U3935 ( .A(n3219), .ZN(n3223) );
  NAND2_X2 U3936 ( .A1(n4524), .A2(memAddr[5]), .ZN(n4404) );
  INV_X8 U3937 ( .A(n4394), .ZN(n4114) );
  NAND2_X1 U3938 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  NAND3_X2 U3939 ( .A1(n4714), .A2(n3216), .A3(n4713), .ZN(n5281) );
  NAND3_X2 U3940 ( .A1(n4430), .A2(n5346), .A3(n3063), .ZN(n4449) );
  NAND3_X2 U3941 ( .A1(n4059), .A2(n4058), .A3(n4057), .ZN(n4246) );
  NAND2_X1 U3942 ( .A1(n5080), .A2(n5369), .ZN(n4713) );
  XNOR2_X2 U3943 ( .A(n2724), .B(n4837), .ZN(n5011) );
  NAND2_X4 U3944 ( .A1(n3363), .A2(n3464), .ZN(n3496) );
  OAI21_X1 U3945 ( .B1(iAddr[12]), .B2(n3734), .A(n3767), .ZN(n3824) );
  INV_X8 U3946 ( .A(n3672), .ZN(n3734) );
  NAND2_X1 U3947 ( .A1(n3231), .A2(n2577), .ZN(n4917) );
  INV_X1 U3948 ( .A(n2577), .ZN(n4921) );
  NAND3_X2 U3949 ( .A1(n5071), .A2(n2577), .A3(n4453), .ZN(n4429) );
  NAND3_X1 U3950 ( .A1(n5554), .A2(n4763), .A3(n2577), .ZN(n4416) );
  INV_X1 U3951 ( .A(n3411), .ZN(n3412) );
  NOR2_X2 U3952 ( .A1(n5764), .A2(n5765), .ZN(n5761) );
  INV_X1 U3953 ( .A(n5725), .ZN(n5239) );
  NAND2_X1 U3954 ( .A1(n5731), .A2(n5725), .ZN(n5242) );
  INV_X2 U3955 ( .A(iAddr[2]), .ZN(n3829) );
  INV_X1 U3956 ( .A(n3747), .ZN(n3748) );
  NAND2_X1 U3957 ( .A1(iAddr[3]), .A2(iAddr[2]), .ZN(n3749) );
  INV_X4 U3958 ( .A(n3747), .ZN(n3670) );
  NOR2_X2 U3959 ( .A1(n4429), .A2(n4428), .ZN(n4436) );
  NOR2_X2 U3960 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  INV_X1 U3961 ( .A(n5889), .ZN(n5025) );
  NOR2_X2 U3962 ( .A1(n5764), .A2(n5769), .ZN(n5759) );
  NAND3_X2 U3963 ( .A1(n5743), .A2(n5742), .A3(n5741), .ZN(n5744) );
  OAI21_X1 U3964 ( .B1(n5699), .B2(n6091), .A(n6016), .ZN(n5717) );
  OAI22_X1 U3965 ( .A1(n5773), .A2(n2592), .B1(n6016), .B2(n2778), .ZN(n5775)
         );
  AOI21_X1 U3966 ( .B1(n6036), .B2(n6016), .A(n2627), .ZN(n6021) );
  NAND3_X2 U3967 ( .A1(n4971), .A2(n4984), .A3(n4970), .ZN(n5436) );
  NOR2_X1 U3968 ( .A1(n5699), .A2(n5698), .ZN(n5703) );
  NAND2_X2 U3969 ( .A1(n5307), .A2(n5306), .ZN(n5312) );
  NAND3_X1 U3970 ( .A1(n5309), .A2(n5308), .A3(n5307), .ZN(n5311) );
  NAND2_X2 U3971 ( .A1(n4362), .A2(n4361), .ZN(n4363) );
  AOI21_X4 U3972 ( .B1(n3361), .B2(n3464), .A(n3360), .ZN(n3364) );
  NAND2_X1 U3973 ( .A1(n4298), .A2(n4297), .ZN(n3092) );
  AOI211_X1 U3974 ( .C1(n2605), .C2(n5712), .A(n5711), .B(n5710), .ZN(n5713)
         );
  NOR2_X1 U3975 ( .A1(n5705), .A2(n3157), .ZN(n5708) );
  NAND2_X2 U3976 ( .A1(n4524), .A2(memAddr[13]), .ZN(n3093) );
  NOR3_X4 U3977 ( .A1(n5664), .A2(n4667), .A3(n4655), .ZN(n4660) );
  OAI21_X2 U3978 ( .B1(n4245), .B2(n4244), .A(n4243), .ZN(n3094) );
  MUX2_X2 U3979 ( .A(n3949), .B(n6622), .S(n3097), .Z(n3096) );
  INV_X4 U3980 ( .A(n3096), .ZN(n5884) );
  NAND3_X2 U3981 ( .A1(n3948), .A2(n3947), .A3(n3946), .ZN(n4230) );
  INV_X8 U3982 ( .A(n3244), .ZN(n3243) );
  NOR2_X1 U3983 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NOR3_X1 U3984 ( .A1(n5529), .A2(n5528), .A3(n5527), .ZN(n5534) );
  INV_X2 U3985 ( .A(n5494), .ZN(n5489) );
  INV_X4 U3986 ( .A(n5494), .ZN(n3098) );
  NAND3_X2 U3987 ( .A1(n5834), .A2(n5921), .A3(n5833), .ZN(n5835) );
  NAND3_X2 U3988 ( .A1(n4248), .A2(n4247), .A3(n4249), .ZN(n3101) );
  INV_X4 U3989 ( .A(n3101), .ZN(n3102) );
  INV_X2 U3990 ( .A(n4250), .ZN(n3925) );
  NAND3_X2 U3991 ( .A1(\wb/dsize_reg/z2 [7]), .A2(n3167), .A3(n4355), .ZN(
        n4247) );
  NAND3_X1 U3992 ( .A1(n4357), .A2(n3167), .A3(n3031), .ZN(n4248) );
  INV_X4 U3993 ( .A(n3103), .ZN(n4331) );
  AOI211_X1 U3994 ( .C1(n5790), .C2(n5789), .A(n5788), .B(n5787), .ZN(n5806)
         );
  OAI21_X1 U3995 ( .B1(n5790), .B2(n3229), .A(n6008), .ZN(n5784) );
  INV_X8 U3996 ( .A(n5790), .ZN(n5005) );
  NAND3_X2 U3997 ( .A1(n3972), .A2(n3971), .A3(n3970), .ZN(n4373) );
  NAND2_X2 U3998 ( .A1(n5670), .A2(n5274), .ZN(n4738) );
  AOI22_X2 U3999 ( .A1(n4129), .A2(n2607), .B1(n4524), .B2(memAddr[24]), .ZN(
        n3961) );
  NOR2_X2 U4000 ( .A1(n5989), .A2(n5988), .ZN(n5992) );
  AOI21_X1 U4001 ( .B1(n5491), .B2(n3226), .A(n5490), .ZN(n5497) );
  NAND2_X1 U4002 ( .A1(n5644), .A2(n5420), .ZN(n5421) );
  NAND2_X1 U4003 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  INV_X2 U4004 ( .A(n5644), .ZN(n5640) );
  AOI21_X4 U4005 ( .B1(n4601), .B2(n5644), .A(n5343), .ZN(n4605) );
  NAND3_X2 U4006 ( .A1(n5490), .A2(n5346), .A3(n4430), .ZN(n4273) );
  INV_X8 U4007 ( .A(n3120), .ZN(n3146) );
  XNOR2_X2 U4008 ( .A(n4680), .B(n4679), .ZN(n4771) );
  OAI221_X4 U4009 ( .B1(n6585), .B2(n3155), .C1(n3185), .C2(n4146), .A(n4145), 
        .ZN(n5196) );
  INV_X1 U4010 ( .A(n5041), .ZN(n4766) );
  NAND3_X2 U4011 ( .A1(n5042), .A2(n5041), .A3(n5040), .ZN(n5841) );
  NAND2_X2 U4012 ( .A1(n2620), .A2(n4610), .ZN(n5041) );
  INV_X2 U4013 ( .A(n4229), .ZN(n4125) );
  OAI21_X1 U4014 ( .B1(n5740), .B2(n5106), .A(n5754), .ZN(n5107) );
  INV_X2 U4015 ( .A(n5740), .ZN(n5742) );
  INV_X2 U4016 ( .A(n4358), .ZN(n4354) );
  XNOR2_X1 U4017 ( .A(n6188), .B(n3745), .ZN(n3746) );
  INV_X4 U4018 ( .A(n3316), .ZN(n3696) );
  XNOR2_X1 U4019 ( .A(n6196), .B(n6188), .ZN(n3517) );
  NAND2_X1 U4020 ( .A1(n4596), .A2(n5397), .ZN(n3106) );
  XNOR2_X1 U4021 ( .A(n5375), .B(n5374), .ZN(n5988) );
  NAND2_X4 U4022 ( .A1(n3633), .A2(n3600), .ZN(n3618) );
  NAND2_X4 U4023 ( .A1(n3407), .A2(n3600), .ZN(n3408) );
  NAND3_X4 U4024 ( .A1(n3370), .A2(n3107), .A3(n3369), .ZN(n3600) );
  NAND4_X2 U4025 ( .A1(n4331), .A2(n3178), .A3(\wb/dsize_reg/z2 [14]), .A4(
        n4355), .ZN(n4335) );
  INV_X4 U4026 ( .A(n5888), .ZN(n5915) );
  NOR2_X1 U4027 ( .A1(n4473), .A2(n4472), .ZN(n4475) );
  NOR2_X1 U4028 ( .A1(n4471), .A2(n4473), .ZN(n4081) );
  OAI211_X4 U4029 ( .C1(n5086), .C2(n3157), .A(n5692), .B(n5085), .ZN(n5298)
         );
  NAND2_X2 U4030 ( .A1(n3483), .A2(n3367), .ZN(n3107) );
  NAND2_X1 U4031 ( .A1(n2577), .A2(n3094), .ZN(n4451) );
  NAND2_X1 U4032 ( .A1(n4763), .A2(n3094), .ZN(n4426) );
  INV_X1 U4033 ( .A(n3094), .ZN(n4816) );
  AOI21_X1 U4034 ( .B1(n4084), .B2(n4329), .A(n3211), .ZN(\ex_mem/N113 ) );
  INV_X2 U4035 ( .A(n4888), .ZN(n4800) );
  XOR2_X1 U4036 ( .A(n3223), .B(n3061), .Z(n3109) );
  INV_X4 U4037 ( .A(n5423), .ZN(n5707) );
  INV_X4 U4038 ( .A(n5750), .ZN(n5046) );
  INV_X1 U4039 ( .A(n5046), .ZN(n3127) );
  INV_X4 U4040 ( .A(n3217), .ZN(n3110) );
  INV_X1 U4041 ( .A(n5392), .ZN(n5402) );
  NAND3_X1 U4042 ( .A1(n3096), .A2(n4838), .A3(n5392), .ZN(n4455) );
  OAI21_X2 U4043 ( .B1(n5402), .B2(n3230), .A(n3227), .ZN(n5403) );
  AOI211_X2 U4044 ( .C1(n5402), .C2(n5408), .A(n5407), .B(n5406), .ZN(n5418)
         );
  AND2_X4 U4045 ( .A1(n3125), .A2(n3120), .ZN(n4075) );
  INV_X8 U4046 ( .A(n5306), .ZN(n5711) );
  NAND3_X2 U4047 ( .A1(n5928), .A2(n5846), .A3(n5925), .ZN(n5027) );
  NAND2_X4 U4048 ( .A1(n3564), .A2(n3459), .ZN(n3568) );
  NAND2_X4 U4049 ( .A1(n3494), .A2(n3458), .ZN(n3564) );
  NAND3_X2 U4050 ( .A1(n3243), .A2(n4350), .A3(n4349), .ZN(n4352) );
  NAND2_X2 U4051 ( .A1(n4129), .A2(n2637), .ZN(n4340) );
  AND2_X2 U4052 ( .A1(n4524), .A2(memAddr[5]), .ZN(n3113) );
  NAND2_X2 U4053 ( .A1(n5839), .A2(n5846), .ZN(n5849) );
  NAND4_X2 U4054 ( .A1(n5034), .A2(n3059), .A3(n5400), .A4(n2587), .ZN(n5035)
         );
  INV_X1 U4055 ( .A(n3175), .ZN(n3181) );
  INV_X4 U4056 ( .A(n3175), .ZN(n3180) );
  NAND4_X1 U4057 ( .A1(n3488), .A2(n3107), .A3(n3486), .A4(n3485), .ZN(n3489)
         );
  OAI21_X1 U4058 ( .B1(n3475), .B2(n3474), .A(n3473), .ZN(n3490) );
  NAND4_X1 U4059 ( .A1(n6024), .A2(n6028), .A3(n6023), .A4(n6027), .ZN(n5771)
         );
  OAI21_X1 U4060 ( .B1(n5068), .B2(n3230), .A(n3227), .ZN(n5069) );
  NAND3_X1 U4061 ( .A1(n4732), .A2(n3216), .A3(n4731), .ZN(n5712) );
  NOR2_X1 U4062 ( .A1(n5377), .A2(n5068), .ZN(n4454) );
  NOR3_X1 U4063 ( .A1(n3180), .A2(n3234), .A3(n3032), .ZN(n5145) );
  NOR3_X2 U4064 ( .A1(n3180), .A2(n3234), .A3(n3022), .ZN(n4191) );
  NOR2_X1 U4065 ( .A1(n3234), .A2(n2977), .ZN(n4128) );
  NOR2_X1 U4066 ( .A1(n3234), .A2(n2978), .ZN(n3952) );
  NOR2_X1 U4067 ( .A1(n3234), .A2(n2979), .ZN(n3960) );
  NOR2_X1 U4068 ( .A1(n3234), .A2(n2874), .ZN(n4094) );
  NOR2_X1 U4069 ( .A1(n3234), .A2(n2922), .ZN(n4103) );
  NAND4_X1 U4070 ( .A1(n4170), .A2(n3178), .A3(\wb/dsize_reg/z2 [16]), .A4(
        n3234), .ZN(n4150) );
  NAND4_X1 U4071 ( .A1(n4170), .A2(n3234), .A3(\wb/dsize_reg/z2 [9]), .A4(
        n3167), .ZN(n4157) );
  NOR2_X2 U4072 ( .A1(n4077), .A2(n4076), .ZN(n4654) );
  INV_X1 U4073 ( .A(n4654), .ZN(regWrData[5]) );
  INV_X1 U4074 ( .A(n3139), .ZN(n3114) );
  AOI21_X2 U4075 ( .B1(n5037), .B2(n5036), .A(n5035), .ZN(n5039) );
  INV_X2 U4076 ( .A(n5625), .ZN(n5301) );
  AOI22_X1 U4077 ( .A1(n5947), .A2(n5771), .B1(n6029), .B2(n5625), .ZN(n5606)
         );
  AOI22_X1 U4078 ( .A1(n5363), .A2(n5626), .B1(n5947), .B2(n5625), .ZN(n5627)
         );
  OAI21_X1 U4079 ( .B1(n4960), .B2(n5274), .A(n6022), .ZN(n5257) );
  AOI21_X1 U4080 ( .B1(n4981), .B2(n5274), .A(n2836), .ZN(n4706) );
  NOR3_X1 U4081 ( .A1(n3180), .A2(n6329), .A3(n3146), .ZN(n4614) );
  NOR2_X1 U4082 ( .A1(n6301), .A2(n3091), .ZN(n4092) );
  XNOR2_X1 U4083 ( .A(n3687), .B(n2684), .ZN(n3688) );
  INV_X4 U4084 ( .A(n3322), .ZN(n3708) );
  OAI211_X4 U4085 ( .C1(n4807), .C2(n5373), .A(n4806), .B(n4805), .ZN(n4808)
         );
  NOR3_X2 U4086 ( .A1(n3180), .A2(n6328), .A3(n3146), .ZN(n4189) );
  XOR2_X2 U4087 ( .A(n3223), .B(n4846), .Z(n3116) );
  OAI21_X1 U4088 ( .B1(n3575), .B2(n3438), .A(n3437), .ZN(n3439) );
  INV_X1 U4089 ( .A(n3397), .ZN(n3395) );
  NOR2_X1 U4090 ( .A1(n3612), .A2(n3409), .ZN(n3410) );
  AOI21_X1 U4091 ( .B1(n4000), .B2(n4164), .A(n3211), .ZN(\ex_mem/N101 ) );
  OAI21_X1 U4092 ( .B1(n5273), .B2(n2589), .A(n5272), .ZN(n5280) );
  NAND3_X1 U4093 ( .A1(n5282), .A2(n2589), .A3(n3156), .ZN(n5286) );
  NAND2_X1 U4094 ( .A1(n6040), .A2(n5610), .ZN(n5510) );
  NOR2_X1 U4095 ( .A1(n6182), .A2(n3148), .ZN(n4138) );
  NOR2_X1 U4096 ( .A1(n6284), .A2(n3148), .ZN(n4018) );
  NOR2_X1 U4097 ( .A1(n6294), .A2(n3148), .ZN(n3967) );
  NOR2_X1 U4098 ( .A1(n6258), .A2(n3148), .ZN(n4062) );
  NOR2_X1 U4099 ( .A1(n6298), .A2(n3148), .ZN(n3935) );
  NOR2_X1 U4100 ( .A1(n6175), .A2(n3148), .ZN(n4111) );
  NOR2_X1 U4101 ( .A1(n6297), .A2(n3148), .ZN(n3942) );
  OAI221_X2 U4102 ( .B1(n4635), .B2(n4636), .C1(n3243), .C2(n4634), .A(n4633), 
        .ZN(n4641) );
  NAND2_X4 U4103 ( .A1(n4661), .A2(n5531), .ZN(n3117) );
  NAND3_X2 U4104 ( .A1(iAddr[17]), .A2(iAddr[16]), .A3(n3772), .ZN(n3775) );
  XNOR2_X1 U4105 ( .A(iAddr[17]), .B(n3782), .ZN(n3915) );
  NOR2_X4 U4106 ( .A1(n3118), .A2(n3119), .ZN(n3120) );
  OAI21_X1 U4107 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n5118) );
  NAND3_X2 U4108 ( .A1(n5114), .A2(n4763), .A3(n4995), .ZN(n4452) );
  NAND3_X2 U4109 ( .A1(n5114), .A2(n4995), .A3(n3096), .ZN(n4427) );
  INV_X32 U4110 ( .A(n3148), .ZN(n4524) );
  NAND2_X4 U4111 ( .A1(n4425), .A2(n5554), .ZN(n4450) );
  INV_X8 U4112 ( .A(n4424), .ZN(n4425) );
  NAND3_X4 U4113 ( .A1(n4957), .A2(n2900), .A3(n4958), .ZN(n5678) );
  AOI22_X2 U4114 ( .A1(n5127), .A2(n5314), .B1(n5505), .B2(n5509), .ZN(n4957)
         );
  NAND4_X4 U4115 ( .A1(n5633), .A2(n3092), .A3(n6091), .A4(n4675), .ZN(n4424)
         );
  INV_X4 U4116 ( .A(n5666), .ZN(n4668) );
  OAI21_X2 U4117 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5478) );
  OAI221_X4 U4118 ( .B1(n2680), .B2(n4495), .C1(n4494), .C2(n4493), .A(n3041), 
        .ZN(n5618) );
  NAND2_X4 U4119 ( .A1(n3995), .A2(n3167), .ZN(n4628) );
  INV_X2 U4120 ( .A(iAddr[4]), .ZN(n3750) );
  OAI21_X1 U4121 ( .B1(n3738), .B2(n3743), .A(n3737), .ZN(n3740) );
  OAI21_X1 U4122 ( .B1(n3742), .B2(n3747), .A(n3741), .ZN(n3744) );
  XNOR2_X1 U4123 ( .A(n3743), .B(iAddr[7]), .ZN(n3827) );
  XNOR2_X1 U4124 ( .A(n3747), .B(iAddr[5]), .ZN(n3823) );
  NAND3_X2 U4125 ( .A1(iAddr[4]), .A2(iAddr[3]), .A3(iAddr[2]), .ZN(n3747) );
  NAND2_X1 U4126 ( .A1(n5127), .A2(n5509), .ZN(n5518) );
  NAND4_X1 U4127 ( .A1(n4576), .A2(n4578), .A3(n4579), .A4(n4577), .ZN(
        regWrData[11]) );
  NAND4_X1 U4128 ( .A1(n5155), .A2(n4577), .A3(n5154), .A4(n4576), .ZN(n4582)
         );
  NAND4_X1 U4129 ( .A1(n3783), .A2(iAddr[21]), .A3(n3784), .A4(iAddr[17]), 
        .ZN(n3786) );
  NAND4_X1 U4130 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  INV_X2 U4131 ( .A(n3472), .ZN(n3473) );
  NAND3_X1 U4132 ( .A1(n3602), .A2(n3601), .A3(n3600), .ZN(n3394) );
  NAND2_X2 U4133 ( .A1(n3159), .A2(n3121), .ZN(n4403) );
  NAND2_X4 U4134 ( .A1(\wb/dsize_reg/z2 [8]), .A2(n4355), .ZN(n4027) );
  NAND2_X1 U4135 ( .A1(n5763), .A2(n5472), .ZN(n5474) );
  NAND3_X2 U4136 ( .A1(n4242), .A2(n3243), .A3(n4241), .ZN(n4244) );
  NAND3_X2 U4137 ( .A1(n4402), .A2(n4400), .A3(n4401), .ZN(n4076) );
  INV_X4 U4138 ( .A(\hazard_detect/eq_83/A[4] ), .ZN(n6411) );
  NAND2_X2 U4139 ( .A1(n6528), .A2(n6492), .ZN(\hazard_detect/eq_83/A[4] ) );
  NOR3_X2 U4140 ( .A1(n2780), .A2(n6420), .A3(n2662), .ZN(n6385) );
  NAND2_X2 U4141 ( .A1(n6587), .A2(n2594), .ZN(n6420) );
  OAI221_X2 U4142 ( .B1(n6491), .B2(n2604), .C1(n6372), .C2(n2837), .A(n6774), 
        .ZN(n6490) );
  NOR4_X2 U4143 ( .A1(n6126), .A2(n6125), .A3(n6135), .A4(n6133), .ZN(n6491)
         );
  NAND2_X4 U4144 ( .A1(n2990), .A2(n5731), .ZN(n5734) );
  OAI22_X2 U4145 ( .A1(n6259), .A2(n3148), .B1(n6556), .B2(n3150), .ZN(n4055)
         );
  INV_X2 U4146 ( .A(n5333), .ZN(n5335) );
  NAND2_X4 U4147 ( .A1(n6103), .A2(n6101), .ZN(n6056) );
  XNOR2_X1 U4148 ( .A(n5593), .B(n5592), .ZN(n5970) );
  INV_X2 U4149 ( .A(n4646), .ZN(n4621) );
  XNOR2_X1 U4150 ( .A(n5553), .B(n5642), .ZN(n5976) );
  NAND2_X4 U4151 ( .A1(n4630), .A2(n3243), .ZN(n4166) );
  NAND2_X4 U4152 ( .A1(n4665), .A2(n5575), .ZN(n4666) );
  INV_X8 U4153 ( .A(n4639), .ZN(n4630) );
  INV_X8 U4154 ( .A(n4161), .ZN(n3151) );
  OAI21_X2 U4155 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n5472) );
  XNOR2_X1 U4156 ( .A(n3732), .B(n2822), .ZN(n3733) );
  NOR2_X1 U4157 ( .A1(n6177), .A2(n3724), .ZN(n3725) );
  INV_X4 U4158 ( .A(n3320), .ZN(n3704) );
  XNOR2_X1 U4159 ( .A(n6197), .B(n6177), .ZN(n3539) );
  INV_X2 U4160 ( .A(n5188), .ZN(n4750) );
  NOR4_X1 U4161 ( .A1(n5386), .A2(n5188), .A3(n5624), .A4(n5187), .ZN(n5192)
         );
  NAND2_X1 U4162 ( .A1(n5887), .A2(n5885), .ZN(n4839) );
  NAND3_X1 U4163 ( .A1(n5920), .A2(n5919), .A3(n5918), .ZN(n5923) );
  NAND4_X1 U4164 ( .A1(n5919), .A2(n5918), .A3(n5920), .A4(n5831), .ZN(n5834)
         );
  OAI221_X4 U4165 ( .B1(n5443), .B2(n2625), .C1(n2843), .C2(n2777), .A(n5442), 
        .ZN(n5864) );
  NOR2_X2 U4166 ( .A1(n2673), .A2(n4073), .ZN(n4074) );
  NAND2_X4 U4167 ( .A1(n4524), .A2(memAddr[10]), .ZN(n4262) );
  OAI21_X1 U4168 ( .B1(n3228), .B2(n5944), .A(n5949), .ZN(n5945) );
  OAI21_X1 U4169 ( .B1(n5949), .B2(n3229), .A(n6008), .ZN(n5950) );
  XNOR2_X1 U4170 ( .A(n3223), .B(n5949), .ZN(n4610) );
  INV_X4 U4171 ( .A(n6311), .ZN(n3236) );
  NAND3_X2 U4172 ( .A1(n5921), .A2(n2720), .A3(n5915), .ZN(n5926) );
  NAND3_X1 U4173 ( .A1(n5923), .A2(n5922), .A3(n5921), .ZN(n5924) );
  INV_X2 U4174 ( .A(n5840), .ZN(n5843) );
  NOR3_X2 U4175 ( .A1(n3180), .A2(n2666), .A3(n4073), .ZN(n4194) );
  XNOR2_X1 U4176 ( .A(n5368), .B(n3222), .ZN(n4556) );
  NAND2_X1 U4177 ( .A1(n4342), .A2(n4348), .ZN(n4346) );
  NAND2_X1 U4178 ( .A1(n4344), .A2(n4348), .ZN(n4345) );
  NAND3_X2 U4179 ( .A1(n4139), .A2(n2848), .A3(n4348), .ZN(n4349) );
  NOR2_X2 U4180 ( .A1(n5002), .A2(n5001), .ZN(n5050) );
  INV_X1 U4181 ( .A(n3134), .ZN(n3126) );
  NAND2_X2 U4182 ( .A1(n4478), .A2(n4477), .ZN(n3133) );
  NAND2_X4 U4183 ( .A1(n4361), .A2(n3105), .ZN(n4358) );
  INV_X16 U4184 ( .A(n3218), .ZN(n3217) );
  NAND3_X2 U4185 ( .A1(n4171), .A2(n4170), .A3(\wb/dsize_reg/z2 [1]), .ZN(
        n4172) );
  NAND2_X2 U4186 ( .A1(n5377), .A2(n4564), .ZN(n3131) );
  NAND2_X4 U4187 ( .A1(n3585), .A2(n3593), .ZN(n3336) );
  INV_X1 U4188 ( .A(n3585), .ZN(n3590) );
  NAND2_X4 U4189 ( .A1(n3599), .A2(n3332), .ZN(n3597) );
  AOI21_X1 U4190 ( .B1(n3787), .B2(n3771), .A(n3784), .ZN(n3916) );
  INV_X1 U4191 ( .A(iAddr[11]), .ZN(n3765) );
  NOR3_X1 U4192 ( .A1(n3788), .A2(n3793), .A3(n3787), .ZN(n3790) );
  INV_X2 U4193 ( .A(n3556), .ZN(n3484) );
  NAND3_X1 U4194 ( .A1(n3142), .A2(n3556), .A3(n3555), .ZN(n3558) );
  INV_X1 U4195 ( .A(n3538), .ZN(n3540) );
  NAND2_X4 U4196 ( .A1(n3556), .A2(n3456), .ZN(n3546) );
  XNOR2_X1 U4197 ( .A(n3698), .B(n2824), .ZN(n3699) );
  XNOR2_X1 U4198 ( .A(n3710), .B(n2681), .ZN(n3711) );
  XNOR2_X1 U4199 ( .A(n3729), .B(n2823), .ZN(n3730) );
  XNOR2_X1 U4200 ( .A(n6187), .B(n3725), .ZN(n3726) );
  XNOR2_X1 U4201 ( .A(n6198), .B(n6187), .ZN(n3449) );
  INV_X1 U4202 ( .A(n5575), .ZN(n5576) );
  NOR2_X1 U4203 ( .A1(n6558), .A2(n3150), .ZN(n4137) );
  NOR2_X1 U4204 ( .A1(n6557), .A2(n3150), .ZN(n4019) );
  NOR2_X1 U4205 ( .A1(n6559), .A2(n3150), .ZN(n3966) );
  NOR2_X1 U4206 ( .A1(n6563), .A2(n3150), .ZN(n4061) );
  NOR2_X1 U4207 ( .A1(n6560), .A2(n3150), .ZN(n3943) );
  NOR2_X1 U4208 ( .A1(n6562), .A2(n3150), .ZN(n4112) );
  NAND2_X1 U4209 ( .A1(n3156), .A2(n5661), .ZN(n4227) );
  INV_X8 U4210 ( .A(n5817), .ZN(n5747) );
  NOR2_X2 U4211 ( .A1(n4902), .A2(n4901), .ZN(n4903) );
  AOI22_X1 U4212 ( .A1(n3225), .A2(n5386), .B1(n6029), .B2(n5385), .ZN(n5389)
         );
  AOI22_X1 U4213 ( .A1(n3225), .A2(n5188), .B1(n5948), .B2(n5385), .ZN(n4787)
         );
  NOR2_X1 U4214 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  NAND2_X2 U4215 ( .A1(n3159), .A2(n3067), .ZN(n4136) );
  OAI21_X2 U4216 ( .B1(n5893), .B2(n5892), .A(n5891), .ZN(n5894) );
  NAND3_X2 U4217 ( .A1(n3170), .A2(n2996), .A3(n4139), .ZN(n4142) );
  NAND3_X2 U4218 ( .A1(n5308), .A2(n5309), .A3(n3157), .ZN(n5313) );
  XNOR2_X2 U4219 ( .A(n4808), .B(n3059), .ZN(n5960) );
  OAI21_X4 U4220 ( .B1(n5917), .B2(n5916), .A(n3069), .ZN(n5892) );
  INV_X4 U4221 ( .A(n4564), .ZN(n3130) );
  INV_X4 U4222 ( .A(n3133), .ZN(n3134) );
  OAI21_X1 U4223 ( .B1(n4960), .B2(n4922), .A(n6022), .ZN(n4923) );
  NAND3_X1 U4224 ( .A1(n6085), .A2(n6084), .A3(n2622), .ZN(n6099) );
  AOI21_X2 U4225 ( .B1(n6080), .B2(n6084), .A(n6079), .ZN(n6081) );
  INV_X2 U4226 ( .A(n6084), .ZN(n6086) );
  NAND2_X1 U4227 ( .A1(n6005), .A2(n6084), .ZN(n5779) );
  AOI211_X2 U4228 ( .C1(n6005), .C2(n6047), .A(n5259), .B(n5258), .ZN(n5320)
         );
  NAND2_X4 U4229 ( .A1(n4298), .A2(n4297), .ZN(n5422) );
  NAND2_X1 U4230 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  NAND2_X1 U4231 ( .A1(n5763), .A2(n5762), .ZN(n5760) );
  INV_X2 U4232 ( .A(n5762), .ZN(n5768) );
  NAND3_X2 U4233 ( .A1(n6067), .A2(n6066), .A3(n6065), .ZN(n6072) );
  INV_X2 U4234 ( .A(n6064), .ZN(n6066) );
  INV_X4 U4235 ( .A(n6063), .ZN(n6067) );
  OAI221_X2 U4236 ( .B1(n3087), .B2(n6320), .C1(n3145), .C2(n2959), .A(n4261), 
        .ZN(n4267) );
  NAND3_X1 U4237 ( .A1(n5756), .A2(n5755), .A3(n5754), .ZN(n5758) );
  NAND2_X4 U4238 ( .A1(n5781), .A2(n5006), .ZN(n5755) );
  NAND2_X1 U4239 ( .A1(n6005), .A2(n5958), .ZN(n5935) );
  NOR2_X2 U4240 ( .A1(n6332), .A2(n3087), .ZN(n3980) );
  NAND2_X1 U4241 ( .A1(n4322), .A2(n4321), .ZN(n4323) );
  NAND2_X4 U4242 ( .A1(n5337), .A2(n5336), .ZN(n5396) );
  INV_X1 U4243 ( .A(n4403), .ZN(n4078) );
  INV_X8 U4244 ( .A(n3787), .ZN(n3772) );
  NAND2_X4 U4245 ( .A1(n3659), .A2(n2902), .ZN(n3527) );
  OAI21_X1 U4246 ( .B1(n5960), .B2(n2718), .A(n4810), .ZN(n4822) );
  OAI21_X1 U4247 ( .B1(n5667), .B2(n5666), .A(n5665), .ZN(n5669) );
  AOI211_X1 U4248 ( .C1(n3171), .C2(regWrData[7]), .A(n4254), .B(n4253), .ZN(
        n3926) );
  AOI211_X1 U4249 ( .C1(n6005), .C2(n6064), .A(n5077), .B(n5076), .ZN(n5097)
         );
  OAI21_X1 U4250 ( .B1(n4679), .B2(n3230), .A(n6008), .ZN(n4547) );
  NAND2_X1 U4251 ( .A1(n5013), .A2(n5042), .ZN(n4767) );
  NAND2_X1 U4252 ( .A1(n5015), .A2(n5013), .ZN(n4840) );
  NAND2_X1 U4253 ( .A1(n5013), .A2(n5041), .ZN(n5219) );
  INV_X2 U4254 ( .A(n5984), .ZN(n5345) );
  NAND2_X4 U4255 ( .A1(n2587), .A2(n4887), .ZN(n4568) );
  NOR4_X4 U4256 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n5987)
         );
  INV_X4 U4257 ( .A(n3126), .ZN(n4885) );
  NAND2_X4 U4258 ( .A1(n3359), .A2(n3358), .ZN(n3464) );
  OAI21_X1 U4259 ( .B1(n4883), .B2(n2776), .A(n3227), .ZN(n4884) );
  INV_X1 U4260 ( .A(n5749), .ZN(n5751) );
  NOR3_X2 U4261 ( .A1(n4424), .A2(n5402), .A3(n4883), .ZN(n4369) );
  NOR2_X2 U4262 ( .A1(n3181), .A2(n3103), .ZN(n4333) );
  NAND2_X4 U4263 ( .A1(n3323), .A2(n2681), .ZN(n3324) );
  AND2_X4 U4264 ( .A1(\wb/dsize_reg/z2 [21]), .A2(n3178), .ZN(n3136) );
  INV_X1 U4265 ( .A(n4773), .ZN(n4430) );
  AOI221_X2 U4266 ( .B1(n5847), .B2(n5846), .C1(n5845), .C2(n5846), .A(n5844), 
        .ZN(n5848) );
  INV_X8 U4267 ( .A(n4135), .ZN(n3147) );
  INV_X2 U4268 ( .A(n5346), .ZN(n5352) );
  NAND2_X1 U4269 ( .A1(n5346), .A2(n3231), .ZN(n5348) );
  NAND2_X1 U4270 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  XNOR2_X1 U4271 ( .A(n5346), .B(n3221), .ZN(n4595) );
  NOR4_X1 U4272 ( .A1(n4839), .A2(n5218), .A3(n5845), .A4(n5832), .ZN(n4844)
         );
  NOR3_X1 U4273 ( .A1(n4767), .A2(n4766), .A3(n5845), .ZN(n4768) );
  NOR4_X2 U4274 ( .A1(n5219), .A2(n5218), .A3(n5845), .A4(n5217), .ZN(n5220)
         );
  NOR3_X1 U4275 ( .A1(n3091), .A2(n6336), .A3(n3173), .ZN(n3950) );
  NOR2_X1 U4276 ( .A1(n6327), .A2(n3091), .ZN(n4009) );
  NOR3_X1 U4277 ( .A1(n3091), .A2(n6335), .A3(n3173), .ZN(n3958) );
  NOR3_X1 U4278 ( .A1(n3180), .A2(n6340), .A3(n3146), .ZN(n5146) );
  NOR2_X1 U4279 ( .A1(n6330), .A2(n3091), .ZN(n3996) );
  NOR3_X1 U4280 ( .A1(n3091), .A2(n6308), .A3(n3173), .ZN(n4127) );
  NOR3_X1 U4281 ( .A1(n3172), .A2(n6319), .A3(n3087), .ZN(n4052) );
  INV_X2 U4282 ( .A(n5997), .ZN(n5824) );
  NOR2_X2 U4283 ( .A1(n2666), .A2(n3073), .ZN(n4015) );
  NAND3_X2 U4284 ( .A1(n4360), .A2(n4359), .A3(n4577), .ZN(n4362) );
  NOR2_X2 U4285 ( .A1(zeroExt_2), .A2(n3030), .ZN(n3137) );
  NAND3_X1 U4286 ( .A1(n5836), .A2(n5890), .A3(n5889), .ZN(n5852) );
  NAND2_X1 U4287 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  NAND3_X1 U4288 ( .A1(n5843), .A2(n5889), .A3(n5842), .ZN(n5847) );
  NOR2_X1 U4289 ( .A1(n4104), .A2(n3232), .ZN(n4105) );
  NOR2_X4 U4290 ( .A1(n3139), .A2(n6314), .ZN(n3138) );
  XNOR2_X1 U4291 ( .A(n6274), .B(n3692), .ZN(n3693) );
  NAND2_X1 U4292 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  INV_X2 U4293 ( .A(n6274), .ZN(n3331) );
  INV_X2 U4294 ( .A(n4276), .ZN(n3991) );
  INV_X1 U4295 ( .A(n5996), .ZN(n5797) );
  AOI21_X1 U4296 ( .B1(n5632), .B2(n3226), .A(n5633), .ZN(n5637) );
  NAND2_X1 U4297 ( .A1(n5633), .A2(n3231), .ZN(n5635) );
  NOR3_X2 U4298 ( .A1(n5965), .A2(n5966), .A3(n3128), .ZN(n3140) );
  AOI22_X1 U4299 ( .A1(n6029), .A2(n5479), .B1(n6005), .B2(n6068), .ZN(n5486)
         );
  NOR3_X2 U4300 ( .A1(n6051), .A2(n6068), .A3(n6064), .ZN(n6053) );
  OAI21_X1 U4301 ( .B1(n5239), .B2(n5470), .A(n5242), .ZN(n5240) );
  INV_X2 U4302 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U4303 ( .A1(n3790), .A2(n3789), .ZN(n3795) );
  NOR2_X1 U4304 ( .A1(n3619), .A2(n3618), .ZN(n3624) );
  XNOR2_X1 U4305 ( .A(n3507), .B(n3506), .ZN(n3510) );
  NAND2_X1 U4306 ( .A1(n3496), .A2(n3495), .ZN(n3497) );
  NAND3_X1 U4307 ( .A1(n3496), .A2(n3456), .A3(n3495), .ZN(n3367) );
  NAND3_X1 U4308 ( .A1(n3766), .A2(iAddr[12]), .A3(iAddr[11]), .ZN(n3767) );
  NAND2_X4 U4309 ( .A1(n3766), .A2(iAddr[11]), .ZN(n3672) );
  NAND2_X1 U4310 ( .A1(reg31Val_3[1]), .A2(n2953), .ZN(n3511) );
  NAND2_X2 U4311 ( .A1(n5042), .A2(n5044), .ZN(n4571) );
  AOI22_X1 U4312 ( .A1(n4129), .A2(n2608), .B1(n4524), .B2(memAddr[27]), .ZN(
        n4130) );
  NAND2_X1 U4313 ( .A1(n4129), .A2(n2654), .ZN(n4313) );
  NAND2_X1 U4314 ( .A1(n4129), .A2(n2660), .ZN(n4175) );
  NAND2_X1 U4315 ( .A1(n4129), .A2(n2658), .ZN(n4199) );
  NAND2_X1 U4316 ( .A1(n4129), .A2(n3021), .ZN(n4304) );
  NAND2_X1 U4317 ( .A1(n4129), .A2(n2655), .ZN(n4251) );
  NAND2_X1 U4318 ( .A1(n4129), .A2(n2653), .ZN(n4232) );
  NAND2_X1 U4319 ( .A1(n4129), .A2(n2659), .ZN(n4163) );
  NOR2_X1 U4320 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  NOR2_X1 U4321 ( .A1(n5977), .A2(n2718), .ZN(n5541) );
  INV_X2 U4322 ( .A(n4635), .ZN(n3998) );
  XNOR2_X1 U4323 ( .A(n5574), .B(n5618), .ZN(n5613) );
  NOR3_X1 U4324 ( .A1(n5701), .A2(n5700), .A3(n3157), .ZN(n5702) );
  NOR3_X1 U4325 ( .A1(n3062), .A2(n5004), .A3(n4975), .ZN(n4937) );
  NOR2_X1 U4326 ( .A1(n3062), .A2(n4948), .ZN(n4952) );
  OAI21_X1 U4327 ( .B1(n5701), .B2(n5700), .A(n3216), .ZN(n4979) );
  NOR3_X1 U4328 ( .A1(n3062), .A2(n5670), .A3(n4735), .ZN(n5271) );
  OAI21_X2 U4329 ( .B1(n5908), .B2(n5700), .A(n3216), .ZN(n5282) );
  INV_X8 U4330 ( .A(n5700), .ZN(n4929) );
  NAND3_X2 U4331 ( .A1(n3059), .A2(n5642), .A3(n5400), .ZN(n4659) );
  NAND2_X1 U4332 ( .A1(n4818), .A2(n4558), .ZN(n5042) );
  INV_X16 U4333 ( .A(n3236), .ZN(n3235) );
  INV_X8 U4334 ( .A(n4607), .ZN(n4661) );
  NOR2_X2 U4335 ( .A1(n4766), .A2(n5839), .ZN(n4678) );
  NOR2_X2 U4336 ( .A1(n5839), .A2(n2714), .ZN(n5821) );
  NOR2_X2 U4337 ( .A1(n5839), .A2(n5791), .ZN(n5794) );
  AOI22_X1 U4338 ( .A1(n4129), .A2(n2610), .B1(n4524), .B2(memAddr[23]), .ZN(
        n3953) );
  NAND2_X1 U4339 ( .A1(n4129), .A2(n2656), .ZN(n4378) );
  AOI22_X1 U4340 ( .A1(n4129), .A2(n2609), .B1(n4524), .B2(memAddr[26]), .ZN(
        n4124) );
  NAND2_X4 U4341 ( .A1(n4404), .A2(n4403), .ZN(n4408) );
  NAND4_X2 U4342 ( .A1(n5754), .A2(n5755), .A3(n5105), .A4(n5249), .ZN(n5108)
         );
  NOR3_X1 U4343 ( .A1(n3988), .A2(n3987), .A3(n4277), .ZN(n3994) );
  INV_X4 U4344 ( .A(n3067), .ZN(n4098) );
  NAND3_X2 U4345 ( .A1(n5400), .A2(n3059), .A3(n4673), .ZN(n5916) );
  NAND3_X2 U4346 ( .A1(n4197), .A2(n4196), .A3(n4195), .ZN(n4201) );
  NAND3_X1 U4347 ( .A1(n4533), .A2(n4153), .A3(n3178), .ZN(n4534) );
  NAND4_X1 U4348 ( .A1(n3243), .A2(n3178), .A3(n4153), .A4(
        \wb/dsize_reg/z2 [17]), .ZN(n4177) );
  NAND3_X2 U4349 ( .A1(n4153), .A2(\wb/dsize_reg/z2 [23]), .A3(n3167), .ZN(
        n3923) );
  NAND2_X4 U4350 ( .A1(n3114), .A2(n3084), .ZN(n4154) );
  NAND2_X4 U4351 ( .A1(n5679), .A2(n4616), .ZN(n5672) );
  OAI221_X4 U4352 ( .B1(n6571), .B2(n3155), .C1(n3185), .C2(n4505), .A(n4504), 
        .ZN(n5679) );
  NAND2_X4 U4353 ( .A1(n5189), .A2(n4445), .ZN(n4935) );
  OAI221_X4 U4354 ( .B1(n3185), .B2(n4654), .C1(n6570), .C2(n3155), .A(n4653), 
        .ZN(n5189) );
  XNOR2_X1 U4355 ( .A(n4914), .B(n4935), .ZN(n5328) );
  NOR3_X1 U4356 ( .A1(n4950), .A2(n4935), .A3(n4975), .ZN(n4936) );
  XNOR2_X1 U4357 ( .A(n3702), .B(n2821), .ZN(n3703) );
  XNOR2_X1 U4358 ( .A(n3690), .B(n2682), .ZN(n3691) );
  XNOR2_X1 U4359 ( .A(n3694), .B(n2700), .ZN(n3695) );
  XNOR2_X1 U4360 ( .A(n3717), .B(n3716), .ZN(n3718) );
  INV_X2 U4361 ( .A(n3817), .ZN(n3818) );
  NOR2_X2 U4362 ( .A1(n6260), .A2(n3817), .ZN(n3326) );
  XNOR2_X1 U4363 ( .A(n6194), .B(n2583), .ZN(n3529) );
  NOR2_X1 U4364 ( .A1(n6194), .A2(n2583), .ZN(n3513) );
  NAND2_X1 U4365 ( .A1(n6194), .A2(n2582), .ZN(n3522) );
  OAI211_X4 U4366 ( .C1(n3563), .C2(n3143), .A(n3562), .B(n3561), .ZN(
        iAddr[10]) );
  NAND2_X4 U4367 ( .A1(n4165), .A2(n3173), .ZN(n4639) );
  OAI211_X4 U4368 ( .C1(n3658), .C2(n3143), .A(n3656), .B(n3655), .ZN(
        iAddr[29]) );
  NAND2_X4 U4369 ( .A1(n3427), .A2(n3425), .ZN(n3378) );
  NAND2_X4 U4370 ( .A1(n3411), .A2(n3414), .ZN(n3427) );
  NAND2_X4 U4371 ( .A1(n3064), .A2(n3054), .ZN(n4104) );
  NAND2_X4 U4372 ( .A1(n3485), .A2(n3487), .ZN(n3475) );
  NAND2_X4 U4373 ( .A1(n3483), .A2(n3367), .ZN(n3487) );
  NAND2_X4 U4374 ( .A1(n3813), .A2(n3802), .ZN(n3805) );
  NAND3_X2 U4375 ( .A1(n5526), .A2(n5397), .A3(n4605), .ZN(n5036) );
  NAND3_X2 U4376 ( .A1(n5400), .A2(n4802), .A3(n5038), .ZN(n5372) );
  OAI211_X2 U4377 ( .C1(n4598), .C2(n5647), .A(n4599), .B(n5339), .ZN(n5526)
         );
  INV_X1 U4378 ( .A(n5638), .ZN(n5325) );
  OAI21_X1 U4379 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n5641) );
  NAND2_X4 U4380 ( .A1(n4567), .A2(n2587), .ZN(n4569) );
  INV_X2 U4381 ( .A(n4262), .ZN(n4050) );
  XNOR2_X1 U4382 ( .A(n5344), .B(n5343), .ZN(n5984) );
  INV_X2 U4383 ( .A(n5343), .ZN(n4603) );
  NAND3_X2 U4384 ( .A1(n4263), .A2(n4262), .A3(n3243), .ZN(n4266) );
  NAND2_X4 U4385 ( .A1(n5770), .A2(n5769), .ZN(n6049) );
  NAND2_X1 U4386 ( .A1(n5302), .A2(n5127), .ZN(n5129) );
  NAND2_X4 U4387 ( .A1(n5505), .A2(n5302), .ZN(n6024) );
  NOR3_X1 U4388 ( .A1(n5270), .A2(n3110), .A3(n5269), .ZN(n5273) );
  INV_X16 U4389 ( .A(n3218), .ZN(n3216) );
  NAND2_X4 U4390 ( .A1(n3218), .A2(n5082), .ZN(n5306) );
  INV_X8 U4391 ( .A(n5688), .ZN(n3218) );
  INV_X4 U4392 ( .A(n6492), .ZN(n6396) );
  OAI22_X2 U4393 ( .A1(n2837), .A2(n6426), .B1(n6421), .B2(n6436), .ZN(n6391)
         );
  NAND3_X1 U4394 ( .A1(n4511), .A2(n4319), .A3(n2997), .ZN(regWrData[12]) );
  AOI21_X1 U4395 ( .B1(n5065), .B2(n5465), .A(n5064), .ZN(n5066) );
  NAND2_X4 U4396 ( .A1(n5081), .A2(n5661), .ZN(n5705) );
  NAND4_X4 U4397 ( .A1(n4956), .A2(n4955), .A3(n4954), .A4(n4953), .ZN(n5509)
         );
  NAND4_X4 U4398 ( .A1(n4460), .A2(n4459), .A3(n4458), .A4(n4457), .ZN(n4950)
         );
  OAI21_X1 U4399 ( .B1(n4836), .B2(n3230), .A(n3227), .ZN(n4834) );
  NOR2_X1 U4400 ( .A1(n5790), .A2(n4836), .ZN(n4433) );
  INV_X8 U4401 ( .A(n4836), .ZN(n4846) );
  NAND2_X4 U4402 ( .A1(n5571), .A2(n4666), .ZN(n5666) );
  XNOR2_X1 U4403 ( .A(n4896), .B(n4895), .ZN(n5989) );
  OAI21_X1 U4404 ( .B1(n4895), .B2(n4892), .A(n4801), .ZN(n4804) );
  MUX2_X1 U4405 ( .A(n2961), .B(n3904), .S(n3162), .Z(n2015) );
  XNOR2_X1 U4406 ( .A(iAddr[29]), .B(n3805), .ZN(n3905) );
  OAI21_X1 U4407 ( .B1(n3461), .B2(n3568), .A(n3460), .ZN(n3469) );
  OAI21_X1 U4408 ( .B1(n3564), .B2(n3466), .A(n2894), .ZN(n3467) );
  NAND3_X2 U4409 ( .A1(n3779), .A2(iAddr[20]), .A3(iAddr[19]), .ZN(n3781) );
  INV_X8 U4410 ( .A(n3739), .ZN(n3761) );
  OAI211_X4 U4411 ( .C1(n3532), .C2(n3657), .A(n3531), .B(n3530), .ZN(iAddr[2]) );
  INV_X8 U4412 ( .A(n3069), .ZN(n5839) );
  NAND2_X4 U4413 ( .A1(n3315), .A2(n2700), .ZN(n3316) );
  NAND2_X4 U4414 ( .A1(n4605), .A2(n4604), .ZN(n5530) );
  NAND4_X2 U4415 ( .A1(n3140), .A2(n6059), .A3(n5999), .A4(n6070), .ZN(n6058)
         );
  NAND3_X2 U4416 ( .A1(n5992), .A2(n5991), .A3(n5990), .ZN(n5993) );
  AOI21_X4 U4417 ( .B1(n6108), .B2(n6107), .A(n6106), .ZN(n6111) );
  AOI211_X1 U4418 ( .C1(n3061), .C2(n5542), .A(n5541), .B(n5540), .ZN(n5550)
         );
  OAI21_X1 U4419 ( .B1(n3061), .B2(n3229), .A(n6008), .ZN(n5537) );
  NOR2_X1 U4420 ( .A1(n5995), .A2(n6063), .ZN(n5999) );
  NOR2_X1 U4421 ( .A1(n5377), .A2(n3061), .ZN(n4368) );
  INV_X4 U4422 ( .A(n6232), .ZN(n3158) );
  OAI22_X2 U4423 ( .A1(n4409), .A2(n4410), .B1(n4408), .B2(n3075), .ZN(n4411)
         );
  AOI21_X2 U4424 ( .B1(n5837), .B2(n5838), .A(n5839), .ZN(n4845) );
  NAND3_X1 U4425 ( .A1(n5846), .A2(n5838), .A3(n5837), .ZN(n5850) );
  NAND3_X1 U4426 ( .A1(n5398), .A2(n5397), .A3(n5642), .ZN(n5399) );
  NAND2_X1 U4427 ( .A1(n4795), .A2(n3117), .ZN(n4888) );
  INV_X8 U4428 ( .A(n4154), .ZN(n3169) );
  NOR2_X1 U4429 ( .A1(n6478), .A2(n3196), .ZN(\id_ex/N40 ) );
  NAND3_X1 U4430 ( .A1(n3847), .A2(n6402), .A3(n3846), .ZN(n2093) );
  NAND3_X1 U4431 ( .A1(n3845), .A2(n6402), .A3(n3844), .ZN(n2092) );
  NAND3_X1 U4432 ( .A1(n3843), .A2(n6402), .A3(n3842), .ZN(n2091) );
  NAND3_X1 U4433 ( .A1(n3841), .A2(n6402), .A3(n3840), .ZN(n2090) );
  NOR2_X1 U4434 ( .A1(n6401), .A2(n3053), .ZN(n3853) );
  NOR2_X1 U4435 ( .A1(n6401), .A2(n3044), .ZN(n3867) );
  NOR2_X1 U4436 ( .A1(n6401), .A2(n3045), .ZN(n3865) );
  NOR2_X1 U4437 ( .A1(n6401), .A2(n3046), .ZN(n3863) );
  NOR2_X1 U4438 ( .A1(n6401), .A2(n3047), .ZN(n3861) );
  NOR2_X1 U4439 ( .A1(n6401), .A2(n3048), .ZN(n3857) );
  NOR2_X1 U4440 ( .A1(n6401), .A2(n3049), .ZN(n3855) );
  NOR2_X1 U4441 ( .A1(n6401), .A2(n3050), .ZN(n3851) );
  NOR2_X1 U4442 ( .A1(n6401), .A2(n3051), .ZN(n3859) );
  OAI211_X1 U4443 ( .C1(n6527), .C2(n3849), .A(n6402), .B(n3848), .ZN(n2094)
         );
  OAI221_X1 U4444 ( .B1(n6553), .B2(n3849), .C1(n6605), .C2(n3193), .A(n6402), 
        .ZN(n2089) );
  OAI221_X1 U4445 ( .B1(n2579), .B2(n3903), .C1(n2628), .C2(n3193), .A(n3839), 
        .ZN(n2088) );
  XNOR2_X2 U4446 ( .A(rd_2[1]), .B(n2579), .ZN(n6501) );
  NAND2_X4 U4447 ( .A1(n3679), .A2(n3789), .ZN(n3800) );
  NAND2_X4 U4448 ( .A1(n3435), .A2(n3410), .ZN(n3610) );
  NAND2_X4 U4449 ( .A1(n3375), .A2(n3472), .ZN(n3602) );
  NAND2_X4 U4450 ( .A1(n5080), .A2(n5661), .ZN(n5700) );
  NAND2_X4 U4451 ( .A1(n4357), .A2(n3177), .ZN(n4390) );
  OAI211_X2 U4452 ( .C1(n5650), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5652)
         );
  NAND2_X4 U4453 ( .A1(n6060), .A2(n6059), .ZN(n6074) );
  NAND2_X4 U4454 ( .A1(n4911), .A2(n4914), .ZN(n5395) );
  NOR2_X1 U4455 ( .A1(n3801), .A2(n3800), .ZN(n3803) );
  XOR2_X1 U4456 ( .A(n6189), .B(n2583), .Z(n3751) );
  NOR2_X1 U4457 ( .A1(n6189), .A2(n2583), .ZN(n3745) );
  NAND3_X2 U4458 ( .A1(n3761), .A2(iAddr[10]), .A3(iAddr[9]), .ZN(n3762) );
  NAND2_X4 U4459 ( .A1(n3319), .A2(n2821), .ZN(n3320) );
  NAND2_X4 U4460 ( .A1(n2586), .A2(n2688), .ZN(n3732) );
  NAND2_X4 U4461 ( .A1(n3696), .A2(n2697), .ZN(n3698) );
  AOI21_X2 U4462 ( .B1(n5250), .B2(n5249), .A(n5248), .ZN(n5252) );
  XNOR2_X1 U4463 ( .A(n5401), .B(n5400), .ZN(n5991) );
  NAND3_X2 U4464 ( .A1(n5755), .A2(n5105), .A3(n5249), .ZN(n5048) );
  NAND2_X1 U4465 ( .A1(n5400), .A2(n5397), .ZN(n4794) );
  NAND3_X1 U4466 ( .A1(n4838), .A2(n5392), .A3(n5368), .ZN(n4428) );
  XNOR2_X1 U4467 ( .A(n5392), .B(n3222), .ZN(n4555) );
  INV_X8 U4468 ( .A(n4439), .ZN(n3144) );
  NAND2_X4 U4469 ( .A1(n5508), .A2(n4445), .ZN(n5494) );
  OAI221_X4 U4470 ( .B1(n6568), .B2(n3155), .C1(n3185), .C2(n4586), .A(n4585), 
        .ZN(n5508) );
  NOR4_X4 U4471 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6083)
         );
  NAND2_X4 U4472 ( .A1(n2849), .A2(n5032), .ZN(n4802) );
  NAND2_X4 U4473 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  INV_X32 U4474 ( .A(n3146), .ZN(n4357) );
  NAND4_X2 U4475 ( .A1(n6496), .A2(n6497), .A3(valid_2), .A4(n6498), .ZN(n6478) );
  AOI211_X2 U4476 ( .C1(op0_1), .C2(n6415), .A(n6416), .B(n6417), .ZN(n6414)
         );
  NOR3_X2 U4477 ( .A1(n6418), .A2(n6592), .A3(n2871), .ZN(n6417) );
  NOR4_X2 U4478 ( .A1(n6499), .A2(n6500), .A3(n6501), .A4(n6502), .ZN(n6498)
         );
  NAND4_X2 U4479 ( .A1(n6386), .A2(n6593), .A3(n6317), .A4(n6129), .ZN(n6418)
         );
  NOR2_X2 U4480 ( .A1(n3197), .A2(n6591), .ZN(n6129) );
  AOI21_X1 U4481 ( .B1(n3226), .B2(n5424), .A(n5423), .ZN(n5425) );
  NOR2_X1 U4482 ( .A1(n5423), .A2(n5705), .ZN(n4980) );
  NAND3_X1 U4483 ( .A1(n5644), .A2(n5647), .A3(n5339), .ZN(n5340) );
  NAND3_X1 U4484 ( .A1(n5325), .A2(n5647), .A3(n5339), .ZN(n5327) );
  NAND2_X4 U4485 ( .A1(n5647), .A2(n5339), .ZN(n4584) );
  NAND2_X4 U4486 ( .A1(n5444), .A2(n4445), .ZN(n5423) );
  NAND4_X1 U4487 ( .A1(n2850), .A2(n3065), .A3(n3234), .A4(n3177), .ZN(n4149)
         );
  NAND4_X1 U4488 ( .A1(n3024), .A2(n3065), .A3(n3234), .A4(n3167), .ZN(n4156)
         );
  NAND2_X1 U4489 ( .A1(n3065), .A2(n3234), .ZN(n3984) );
  NOR2_X1 U4490 ( .A1(n3065), .A2(n3233), .ZN(n4028) );
  NAND2_X4 U4491 ( .A1(n2585), .A2(n2691), .ZN(n3690) );
  NAND2_X4 U4492 ( .A1(n3704), .A2(n2825), .ZN(n3706) );
  NAND3_X2 U4493 ( .A1(n5125), .A2(n5126), .A3(n5124), .ZN(n5302) );
  NAND2_X4 U4494 ( .A1(n4355), .A2(n3177), .ZN(n4394) );
  NAND2_X4 U4495 ( .A1(n5047), .A2(n5465), .ZN(n5249) );
  NAND2_X4 U4496 ( .A1(n5017), .A2(n3116), .ZN(n5921) );
  AOI22_X1 U4497 ( .A1(n5947), .A2(n5802), .B1(n6005), .B2(n6063), .ZN(n5049)
         );
  NAND2_X1 U4498 ( .A1(n2895), .A2(n3069), .ZN(n5943) );
  NAND3_X1 U4499 ( .A1(n3069), .A2(n4769), .A3(n4768), .ZN(n4772) );
  NAND3_X1 U4500 ( .A1(n5751), .A2(n3069), .A3(n3127), .ZN(n5752) );
  NAND2_X4 U4501 ( .A1(n5820), .A2(n3069), .ZN(n5465) );
  NAND3_X1 U4502 ( .A1(n3159), .A2(memAddr[17]), .A3(n4098), .ZN(n4100) );
  NAND3_X1 U4503 ( .A1(n3067), .A2(n2651), .A3(n3159), .ZN(n4099) );
  NAND3_X1 U4504 ( .A1(n3067), .A2(n2652), .A3(n3159), .ZN(n4531) );
  NOR3_X1 U4505 ( .A1(n3159), .A2(n2703), .A3(n4098), .ZN(n3990) );
  NOR4_X1 U4506 ( .A1(n3984), .A2(n4098), .A3(n6331), .A4(n3159), .ZN(n3985)
         );
  NAND3_X1 U4507 ( .A1(n3067), .A2(n6367), .A3(n3159), .ZN(n4360) );
  NAND3_X1 U4508 ( .A1(n3067), .A2(n6366), .A3(n3159), .ZN(n4328) );
  NOR2_X1 U4509 ( .A1(n6176), .A2(n3067), .ZN(n4083) );
  NAND2_X4 U4510 ( .A1(n4170), .A2(n3235), .ZN(n4439) );
  INV_X32 U4511 ( .A(n3147), .ZN(n3148) );
  NAND2_X4 U4512 ( .A1(n3159), .A2(n4098), .ZN(n4135) );
  NAND2_X4 U4513 ( .A1(n4355), .A2(n3167), .ZN(n4161) );
  NAND2_X4 U4514 ( .A1(n3167), .A2(n3233), .ZN(n4343) );
  NAND2_X4 U4515 ( .A1(n4357), .A2(n3168), .ZN(n4162) );
  INV_X16 U4516 ( .A(n3062), .ZN(n5080) );
  INV_X16 U4517 ( .A(n4950), .ZN(n5081) );
  INV_X32 U4518 ( .A(n3169), .ZN(n3167) );
  INV_X32 U4519 ( .A(n3174), .ZN(n3173) );
  INV_X4 U4520 ( .A(n6257), .ZN(n3300) );
  XNOR2_X2 U4521 ( .A(op0_3), .B(n3300), .ZN(n3301) );
  NOR2_X4 U4522 ( .A1(n3196), .A2(n6594), .ZN(n6137) );
  INV_X4 U4523 ( .A(n6421), .ZN(n6136) );
  NAND2_X2 U4524 ( .A1(n3194), .A2(n6316), .ZN(n6776) );
  INV_X4 U4525 ( .A(n6776), .ZN(n6135) );
  NAND4_X2 U4526 ( .A1(n6403), .A2(n6399), .A3(n6134), .A4(n6404), .ZN(n6402)
         );
  INV_X4 U4527 ( .A(n6388), .ZN(n6416) );
  INV_X4 U4528 ( .A(n6133), .ZN(\id_ex/N4 ) );
  NAND2_X2 U4529 ( .A1(n6444), .A2(n6588), .ZN(n3302) );
  INV_X4 U4530 ( .A(n6132), .ZN(n6433) );
  MUX2_X2 U4531 ( .A(n6603), .B(n6438), .S(n3193), .Z(n6427) );
  NAND2_X2 U4532 ( .A1(n3194), .A2(n6317), .ZN(n6774) );
  INV_X4 U4533 ( .A(n6774), .ZN(n6434) );
  MUX2_X2 U4534 ( .A(n6600), .B(n6443), .S(n3193), .Z(n6440) );
  INV_X4 U4535 ( .A(n6418), .ZN(n6138) );
  NAND2_X2 U4536 ( .A1(n3194), .A2(n6369), .ZN(n3849) );
  NAND2_X2 U4537 ( .A1(n3194), .A2(n2662), .ZN(n3303) );
  INV_X4 U4538 ( .A(n3303), .ZN(n6130) );
  NAND2_X2 U4539 ( .A1(n6594), .A2(n6130), .ZN(n6371) );
  INV_X4 U4540 ( .A(n6129), .ZN(n6372) );
  OAI22_X2 U4541 ( .A1(n6437), .A2(n3197), .B1(n6446), .B2(n6421), .ZN(n6383)
         );
  INV_X4 U4542 ( .A(n6127), .ZN(n6483) );
  NAND2_X2 U4543 ( .A1(n6444), .A2(n6130), .ZN(n6398) );
  INV_X4 U4544 ( .A(n2582), .ZN(n3305) );
  INV_X4 U4545 ( .A(n3717), .ZN(n3309) );
  INV_X4 U4546 ( .A(n6184), .ZN(n3716) );
  INV_X4 U4547 ( .A(n3310), .ZN(n3712) );
  INV_X4 U4548 ( .A(n3714), .ZN(n3311) );
  INV_X4 U4549 ( .A(n3690), .ZN(n3313) );
  INV_X4 U4550 ( .A(n3314), .ZN(n3692) );
  INV_X4 U4551 ( .A(n3694), .ZN(n3315) );
  INV_X4 U4552 ( .A(n3698), .ZN(n3317) );
  INV_X4 U4553 ( .A(n3702), .ZN(n3319) );
  INV_X4 U4554 ( .A(n3706), .ZN(n3321) );
  INV_X4 U4555 ( .A(n3710), .ZN(n3323) );
  INV_X4 U4556 ( .A(n3732), .ZN(n3325) );
  XNOR2_X2 U4557 ( .A(n3326), .B(n6159), .ZN(n3327) );
  MUX2_X2 U4558 ( .A(reg31Val_0[31]), .B(n3327), .S(n3282), .Z(n1915) );
  XNOR2_X2 U4559 ( .A(\mem/addImm/mux_map1/M1/M3/z2[31] ), .B(n6159), .ZN(
        n3388) );
  XNOR2_X2 U4560 ( .A(n6222), .B(n6260), .ZN(n3661) );
  INV_X4 U4561 ( .A(n3661), .ZN(n3386) );
  NAND2_X2 U4562 ( .A1(n2688), .A2(n2909), .ZN(n3653) );
  INV_X4 U4563 ( .A(n3653), .ZN(n3382) );
  NAND2_X2 U4564 ( .A1(n2696), .A2(n2910), .ZN(n3379) );
  XNOR2_X2 U4565 ( .A(n6217), .B(n6265), .ZN(n3444) );
  NAND2_X2 U4566 ( .A1(n2681), .A2(n2911), .ZN(n3428) );
  NAND2_X2 U4567 ( .A1(n3444), .A2(n3428), .ZN(n3329) );
  XNOR2_X2 U4568 ( .A(n6218), .B(n6264), .ZN(n3429) );
  INV_X4 U4569 ( .A(n3429), .ZN(n3328) );
  NAND2_X2 U4570 ( .A1(n3329), .A2(n3328), .ZN(n3422) );
  NAND2_X2 U4571 ( .A1(n3379), .A2(n3422), .ZN(n3637) );
  XNOR2_X2 U4572 ( .A(n6219), .B(n6263), .ZN(n3639) );
  INV_X4 U4573 ( .A(n3639), .ZN(n3380) );
  NAND2_X2 U4574 ( .A1(n2689), .A2(n2912), .ZN(n3426) );
  XNOR2_X2 U4575 ( .A(n6215), .B(n6267), .ZN(n3403) );
  XNOR2_X2 U4576 ( .A(n6214), .B(n6268), .ZN(n3580) );
  XNOR2_X2 U4577 ( .A(n6213), .B(n6269), .ZN(n3625) );
  NAND2_X2 U4578 ( .A1(n2697), .A2(n2913), .ZN(n3611) );
  NAND2_X2 U4579 ( .A1(n2700), .A2(n2998), .ZN(n3598) );
  XNOR2_X2 U4580 ( .A(n6208), .B(n6274), .ZN(n3397) );
  INV_X4 U4581 ( .A(n6208), .ZN(n3330) );
  NAND2_X2 U4582 ( .A1(n3331), .A2(n3330), .ZN(n3631) );
  XNOR2_X2 U4583 ( .A(n6209), .B(n6273), .ZN(n3343) );
  INV_X4 U4584 ( .A(n3343), .ZN(n3633) );
  INV_X4 U4585 ( .A(n3409), .ZN(n3599) );
  NAND2_X2 U4586 ( .A1(n2682), .A2(n2914), .ZN(n3393) );
  NAND2_X2 U4587 ( .A1(n3631), .A2(n3393), .ZN(n3332) );
  XNOR2_X2 U4588 ( .A(n6210), .B(n6272), .ZN(n3612) );
  NAND2_X2 U4589 ( .A1(n3612), .A2(n3611), .ZN(n3333) );
  XNOR2_X2 U4590 ( .A(n6211), .B(n6271), .ZN(n3614) );
  INV_X4 U4591 ( .A(n3614), .ZN(n3436) );
  OAI21_X4 U4592 ( .B1(n6211), .B2(n6271), .A(n3335), .ZN(n3585) );
  XNOR2_X2 U4593 ( .A(n6212), .B(n6270), .ZN(n3572) );
  INV_X4 U4594 ( .A(n3572), .ZN(n3593) );
  OAI21_X4 U4595 ( .B1(n6212), .B2(n6270), .A(n3336), .ZN(n3622) );
  NOR2_X4 U4596 ( .A1(n3625), .A2(n3337), .ZN(n3339) );
  NOR2_X4 U4597 ( .A1(n3339), .A2(n3338), .ZN(n3574) );
  XNOR2_X2 U4598 ( .A(n6216), .B(n6266), .ZN(n3417) );
  INV_X4 U4599 ( .A(n3417), .ZN(n3414) );
  NAND2_X2 U4600 ( .A1(n3593), .A2(n3436), .ZN(n3620) );
  INV_X4 U4601 ( .A(n3403), .ZN(n3440) );
  INV_X4 U4602 ( .A(n3612), .ZN(n3606) );
  INV_X4 U4603 ( .A(n3580), .ZN(n3577) );
  INV_X4 U4604 ( .A(n3625), .ZN(n3405) );
  XNOR2_X2 U4605 ( .A(n6207), .B(n6275), .ZN(n3478) );
  INV_X4 U4606 ( .A(n3539), .ZN(n3451) );
  NAND2_X2 U4607 ( .A1(n2710), .A2(n2915), .ZN(n3347) );
  INV_X4 U4608 ( .A(n3755), .ZN(n3345) );
  XNOR2_X2 U4609 ( .A(reg31Val_3[1]), .B(n6193), .ZN(n3752) );
  NAND4_X2 U4610 ( .A1(n3514), .A2(n3347), .A3(n3511), .A4(n3512), .ZN(n3346)
         );
  INV_X4 U4611 ( .A(n3346), .ZN(n3352) );
  INV_X4 U4612 ( .A(n3347), .ZN(n3515) );
  XNOR2_X2 U4613 ( .A(n6195), .B(n6189), .ZN(n3524) );
  INV_X4 U4614 ( .A(n3524), .ZN(n3348) );
  NAND2_X2 U4615 ( .A1(n3348), .A2(n3522), .ZN(n3349) );
  INV_X4 U4616 ( .A(n3349), .ZN(n3516) );
  INV_X4 U4617 ( .A(n3517), .ZN(n3350) );
  OAI21_X4 U4618 ( .B1(n3352), .B2(n3351), .A(n2904), .ZN(n3538) );
  NAND2_X2 U4619 ( .A1(n2669), .A2(n2951), .ZN(n3448) );
  NAND2_X2 U4620 ( .A1(n3542), .A2(n3448), .ZN(n3533) );
  INV_X4 U4621 ( .A(n3533), .ZN(n3353) );
  NAND2_X2 U4622 ( .A1(n2671), .A2(n2952), .ZN(n3454) );
  INV_X4 U4623 ( .A(n3474), .ZN(n3370) );
  XNOR2_X2 U4624 ( .A(n6200), .B(n6185), .ZN(n3547) );
  XNOR2_X2 U4625 ( .A(n6204), .B(n6183), .ZN(n3463) );
  NAND2_X2 U4626 ( .A1(n2631), .A2(n2896), .ZN(n3460) );
  NAND2_X2 U4627 ( .A1(n3716), .A2(n2916), .ZN(n3504) );
  INV_X4 U4628 ( .A(n3504), .ZN(n3355) );
  NAND2_X2 U4629 ( .A1(n6202), .A2(n6279), .ZN(n3356) );
  XNOR2_X2 U4630 ( .A(n6203), .B(n6278), .ZN(n3506) );
  INV_X4 U4631 ( .A(n3506), .ZN(n3357) );
  INV_X4 U4632 ( .A(n3461), .ZN(n3354) );
  OAI21_X4 U4633 ( .B1(n3355), .B2(n3505), .A(n3354), .ZN(n3462) );
  NAND2_X2 U4634 ( .A1(n3460), .A2(n3462), .ZN(n3466) );
  INV_X4 U4635 ( .A(n3466), .ZN(n3359) );
  XNOR2_X2 U4636 ( .A(n6201), .B(n6184), .ZN(n3565) );
  INV_X4 U4637 ( .A(n3565), .ZN(n3459) );
  NAND2_X2 U4638 ( .A1(n2698), .A2(n2917), .ZN(n3495) );
  INV_X4 U4639 ( .A(n3495), .ZN(n3360) );
  NAND2_X2 U4640 ( .A1(n2690), .A2(n2918), .ZN(n3458) );
  NAND3_X2 U4641 ( .A1(n3462), .A2(n3458), .A3(n3460), .ZN(n3362) );
  INV_X4 U4642 ( .A(n3463), .ZN(n3465) );
  AND2_X2 U4643 ( .A1(n3362), .A2(n3465), .ZN(n3363) );
  XNOR2_X2 U4644 ( .A(n6205), .B(n6277), .ZN(n3499) );
  INV_X4 U4645 ( .A(n3499), .ZN(n3365) );
  INV_X4 U4646 ( .A(n3366), .ZN(n3483) );
  NAND2_X2 U4647 ( .A1(n2684), .A2(n2920), .ZN(n3485) );
  INV_X4 U4648 ( .A(n3485), .ZN(n3368) );
  NAND2_X2 U4649 ( .A1(n2691), .A2(n2921), .ZN(n3375) );
  INV_X4 U4650 ( .A(n3375), .ZN(n3476) );
  XNOR2_X2 U4651 ( .A(n6199), .B(n6186), .ZN(n3553) );
  XNOR2_X2 U4652 ( .A(n6206), .B(n6276), .ZN(n3488) );
  INV_X4 U4653 ( .A(n3488), .ZN(n3373) );
  OAI21_X4 U4654 ( .B1(n3475), .B2(n3374), .A(n3373), .ZN(n3472) );
  NAND4_X2 U4655 ( .A1(n3377), .A2(n3376), .A3(n3600), .A4(n3602), .ZN(n3425)
         );
  NAND3_X4 U4656 ( .A1(n3379), .A2(n2692), .A3(n3423), .ZN(n3638) );
  NAND3_X4 U4657 ( .A1(n3637), .A2(n3380), .A3(n3638), .ZN(n3381) );
  OAI21_X4 U4658 ( .B1(n6219), .B2(n6263), .A(n3381), .ZN(n3645) );
  XNOR2_X2 U4659 ( .A(n6220), .B(n6262), .ZN(n3646) );
  NAND2_X2 U4660 ( .A1(n3646), .A2(n3653), .ZN(n3383) );
  NAND2_X2 U4661 ( .A1(n3383), .A2(n2870), .ZN(n3384) );
  OAI21_X4 U4662 ( .B1(n3385), .B2(n3384), .A(n2954), .ZN(n3660) );
  NAND2_X2 U4663 ( .A1(n3386), .A2(n3660), .ZN(n3807) );
  XNOR2_X2 U4664 ( .A(n3388), .B(n3387), .ZN(n3392) );
  NAND2_X2 U4665 ( .A1(n3161), .A2(n2999), .ZN(n3402) );
  INV_X4 U4666 ( .A(n3478), .ZN(n3601) );
  NAND2_X2 U4667 ( .A1(n3394), .A2(n3393), .ZN(n3396) );
  NAND2_X2 U4668 ( .A1(n3396), .A2(n3395), .ZN(n3630) );
  INV_X4 U4669 ( .A(n3396), .ZN(n3398) );
  NAND3_X2 U4670 ( .A1(n3142), .A2(n3630), .A3(n3399), .ZN(n3401) );
  NAND2_X2 U4671 ( .A1(n3214), .A2(n2771), .ZN(n3400) );
  NAND3_X2 U4672 ( .A1(n3402), .A2(n3401), .A3(n3400), .ZN(iAddr[16]) );
  INV_X4 U4673 ( .A(n3620), .ZN(n3406) );
  NAND3_X2 U4674 ( .A1(n3406), .A2(n3405), .A3(n3404), .ZN(n3413) );
  INV_X4 U4675 ( .A(n3619), .ZN(n3407) );
  INV_X4 U4676 ( .A(n3408), .ZN(n3435) );
  INV_X4 U4677 ( .A(n3415), .ZN(n3416) );
  NAND2_X2 U4678 ( .A1(n3161), .A2(n3000), .ZN(n3419) );
  NAND2_X2 U4679 ( .A1(n3215), .A2(n2966), .ZN(n3418) );
  OAI211_X2 U4680 ( .C1(n3421), .C2(n3420), .A(n3419), .B(n3418), .ZN(
        iAddr[24]) );
  OAI211_X2 U4681 ( .C1(n3444), .C2(n2881), .A(n3429), .B(n3428), .ZN(n3431)
         );
  NAND2_X2 U4682 ( .A1(n3214), .A2(n2968), .ZN(n3433) );
  NAND2_X2 U4683 ( .A1(n3434), .A2(n3433), .ZN(iAddr[26]) );
  NAND2_X2 U4684 ( .A1(n3435), .A2(n3599), .ZN(n3575) );
  XNOR2_X2 U4685 ( .A(n3440), .B(n3439), .ZN(n3443) );
  NAND2_X2 U4686 ( .A1(n3161), .A2(n3001), .ZN(n3442) );
  NAND2_X2 U4687 ( .A1(n3215), .A2(n2965), .ZN(n3441) );
  OAI211_X2 U4688 ( .C1(n3443), .C2(n3143), .A(n3442), .B(n3441), .ZN(
        iAddr[23]) );
  XNOR2_X2 U4689 ( .A(n2881), .B(n3444), .ZN(n3447) );
  NAND2_X2 U4690 ( .A1(n3161), .A2(n3002), .ZN(n3446) );
  NAND2_X2 U4691 ( .A1(n3215), .A2(n2967), .ZN(n3445) );
  OAI211_X2 U4692 ( .C1(n3447), .C2(n3143), .A(n3446), .B(n3445), .ZN(
        iAddr[25]) );
  NAND2_X2 U4693 ( .A1(n3215), .A2(n2962), .ZN(n3471) );
  INV_X4 U4694 ( .A(n3448), .ZN(n3450) );
  INV_X4 U4695 ( .A(n3449), .ZN(n3534) );
  NAND2_X2 U4696 ( .A1(n3450), .A2(n3534), .ZN(n3453) );
  NAND3_X4 U4697 ( .A1(n3451), .A2(n3534), .A3(n3538), .ZN(n3452) );
  NAND3_X4 U4698 ( .A1(n3454), .A2(n3453), .A3(n3452), .ZN(n3552) );
  INV_X4 U4699 ( .A(n3553), .ZN(n3455) );
  NAND2_X2 U4700 ( .A1(n3552), .A2(n3455), .ZN(n3556) );
  INV_X4 U4701 ( .A(n3547), .ZN(n3457) );
  OAI211_X2 U4702 ( .C1(n3469), .C2(n3468), .A(n3467), .B(n3142), .ZN(n3470)
         );
  INV_X4 U4703 ( .A(n3490), .ZN(n3477) );
  XNOR2_X2 U4704 ( .A(n3479), .B(n3478), .ZN(n3482) );
  NAND2_X2 U4705 ( .A1(n3659), .A2(n3003), .ZN(n3481) );
  NAND2_X2 U4706 ( .A1(n3215), .A2(n2770), .ZN(n3480) );
  OAI211_X2 U4707 ( .C1(n3482), .C2(n3143), .A(n3481), .B(n3480), .ZN(
        iAddr[15]) );
  NAND2_X2 U4708 ( .A1(n3659), .A2(n3004), .ZN(n3493) );
  NAND3_X2 U4709 ( .A1(n3142), .A2(n3490), .A3(n3489), .ZN(n3492) );
  NAND2_X2 U4710 ( .A1(n3214), .A2(n2769), .ZN(n3491) );
  NAND3_X2 U4711 ( .A1(n3493), .A2(n3492), .A3(n3491), .ZN(iAddr[14]) );
  XNOR2_X2 U4712 ( .A(n3500), .B(n3499), .ZN(n3503) );
  NAND2_X2 U4713 ( .A1(n3659), .A2(n3005), .ZN(n3502) );
  NAND2_X2 U4714 ( .A1(n3215), .A2(n2768), .ZN(n3501) );
  OAI211_X2 U4715 ( .C1(n3503), .C2(n3143), .A(n3502), .B(n3501), .ZN(
        iAddr[13]) );
  NAND2_X2 U4716 ( .A1(n3659), .A2(n3006), .ZN(n3509) );
  NAND2_X2 U4717 ( .A1(n3215), .A2(n2767), .ZN(n3508) );
  INV_X4 U4718 ( .A(n3513), .ZN(n3514) );
  NAND2_X2 U4719 ( .A1(n2897), .A2(n3514), .ZN(n3523) );
  XNOR2_X2 U4720 ( .A(n3518), .B(n3517), .ZN(n3521) );
  NAND2_X2 U4721 ( .A1(n3215), .A2(n3034), .ZN(n3519) );
  NAND2_X2 U4722 ( .A1(n3523), .A2(n3522), .ZN(n3525) );
  XNOR2_X2 U4723 ( .A(n3525), .B(n3524), .ZN(n3528) );
  NAND2_X2 U4724 ( .A1(n3215), .A2(n3035), .ZN(n3526) );
  XNOR2_X2 U4725 ( .A(n2897), .B(n3529), .ZN(n3532) );
  NAND2_X2 U4726 ( .A1(n3215), .A2(n2765), .ZN(n3530) );
  XNOR2_X2 U4727 ( .A(n3534), .B(n3533), .ZN(n3537) );
  NAND2_X2 U4728 ( .A1(n3659), .A2(n3007), .ZN(n3536) );
  NAND2_X2 U4729 ( .A1(n3215), .A2(n3036), .ZN(n3535) );
  OAI211_X2 U4730 ( .C1(n3537), .C2(n3657), .A(n3536), .B(n3535), .ZN(iAddr[6]) );
  NAND2_X2 U4731 ( .A1(n3659), .A2(n3008), .ZN(n3545) );
  NAND2_X2 U4732 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  NAND3_X2 U4733 ( .A1(n3142), .A2(n3542), .A3(n3541), .ZN(n3544) );
  NAND2_X2 U4734 ( .A1(n3215), .A2(n3037), .ZN(n3543) );
  INV_X4 U4735 ( .A(n3546), .ZN(n3548) );
  XNOR2_X2 U4736 ( .A(n3548), .B(n3547), .ZN(n3551) );
  NAND2_X2 U4737 ( .A1(n3161), .A2(n3009), .ZN(n3550) );
  NAND2_X2 U4738 ( .A1(n3213), .A2(n3038), .ZN(n3549) );
  OAI211_X2 U4739 ( .C1(n3551), .C2(n2580), .A(n3550), .B(n3549), .ZN(iAddr[8]) );
  NAND2_X2 U4740 ( .A1(n3659), .A2(n3010), .ZN(n3559) );
  INV_X4 U4741 ( .A(n3552), .ZN(n3554) );
  NAND2_X2 U4742 ( .A1(n3554), .A2(n3553), .ZN(n3555) );
  NAND2_X2 U4743 ( .A1(n3213), .A2(n3039), .ZN(n3557) );
  XNOR2_X2 U4744 ( .A(n2847), .B(n3560), .ZN(n3563) );
  NAND2_X2 U4745 ( .A1(n3161), .A2(n2624), .ZN(n3562) );
  NAND2_X2 U4746 ( .A1(n3212), .A2(n2766), .ZN(n3561) );
  NAND2_X2 U4747 ( .A1(n3161), .A2(n3011), .ZN(n3571) );
  INV_X4 U4748 ( .A(n3564), .ZN(n3566) );
  NAND2_X2 U4749 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  NAND3_X2 U4750 ( .A1(n3142), .A2(n3568), .A3(n3567), .ZN(n3570) );
  NAND2_X2 U4751 ( .A1(n3212), .A2(n3040), .ZN(n3569) );
  NAND2_X2 U4752 ( .A1(n2851), .A2(n3573), .ZN(n3576) );
  INV_X4 U4753 ( .A(n3578), .ZN(n3579) );
  NAND2_X2 U4754 ( .A1(n3161), .A2(n3012), .ZN(n3582) );
  NAND2_X2 U4755 ( .A1(n3214), .A2(n2964), .ZN(n3581) );
  OAI211_X2 U4756 ( .C1(n3584), .C2(n3583), .A(n3582), .B(n3581), .ZN(
        iAddr[22]) );
  NAND2_X2 U4757 ( .A1(n3161), .A2(n3013), .ZN(n3596) );
  INV_X4 U4758 ( .A(n3618), .ZN(n3588) );
  NAND4_X2 U4759 ( .A1(n3602), .A2(n3601), .A3(n3588), .A4(n3587), .ZN(n3589)
         );
  OAI21_X2 U4760 ( .B1(n3593), .B2(n3592), .A(n3591), .ZN(n3595) );
  NAND2_X2 U4761 ( .A1(n3214), .A2(n2775), .ZN(n3594) );
  NAND2_X2 U4762 ( .A1(n3161), .A2(n3014), .ZN(n3609) );
  NAND2_X2 U4763 ( .A1(n2857), .A2(n3603), .ZN(n3605) );
  OAI21_X2 U4764 ( .B1(n3606), .B2(n3605), .A(n3604), .ZN(n3608) );
  NAND2_X2 U4765 ( .A1(n3212), .A2(n2773), .ZN(n3607) );
  XNOR2_X2 U4766 ( .A(n3614), .B(n3613), .ZN(n3615) );
  NAND2_X2 U4767 ( .A1(n3214), .A2(n2774), .ZN(n3616) );
  NAND3_X4 U4768 ( .A1(n3617), .A2(n3616), .A3(n2880), .ZN(iAddr[19]) );
  XNOR2_X2 U4769 ( .A(n3626), .B(n3625), .ZN(n3629) );
  NAND2_X2 U4770 ( .A1(n3161), .A2(n3015), .ZN(n3628) );
  NAND2_X2 U4771 ( .A1(n3212), .A2(n2963), .ZN(n3627) );
  OAI211_X2 U4772 ( .C1(n3629), .C2(n3143), .A(n3628), .B(n3627), .ZN(
        iAddr[21]) );
  NAND2_X2 U4773 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  XNOR2_X2 U4774 ( .A(n3633), .B(n3632), .ZN(n3636) );
  NAND2_X2 U4775 ( .A1(n3161), .A2(n3016), .ZN(n3635) );
  NAND2_X2 U4776 ( .A1(n3214), .A2(n2772), .ZN(n3634) );
  OAI211_X2 U4777 ( .C1(n3636), .C2(n3143), .A(n3635), .B(n3634), .ZN(
        iAddr[17]) );
  NAND2_X2 U4778 ( .A1(n3638), .A2(n3637), .ZN(n3640) );
  XNOR2_X2 U4779 ( .A(n3640), .B(n3639), .ZN(n3643) );
  NAND2_X2 U4780 ( .A1(n3161), .A2(n3017), .ZN(n3642) );
  NAND2_X2 U4781 ( .A1(n3213), .A2(n2969), .ZN(n3641) );
  OAI211_X2 U4782 ( .C1(n3643), .C2(n3143), .A(n3642), .B(n3641), .ZN(
        iAddr[27]) );
  NAND2_X2 U4783 ( .A1(n3161), .A2(n3018), .ZN(n3651) );
  INV_X4 U4784 ( .A(n3646), .ZN(n3644) );
  NAND2_X2 U4785 ( .A1(n3647), .A2(n3646), .ZN(n3648) );
  NAND2_X2 U4786 ( .A1(n3212), .A2(n2970), .ZN(n3649) );
  NAND3_X2 U4787 ( .A1(n3651), .A2(n3650), .A3(n3649), .ZN(iAddr[28]) );
  NAND2_X2 U4788 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  XNOR2_X2 U4789 ( .A(n2870), .B(n3654), .ZN(n3658) );
  NAND2_X2 U4790 ( .A1(n3161), .A2(n3019), .ZN(n3656) );
  NAND2_X2 U4791 ( .A1(n3214), .A2(n2971), .ZN(n3655) );
  NAND2_X2 U4792 ( .A1(n3161), .A2(n3020), .ZN(n3809) );
  NAND2_X2 U4793 ( .A1(n3213), .A2(n2961), .ZN(n3808) );
  NAND2_X2 U4794 ( .A1(n3809), .A2(n3808), .ZN(n3665) );
  INV_X4 U4795 ( .A(n3660), .ZN(n3662) );
  NAND2_X2 U4796 ( .A1(n3662), .A2(n3661), .ZN(n3806) );
  INV_X4 U4797 ( .A(iAddr[28]), .ZN(n3666) );
  NAND2_X2 U4798 ( .A1(iAddr[13]), .A2(iAddr[14]), .ZN(n3669) );
  INV_X4 U4799 ( .A(iAddr[12]), .ZN(n3668) );
  NAND3_X4 U4800 ( .A1(n3673), .A2(iAddr[15]), .A3(n3734), .ZN(n3787) );
  NAND3_X2 U4801 ( .A1(iAddr[25]), .A2(iAddr[23]), .A3(n3772), .ZN(n3674) );
  INV_X4 U4802 ( .A(iAddr[26]), .ZN(n3798) );
  NAND2_X2 U4803 ( .A1(iAddr[24]), .A2(iAddr[16]), .ZN(n3788) );
  NOR3_X4 U4804 ( .A1(n3674), .A2(n3798), .A3(n3788), .ZN(n3679) );
  INV_X4 U4805 ( .A(iAddr[22]), .ZN(n3677) );
  INV_X4 U4806 ( .A(iAddr[18]), .ZN(n3774) );
  INV_X4 U4807 ( .A(iAddr[20]), .ZN(n3776) );
  NOR3_X4 U4808 ( .A1(n3675), .A2(n3774), .A3(n3776), .ZN(n3783) );
  INV_X4 U4809 ( .A(n3783), .ZN(n3676) );
  NOR3_X4 U4810 ( .A1(n3678), .A2(n3677), .A3(n3676), .ZN(n3789) );
  XNOR2_X2 U4811 ( .A(iAddr[31]), .B(n3682), .ZN(n3822) );
  NAND2_X2 U4812 ( .A1(not_trap_3), .A2(n3816), .ZN(n3759) );
  MUX2_X2 U4813 ( .A(n3029), .B(n3822), .S(n3163), .Z(n1918) );
  MUX2_X2 U4814 ( .A(reg31Val_0[12]), .B(n3686), .S(n3280), .Z(n1919) );
  MUX2_X2 U4815 ( .A(reg31Val_0[13]), .B(n3688), .S(n3280), .Z(n1920) );
  XNOR2_X2 U4816 ( .A(n6276), .B(n2585), .ZN(n3689) );
  MUX2_X2 U4817 ( .A(reg31Val_0[14]), .B(n3689), .S(n3280), .Z(n1926) );
  MUX2_X2 U4818 ( .A(reg31Val_0[15]), .B(n3691), .S(n3280), .Z(n1927) );
  MUX2_X2 U4819 ( .A(reg31Val_0[16]), .B(n3693), .S(n3280), .Z(n1928) );
  MUX2_X2 U4820 ( .A(reg31Val_0[17]), .B(n3695), .S(n3280), .Z(n1929) );
  MUX2_X2 U4821 ( .A(reg31Val_0[18]), .B(n3697), .S(n3280), .Z(n1930) );
  MUX2_X2 U4822 ( .A(reg31Val_0[19]), .B(n3699), .S(n3280), .Z(n1931) );
  MUX2_X2 U4823 ( .A(reg31Val_0[20]), .B(n3701), .S(n3280), .Z(n1932) );
  MUX2_X2 U4824 ( .A(reg31Val_0[21]), .B(n3703), .S(n3280), .Z(n1933) );
  MUX2_X2 U4825 ( .A(reg31Val_0[22]), .B(n3705), .S(n3281), .Z(n1934) );
  MUX2_X2 U4826 ( .A(reg31Val_0[23]), .B(n3707), .S(n3281), .Z(n1935) );
  XNOR2_X2 U4827 ( .A(n6266), .B(n3708), .ZN(n3709) );
  MUX2_X2 U4828 ( .A(reg31Val_0[24]), .B(n3709), .S(n3281), .Z(n1936) );
  MUX2_X2 U4829 ( .A(reg31Val_0[25]), .B(n3711), .S(n3281), .Z(n1937) );
  MUX2_X2 U4830 ( .A(reg31Val_0[10]), .B(n3713), .S(n3281), .Z(n1938) );
  MUX2_X2 U4831 ( .A(reg31Val_0[11]), .B(n3715), .S(n3281), .Z(n1939) );
  MUX2_X2 U4832 ( .A(reg31Val_0[9]), .B(n3718), .S(n3281), .Z(n1940) );
  MUX2_X2 U4833 ( .A(reg31Val_0[7]), .B(n3720), .S(n3281), .Z(n1941) );
  XNOR2_X2 U4834 ( .A(n6185), .B(n3721), .ZN(n3722) );
  MUX2_X2 U4835 ( .A(reg31Val_0[8]), .B(n3722), .S(n3281), .Z(n1942) );
  NAND2_X2 U4836 ( .A1(n3745), .A2(n2852), .ZN(n3724) );
  XNOR2_X2 U4837 ( .A(n3724), .B(n2669), .ZN(n3723) );
  MUX2_X2 U4838 ( .A(reg31Val_0[5]), .B(n3723), .S(n3281), .Z(n1943) );
  MUX2_X2 U4839 ( .A(reg31Val_0[6]), .B(n3726), .S(n3281), .Z(n1944) );
  MUX2_X2 U4840 ( .A(n3037), .B(n3823), .S(n3163), .Z(n1947) );
  MUX2_X2 U4841 ( .A(reg31Val_0[26]), .B(n3728), .S(n3281), .Z(n1950) );
  MUX2_X2 U4842 ( .A(reg31Val_0[27]), .B(n3730), .S(n3281), .Z(n1952) );
  XNOR2_X2 U4843 ( .A(n6262), .B(n2586), .ZN(n3731) );
  MUX2_X2 U4844 ( .A(reg31Val_0[28]), .B(n3731), .S(n3281), .Z(n1954) );
  MUX2_X2 U4845 ( .A(reg31Val_0[29]), .B(n3733), .S(n3282), .Z(n1955) );
  INV_X4 U4846 ( .A(n3824), .ZN(n3735) );
  MUX2_X2 U4847 ( .A(n2962), .B(n3735), .S(n3163), .Z(n1958) );
  INV_X4 U4848 ( .A(iAddr[9]), .ZN(n3736) );
  XNOR2_X2 U4849 ( .A(n3736), .B(n3761), .ZN(n3826) );
  MUX2_X2 U4850 ( .A(n3040), .B(n3826), .S(n3163), .Z(n1961) );
  INV_X4 U4851 ( .A(iAddr[7]), .ZN(n3738) );
  INV_X4 U4852 ( .A(iAddr[8]), .ZN(n3737) );
  MUX2_X2 U4853 ( .A(n3038), .B(n2906), .S(n3163), .Z(n1964) );
  MUX2_X2 U4854 ( .A(n3039), .B(n3827), .S(n3163), .Z(n1967) );
  INV_X4 U4855 ( .A(iAddr[5]), .ZN(n3742) );
  INV_X4 U4856 ( .A(iAddr[6]), .ZN(n3741) );
  MUX2_X2 U4857 ( .A(n3036), .B(n2907), .S(n3163), .Z(n1970) );
  MUX2_X2 U4858 ( .A(reg31Val_0[4]), .B(n3746), .S(n3282), .Z(n1971) );
  MUX2_X2 U4859 ( .A(n3034), .B(n3828), .S(n3163), .Z(n1974) );
  MUX2_X2 U4860 ( .A(reg31Val_0[3]), .B(n3751), .S(n3282), .Z(n1975) );
  MUX2_X2 U4861 ( .A(n3035), .B(n2721), .S(n3162), .Z(n1978) );
  MUX2_X2 U4862 ( .A(n2765), .B(n3829), .S(n3162), .Z(n6756) );
  OAI22_X2 U4863 ( .A1(n6522), .A2(n3760), .B1(n3830), .B2(n3759), .ZN(n1986)
         );
  INV_X4 U4864 ( .A(n3758), .ZN(n3831) );
  OAI22_X2 U4865 ( .A1(n6523), .A2(n3760), .B1(n3831), .B2(n3759), .ZN(n1990)
         );
  MUX2_X2 U4866 ( .A(n3064), .B(n2635), .S(n3282), .Z(n6644) );
  MUX2_X2 U4867 ( .A(n3233), .B(link_3), .S(n3282), .Z(n1992) );
  NAND2_X2 U4868 ( .A1(n3761), .A2(iAddr[9]), .ZN(n3764) );
  MUX2_X2 U4869 ( .A(n2766), .B(n3922), .S(n3163), .Z(n1996) );
  MUX2_X2 U4870 ( .A(n2767), .B(n3920), .S(n3163), .Z(n1997) );
  XNOR2_X2 U4871 ( .A(n3767), .B(iAddr[13]), .ZN(n3919) );
  MUX2_X2 U4872 ( .A(n2768), .B(n3919), .S(n3163), .Z(n1998) );
  INV_X4 U4873 ( .A(n3767), .ZN(n3768) );
  NAND2_X2 U4874 ( .A1(n2876), .A2(iAddr[14]), .ZN(n3770) );
  INV_X4 U4875 ( .A(n3769), .ZN(n3918) );
  MUX2_X2 U4876 ( .A(n2769), .B(n3918), .S(n3163), .Z(n1999) );
  XNOR2_X2 U4877 ( .A(iAddr[15]), .B(n3770), .ZN(n3917) );
  MUX2_X2 U4878 ( .A(n2770), .B(n3917), .S(n3163), .Z(n2000) );
  INV_X4 U4879 ( .A(iAddr[16]), .ZN(n3771) );
  NAND2_X2 U4880 ( .A1(n3772), .A2(iAddr[16]), .ZN(n3782) );
  MUX2_X2 U4881 ( .A(n2771), .B(n3916), .S(n3163), .Z(n2001) );
  MUX2_X2 U4882 ( .A(n2772), .B(n3915), .S(n3163), .Z(n2002) );
  MUX2_X2 U4883 ( .A(n2773), .B(n3914), .S(n3162), .Z(n2003) );
  INV_X4 U4884 ( .A(n3777), .ZN(n3779) );
  INV_X4 U4885 ( .A(iAddr[19]), .ZN(n3778) );
  XNOR2_X2 U4886 ( .A(n3779), .B(n3778), .ZN(n3913) );
  MUX2_X2 U4887 ( .A(n2774), .B(n3913), .S(n3163), .Z(n2004) );
  MUX2_X2 U4888 ( .A(n2775), .B(n2984), .S(n3162), .Z(n2005) );
  XNOR2_X2 U4889 ( .A(iAddr[21]), .B(n3781), .ZN(n3912) );
  MUX2_X2 U4890 ( .A(n2963), .B(n3912), .S(n3162), .Z(n2006) );
  INV_X4 U4891 ( .A(n3782), .ZN(n3784) );
  INV_X4 U4892 ( .A(n3792), .ZN(n3785) );
  MUX2_X2 U4893 ( .A(n2964), .B(n3911), .S(n3162), .Z(n2007) );
  INV_X4 U4894 ( .A(iAddr[23]), .ZN(n3793) );
  XNOR2_X2 U4895 ( .A(n3785), .B(n3793), .ZN(n3910) );
  MUX2_X2 U4896 ( .A(n2965), .B(n3910), .S(n3162), .Z(n2008) );
  INV_X4 U4897 ( .A(iAddr[24]), .ZN(n3791) );
  MUX2_X2 U4898 ( .A(n2966), .B(n2760), .S(n3162), .Z(n2009) );
  INV_X4 U4899 ( .A(n3795), .ZN(n3797) );
  INV_X4 U4900 ( .A(iAddr[25]), .ZN(n3796) );
  XNOR2_X2 U4901 ( .A(n3797), .B(n3796), .ZN(n3909) );
  MUX2_X2 U4902 ( .A(n2967), .B(n3909), .S(n3162), .Z(n2010) );
  NAND2_X2 U4903 ( .A1(n3797), .A2(iAddr[25]), .ZN(n3799) );
  MUX2_X2 U4904 ( .A(n2968), .B(n3908), .S(n3162), .Z(n2011) );
  INV_X4 U4905 ( .A(iAddr[27]), .ZN(n3801) );
  XNOR2_X2 U4906 ( .A(n3813), .B(n3801), .ZN(n3907) );
  MUX2_X2 U4907 ( .A(n2969), .B(n3907), .S(n3162), .Z(n2012) );
  NAND2_X2 U4908 ( .A1(iAddr[28]), .A2(iAddr[27]), .ZN(n3811) );
  INV_X4 U4909 ( .A(n3811), .ZN(n3802) );
  INV_X4 U4910 ( .A(n3804), .ZN(n3906) );
  MUX2_X2 U4911 ( .A(n2970), .B(n3906), .S(n3162), .Z(n2013) );
  MUX2_X2 U4912 ( .A(n2971), .B(n3905), .S(n3162), .Z(n2014) );
  NAND3_X2 U4913 ( .A1(n3810), .A2(n3809), .A3(n3808), .ZN(iAddr[30]) );
  INV_X4 U4914 ( .A(iAddr[29]), .ZN(n3812) );
  XNOR2_X2 U4915 ( .A(n3815), .B(iAddr[30]), .ZN(n3904) );
  MUX2_X2 U4916 ( .A(n2722), .B(dSize[1]), .S(n3282), .Z(n2121) );
  MUX2_X2 U4917 ( .A(dSize[1]), .B(n2757), .S(n2623), .Z(n2122) );
  INV_X4 U4918 ( .A(n6313), .ZN(n4029) );
  MUX2_X2 U4919 ( .A(n4029), .B(dSize[0]), .S(n3282), .Z(n2124) );
  MUX2_X2 U4920 ( .A(dSize[0]), .B(n2758), .S(n2623), .Z(n2125) );
  MUX2_X2 U4921 ( .A(n3084), .B(fp_3), .S(n3282), .Z(n2128) );
  INV_X4 U4922 ( .A(n3816), .ZN(n3921) );
  MUX2_X2 U4923 ( .A(instruction[0]), .B(n2837), .S(n3166), .Z(n2139) );
  MUX2_X2 U4924 ( .A(instruction[2]), .B(n2871), .S(n3165), .Z(n2141) );
  MUX2_X2 U4925 ( .A(instruction[4]), .B(n2712), .S(n3166), .Z(n2143) );
  XNOR2_X2 U4926 ( .A(n6260), .B(n3818), .ZN(n3819) );
  MUX2_X2 U4927 ( .A(reg31Val_0[30]), .B(n3819), .S(n3282), .Z(n2174) );
  NAND2_X2 U4928 ( .A1(n6341), .A2(n3215), .ZN(\ex_mem/N242 ) );
  INV_X4 U4929 ( .A(n6449), .ZN(n3821) );
  INV_X4 U4930 ( .A(n6406), .ZN(n3820) );
  MUX2_X2 U4931 ( .A(n2725), .B(n2929), .S(n3193), .Z(n1916) );
  MUX2_X2 U4932 ( .A(n3822), .B(n2929), .S(n3921), .Z(n1917) );
  MUX2_X2 U4933 ( .A(n2726), .B(n2611), .S(n3193), .Z(n1945) );
  MUX2_X2 U4934 ( .A(n3823), .B(n2611), .S(n3166), .Z(n1946) );
  MUX2_X2 U4935 ( .A(n2727), .B(n2983), .S(n3193), .Z(n1956) );
  MUX2_X2 U4936 ( .A(n3824), .B(n6514), .S(n3165), .Z(n3825) );
  INV_X4 U4937 ( .A(n3825), .ZN(n1957) );
  MUX2_X2 U4938 ( .A(n2728), .B(n2612), .S(n3193), .Z(n1959) );
  MUX2_X2 U4939 ( .A(n3826), .B(n2612), .S(n3165), .Z(n1960) );
  MUX2_X2 U4940 ( .A(n2729), .B(n2613), .S(n3193), .Z(n1962) );
  MUX2_X2 U4941 ( .A(n2906), .B(n2613), .S(n3166), .Z(n1963) );
  MUX2_X2 U4942 ( .A(n2730), .B(n2614), .S(n3193), .Z(n1965) );
  MUX2_X2 U4943 ( .A(n3827), .B(n2614), .S(n3165), .Z(n1966) );
  MUX2_X2 U4944 ( .A(n2731), .B(n2615), .S(n3193), .Z(n1968) );
  MUX2_X2 U4945 ( .A(n2907), .B(n2615), .S(n3166), .Z(n1969) );
  MUX2_X2 U4946 ( .A(n2732), .B(n2616), .S(n3193), .Z(n1972) );
  MUX2_X2 U4947 ( .A(n3828), .B(n2616), .S(n3165), .Z(n1973) );
  MUX2_X2 U4948 ( .A(n2733), .B(n2617), .S(n3193), .Z(n1976) );
  MUX2_X2 U4949 ( .A(n2721), .B(n2617), .S(n3164), .Z(n1977) );
  MUX2_X2 U4950 ( .A(n2734), .B(n2930), .S(n3193), .Z(n1980) );
  MUX2_X2 U4951 ( .A(n3829), .B(n2930), .S(n3164), .Z(n1981) );
  MUX2_X2 U4952 ( .A(n2735), .B(n2618), .S(n3193), .Z(n6763) );
  MUX2_X2 U4953 ( .A(iAddr[1]), .B(n2618), .S(n3164), .Z(n6752) );
  MUX2_X2 U4954 ( .A(n2736), .B(n2619), .S(n3193), .Z(n6764) );
  MUX2_X2 U4955 ( .A(iAddr[0]), .B(n2619), .S(n3164), .Z(n6753) );
  NAND2_X2 U4956 ( .A1(n6424), .A2(n2837), .ZN(n3834) );
  NAND2_X2 U4957 ( .A1(n6423), .A2(n6132), .ZN(n3833) );
  NAND2_X2 U4958 ( .A1(n3197), .A2(n2787), .ZN(n3832) );
  NAND4_X2 U4959 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n6414), .ZN(n2018)
         );
  MUX2_X2 U4960 ( .A(n3021), .B(busB[31]), .S(n3193), .Z(n6701) );
  MUX2_X2 U4961 ( .A(n2812), .B(busB[30]), .S(n3193), .Z(n6702) );
  MUX2_X2 U4962 ( .A(n2815), .B(busB[29]), .S(n3192), .Z(n6703) );
  MUX2_X2 U4963 ( .A(n2816), .B(busB[28]), .S(n3193), .Z(n6704) );
  MUX2_X2 U4964 ( .A(n2608), .B(busB[27]), .S(n3192), .Z(n6705) );
  MUX2_X2 U4965 ( .A(n2609), .B(busB[26]), .S(n3192), .Z(n6706) );
  MUX2_X2 U4966 ( .A(n2817), .B(busB[25]), .S(n3193), .Z(n6707) );
  MUX2_X2 U4967 ( .A(n2607), .B(busB[24]), .S(n3193), .Z(n6708) );
  MUX2_X2 U4968 ( .A(n2610), .B(busB[23]), .S(n3192), .Z(n6709) );
  MUX2_X2 U4969 ( .A(n2818), .B(busB[22]), .S(n3192), .Z(n6710) );
  MUX2_X2 U4970 ( .A(n2814), .B(busB[21]), .S(n3192), .Z(n6711) );
  MUX2_X2 U4971 ( .A(n2819), .B(busB[20]), .S(n3192), .Z(n6712) );
  MUX2_X2 U4972 ( .A(n2820), .B(busB[19]), .S(n3192), .Z(n6713) );
  MUX2_X2 U4973 ( .A(n2606), .B(busB[18]), .S(n3192), .Z(n6714) );
  MUX2_X2 U4974 ( .A(n2651), .B(busB[17]), .S(n3192), .Z(n6715) );
  MUX2_X2 U4975 ( .A(n2813), .B(busB[16]), .S(n3192), .Z(n6716) );
  MUX2_X2 U4976 ( .A(n2653), .B(busB[15]), .S(n3192), .Z(n6717) );
  MUX2_X2 U4977 ( .A(n6366), .B(busB[14]), .S(n3192), .Z(n6718) );
  MUX2_X2 U4978 ( .A(n2637), .B(busB[13]), .S(n3192), .Z(n6719) );
  MUX2_X2 U4979 ( .A(n2654), .B(busB[12]), .S(n3192), .Z(n6720) );
  MUX2_X2 U4980 ( .A(n6367), .B(busB[11]), .S(n3192), .Z(n6721) );
  MUX2_X2 U4981 ( .A(n2634), .B(busB[10]), .S(n3191), .Z(n6722) );
  MUX2_X2 U4982 ( .A(n2677), .B(busB[9]), .S(n3192), .Z(n6723) );
  MUX2_X2 U4983 ( .A(n2638), .B(busB[8]), .S(n3191), .Z(n6724) );
  MUX2_X2 U4984 ( .A(n2655), .B(busB[7]), .S(n3192), .Z(n6725) );
  MUX2_X2 U4985 ( .A(n2656), .B(busB[6]), .S(n3191), .Z(n6726) );
  MUX2_X2 U4986 ( .A(n2672), .B(busB[5]), .S(n3192), .Z(n6727) );
  MUX2_X2 U4987 ( .A(n2657), .B(busB[4]), .S(n3191), .Z(n6728) );
  MUX2_X2 U4988 ( .A(n2658), .B(busB[3]), .S(n3192), .Z(n6729) );
  MUX2_X2 U4989 ( .A(n2659), .B(busB[2]), .S(n3188), .Z(n6730) );
  MUX2_X2 U4990 ( .A(n2660), .B(busB[1]), .S(n3191), .Z(n6731) );
  MUX2_X2 U4991 ( .A(n2652), .B(busB[0]), .S(n3192), .Z(n6732) );
  MUX2_X2 U4992 ( .A(n2639), .B(busA[31]), .S(n3190), .Z(n6669) );
  MUX2_X2 U4993 ( .A(n2640), .B(busA[30]), .S(n3189), .Z(n6670) );
  MUX2_X2 U4994 ( .A(n2674), .B(busA[29]), .S(n3188), .Z(n6671) );
  MUX2_X2 U4995 ( .A(n2675), .B(busA[28]), .S(n3191), .Z(n6672) );
  MUX2_X2 U4996 ( .A(n2676), .B(busA[27]), .S(n3192), .Z(n6673) );
  MUX2_X2 U4997 ( .A(n2799), .B(busA[26]), .S(n3191), .Z(n6674) );
  MUX2_X2 U4998 ( .A(n2800), .B(busA[25]), .S(n3191), .Z(n6675) );
  MUX2_X2 U4999 ( .A(n2801), .B(busA[24]), .S(n3191), .Z(n6676) );
  MUX2_X2 U5000 ( .A(n2802), .B(busA[23]), .S(n3191), .Z(n6677) );
  MUX2_X2 U5001 ( .A(n2803), .B(busA[22]), .S(n3191), .Z(n6678) );
  MUX2_X2 U5002 ( .A(n2804), .B(busA[21]), .S(n3191), .Z(n6679) );
  MUX2_X2 U5003 ( .A(n2805), .B(busA[20]), .S(n3191), .Z(n6680) );
  MUX2_X2 U5004 ( .A(n2806), .B(busA[19]), .S(n3191), .Z(n6681) );
  MUX2_X2 U5005 ( .A(n2807), .B(busA[18]), .S(n3191), .Z(n6682) );
  MUX2_X2 U5006 ( .A(n2792), .B(busA[17]), .S(n3191), .Z(n6683) );
  MUX2_X2 U5007 ( .A(n2599), .B(busA[16]), .S(n3191), .Z(n6684) );
  MUX2_X2 U5008 ( .A(n2808), .B(busA[15]), .S(n3191), .Z(n6685) );
  MUX2_X2 U5009 ( .A(n2641), .B(busA[14]), .S(n3191), .Z(n6686) );
  MUX2_X2 U5010 ( .A(n2642), .B(busA[13]), .S(n3191), .Z(n6687) );
  MUX2_X2 U5011 ( .A(n2643), .B(busA[12]), .S(n3191), .Z(n6688) );
  MUX2_X2 U5012 ( .A(n2644), .B(busA[11]), .S(n3190), .Z(n6689) );
  MUX2_X2 U5013 ( .A(n2645), .B(busA[10]), .S(n3190), .Z(n6690) );
  MUX2_X2 U5014 ( .A(n2600), .B(busA[9]), .S(n3190), .Z(n6691) );
  MUX2_X2 U5015 ( .A(n2793), .B(busA[8]), .S(n3190), .Z(n6692) );
  MUX2_X2 U5016 ( .A(n2794), .B(busA[7]), .S(n3190), .Z(n6693) );
  MUX2_X2 U5017 ( .A(n2795), .B(busA[6]), .S(n3190), .Z(n6694) );
  MUX2_X2 U5018 ( .A(n2791), .B(busA[5]), .S(n3190), .Z(n6695) );
  MUX2_X2 U5019 ( .A(n2796), .B(busA[4]), .S(n3190), .Z(n6696) );
  MUX2_X2 U5020 ( .A(n2809), .B(busA[3]), .S(n3190), .Z(n6697) );
  MUX2_X2 U5021 ( .A(n2646), .B(busA[2]), .S(n3190), .Z(n6698) );
  MUX2_X2 U5022 ( .A(n2647), .B(busA[1]), .S(n3190), .Z(n6699) );
  MUX2_X2 U5023 ( .A(n2648), .B(busA[0]), .S(n3190), .Z(n6700) );
  NAND2_X2 U5024 ( .A1(n6134), .A2(n2788), .ZN(n3836) );
  OAI221_X2 U5025 ( .B1(n6411), .B2(n3903), .C1(n2782), .C2(n3193), .A(n3836), 
        .ZN(n2083) );
  NAND2_X2 U5026 ( .A1(n3193), .A2(n2883), .ZN(n3873) );
  INV_X4 U5027 ( .A(n3873), .ZN(n6124) );
  NAND2_X2 U5028 ( .A1(n6124), .A2(n2788), .ZN(n3837) );
  OAI221_X2 U5029 ( .B1(n6410), .B2(n3903), .C1(n2593), .C2(n3193), .A(n3837), 
        .ZN(n2084) );
  NAND2_X2 U5030 ( .A1(n3194), .A2(n2884), .ZN(n3874) );
  INV_X4 U5031 ( .A(n3874), .ZN(n6123) );
  NAND2_X2 U5032 ( .A1(n6123), .A2(n2788), .ZN(n3838) );
  OAI221_X2 U5033 ( .B1(n6409), .B2(n3903), .C1(n2629), .C2(n3193), .A(n3838), 
        .ZN(n2086) );
  NAND2_X2 U5034 ( .A1(n3193), .A2(n2885), .ZN(n3875) );
  INV_X4 U5035 ( .A(n3875), .ZN(n6122) );
  NAND2_X2 U5036 ( .A1(n6122), .A2(n2788), .ZN(n3839) );
  NAND2_X2 U5037 ( .A1(n3197), .A2(n2713), .ZN(n3841) );
  NAND2_X2 U5038 ( .A1(n6131), .A2(n2883), .ZN(n3840) );
  NAND2_X2 U5039 ( .A1(n3198), .A2(n2864), .ZN(n3843) );
  NAND2_X2 U5040 ( .A1(n6131), .A2(n2884), .ZN(n3842) );
  NAND2_X2 U5041 ( .A1(n3197), .A2(n2858), .ZN(n3845) );
  NAND2_X2 U5042 ( .A1(n6131), .A2(n2885), .ZN(n3844) );
  NAND2_X2 U5043 ( .A1(n3197), .A2(n2869), .ZN(n3847) );
  NAND2_X2 U5044 ( .A1(n6131), .A2(n2886), .ZN(n3846) );
  NAND2_X2 U5045 ( .A1(n3197), .A2(n2859), .ZN(n3848) );
  AOI22_X2 U5046 ( .A1(n6121), .A2(n6400), .B1(n6131), .B2(n2955), .ZN(n3850)
         );
  NAND2_X2 U5047 ( .A1(n3851), .A2(n3850), .ZN(n2095) );
  AOI22_X2 U5048 ( .A1(n6400), .A2(n6127), .B1(n6131), .B2(n2956), .ZN(n3852)
         );
  NAND2_X2 U5049 ( .A1(n3853), .A2(n3852), .ZN(n2096) );
  AOI22_X2 U5050 ( .A1(n6120), .A2(n6400), .B1(n6131), .B2(n2957), .ZN(n3854)
         );
  NAND2_X2 U5051 ( .A1(n3855), .A2(n3854), .ZN(n2097) );
  AOI22_X2 U5052 ( .A1(n6119), .A2(n6400), .B1(n6131), .B2(n2958), .ZN(n3856)
         );
  NAND2_X2 U5053 ( .A1(n3857), .A2(n3856), .ZN(n2098) );
  AOI22_X2 U5054 ( .A1(n6129), .A2(n6369), .B1(n6118), .B2(n6400), .ZN(n3858)
         );
  NAND2_X2 U5055 ( .A1(n3859), .A2(n3858), .ZN(n2099) );
  AOI22_X2 U5056 ( .A1(n2960), .A2(n6400), .B1(n6131), .B2(n2712), .ZN(n3860)
         );
  NAND2_X2 U5057 ( .A1(n3861), .A2(n3860), .ZN(n2100) );
  AOI22_X2 U5058 ( .A1(n2764), .A2(n6400), .B1(n6131), .B2(n2649), .ZN(n3862)
         );
  NAND2_X2 U5059 ( .A1(n3863), .A2(n3862), .ZN(n2101) );
  AOI22_X2 U5060 ( .A1(n2763), .A2(n6400), .B1(n6131), .B2(n2871), .ZN(n3864)
         );
  NAND2_X2 U5061 ( .A1(n3865), .A2(n3864), .ZN(n2102) );
  AOI22_X2 U5062 ( .A1(n2762), .A2(n6400), .B1(n6131), .B2(n2636), .ZN(n3866)
         );
  NAND2_X2 U5063 ( .A1(n3867), .A2(n3866), .ZN(n2103) );
  NAND2_X2 U5064 ( .A1(n6400), .A2(n2981), .ZN(n3871) );
  NAND2_X2 U5065 ( .A1(n3197), .A2(n2861), .ZN(n3870) );
  NAND2_X2 U5066 ( .A1(n6131), .A2(n2837), .ZN(n3869) );
  INV_X4 U5067 ( .A(n6401), .ZN(n3868) );
  NAND4_X2 U5068 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n2104)
         );
  NAND2_X2 U5069 ( .A1(n6134), .A2(n6399), .ZN(n3872) );
  OAI22_X2 U5070 ( .A1(n6608), .A2(n3193), .B1(n6369), .B2(n3873), .ZN(n2106)
         );
  OAI22_X2 U5071 ( .A1(n6604), .A2(n3193), .B1(n6369), .B2(n3874), .ZN(n2107)
         );
  OAI22_X2 U5072 ( .A1(n6607), .A2(n3193), .B1(n6369), .B2(n3875), .ZN(n2108)
         );
  NAND2_X2 U5073 ( .A1(n3194), .A2(n2886), .ZN(n3901) );
  OAI22_X2 U5074 ( .A1(n6606), .A2(n3193), .B1(n6369), .B2(n3901), .ZN(n2109)
         );
  NAND2_X2 U5075 ( .A1(n6116), .A2(n6399), .ZN(n3876) );
  NAND2_X2 U5076 ( .A1(n6115), .A2(n6399), .ZN(n3877) );
  NAND2_X2 U5077 ( .A1(n6114), .A2(n6399), .ZN(n3878) );
  NAND2_X2 U5078 ( .A1(n3197), .A2(n2839), .ZN(n3880) );
  NAND2_X2 U5079 ( .A1(n6113), .A2(n6399), .ZN(n3879) );
  NAND2_X2 U5080 ( .A1(n3880), .A2(n3879), .ZN(n6767) );
  NAND2_X2 U5081 ( .A1(n6112), .A2(n6399), .ZN(n3881) );
  NAND2_X2 U5082 ( .A1(n6129), .A2(n6399), .ZN(n3882) );
  NAND2_X2 U5083 ( .A1(n3889), .A2(n2712), .ZN(n3884) );
  NAND2_X2 U5084 ( .A1(n3197), .A2(n2838), .ZN(n3883) );
  NAND2_X2 U5085 ( .A1(n3884), .A2(n3883), .ZN(n2116) );
  NAND2_X2 U5086 ( .A1(n6126), .A2(n6399), .ZN(n3885) );
  NAND2_X2 U5087 ( .A1(n3889), .A2(n2871), .ZN(n3887) );
  NAND2_X2 U5088 ( .A1(n3198), .A2(n2833), .ZN(n3886) );
  NAND2_X2 U5089 ( .A1(n3887), .A2(n3886), .ZN(n2118) );
  NAND2_X2 U5090 ( .A1(n6125), .A2(n6399), .ZN(n3888) );
  NAND2_X2 U5091 ( .A1(n3889), .A2(n2837), .ZN(n3890) );
  NAND2_X2 U5092 ( .A1(n3198), .A2(n2757), .ZN(n3891) );
  OAI221_X2 U5093 ( .B1(n6589), .B2(n6371), .C1(n2603), .C2(n6398), .A(n3891), 
        .ZN(n2123) );
  NAND2_X2 U5094 ( .A1(n3198), .A2(n2758), .ZN(n3892) );
  OAI221_X2 U5095 ( .B1(n2630), .B2(n6371), .C1(n6397), .C2(n6398), .A(n3892), 
        .ZN(n2126) );
  NAND2_X2 U5096 ( .A1(n3194), .A2(op0_1), .ZN(n5170) );
  NAND2_X2 U5097 ( .A1(op0_2), .A2(n3198), .ZN(n3893) );
  NAND2_X2 U5098 ( .A1(n5170), .A2(n3893), .ZN(n2127) );
  NAND2_X2 U5099 ( .A1(n2712), .A2(n6386), .ZN(n3895) );
  NAND2_X2 U5100 ( .A1(n3198), .A2(n2872), .ZN(n3894) );
  MUX2_X2 U5101 ( .A(n2798), .B(n6396), .S(n3190), .Z(n2130) );
  MUX2_X2 U5102 ( .A(n2737), .B(n6400), .S(n3190), .Z(n2131) );
  INV_X4 U5103 ( .A(n6137), .ZN(n3896) );
  OAI22_X2 U5104 ( .A1(n6597), .A2(n3193), .B1(n6370), .B2(n3896), .ZN(n6771)
         );
  INV_X4 U5105 ( .A(n6128), .ZN(n3897) );
  OAI22_X2 U5106 ( .A1(n6526), .A2(n3193), .B1(n6394), .B2(n3897), .ZN(n2133)
         );
  NAND2_X2 U5107 ( .A1(n6442), .A2(n6590), .ZN(n5169) );
  MUX2_X2 U5108 ( .A(n3245), .B(n6384), .S(n3190), .Z(n2136) );
  INV_X4 U5109 ( .A(n6383), .ZN(n3899) );
  NAND2_X2 U5110 ( .A1(n3198), .A2(n2595), .ZN(n3898) );
  AND3_X2 U5111 ( .A1(n6382), .A2(n3899), .A3(n3898), .ZN(n3900) );
  OAI221_X2 U5112 ( .B1(n6433), .B2(n2603), .C1(n6418), .C2(n6316), .A(n3900), 
        .ZN(n2137) );
  INV_X4 U5113 ( .A(n3901), .ZN(n6117) );
  NAND2_X2 U5114 ( .A1(n6117), .A2(n2788), .ZN(n3902) );
  OAI221_X2 U5115 ( .B1(n6381), .B2(n3903), .C1(n2781), .C2(n3193), .A(n3902), 
        .ZN(n2138) );
  MUX2_X2 U5116 ( .A(instruction[1]), .B(n2636), .S(n3164), .Z(n2140) );
  MUX2_X2 U5117 ( .A(instruction[3]), .B(n2649), .S(n3164), .Z(n2142) );
  MUX2_X2 U5118 ( .A(instruction[5]), .B(n2604), .S(n3164), .Z(n2144) );
  MUX2_X2 U5119 ( .A(instruction[6]), .B(n2958), .S(n3164), .Z(n2145) );
  MUX2_X2 U5120 ( .A(instruction[7]), .B(n2957), .S(n3164), .Z(n2146) );
  MUX2_X2 U5121 ( .A(instruction[8]), .B(n2956), .S(n3164), .Z(n2147) );
  MUX2_X2 U5122 ( .A(instruction[9]), .B(n2955), .S(n3164), .Z(n2148) );
  MUX2_X2 U5123 ( .A(instruction[10]), .B(n2678), .S(n3164), .Z(n2149) );
  MUX2_X2 U5124 ( .A(instruction[11]), .B(n2886), .S(n3164), .Z(n2150) );
  MUX2_X2 U5125 ( .A(instruction[12]), .B(n2885), .S(n3164), .Z(n2151) );
  MUX2_X2 U5126 ( .A(instruction[13]), .B(n2884), .S(n3164), .Z(n2152) );
  MUX2_X2 U5127 ( .A(instruction[14]), .B(n2883), .S(n3164), .Z(n2153) );
  MUX2_X2 U5128 ( .A(instruction[15]), .B(n2679), .S(n3164), .Z(n2154) );
  MUX2_X2 U5129 ( .A(instruction[16]), .B(n2975), .S(n3164), .Z(n2155) );
  MUX2_X2 U5130 ( .A(instruction[17]), .B(n2974), .S(n3164), .Z(n2156) );
  MUX2_X2 U5131 ( .A(instruction[18]), .B(n2973), .S(n3164), .Z(n2157) );
  MUX2_X2 U5132 ( .A(instruction[19]), .B(n2972), .S(n3164), .Z(n2158) );
  MUX2_X2 U5133 ( .A(instruction[20]), .B(n2661), .S(n3164), .Z(n2159) );
  MUX2_X2 U5134 ( .A(instruction[21]), .B(rs1[0]), .S(n3165), .Z(n2160) );
  MUX2_X2 U5135 ( .A(instruction[22]), .B(rs1[1]), .S(n3165), .Z(n2161) );
  MUX2_X2 U5136 ( .A(instruction[23]), .B(rs1[2]), .S(n3165), .Z(n2162) );
  MUX2_X2 U5137 ( .A(instruction[24]), .B(rs1[3]), .S(n3165), .Z(n2163) );
  MUX2_X2 U5138 ( .A(instruction[25]), .B(rs1[4]), .S(n3165), .Z(n2164) );
  MUX2_X2 U5139 ( .A(instruction[26]), .B(op0_1), .S(n3165), .Z(n2165) );
  MUX2_X2 U5140 ( .A(instruction[27]), .B(n2594), .S(n3165), .Z(n2166) );
  MUX2_X2 U5141 ( .A(instruction[28]), .B(n2597), .S(n3165), .Z(n2167) );
  MUX2_X2 U5142 ( .A(instruction[29]), .B(n2780), .S(n3165), .Z(n2168) );
  MUX2_X2 U5143 ( .A(instruction[30]), .B(n2650), .S(n3165), .Z(n2169) );
  MUX2_X2 U5144 ( .A(instruction[31]), .B(n2662), .S(n3165), .Z(n2170) );
  MUX2_X2 U5145 ( .A(n2738), .B(n2931), .S(n3190), .Z(n2175) );
  MUX2_X2 U5146 ( .A(n3904), .B(n2931), .S(n3166), .Z(n2176) );
  MUX2_X2 U5147 ( .A(n2739), .B(n2932), .S(n3189), .Z(n2177) );
  MUX2_X2 U5148 ( .A(n3905), .B(n2932), .S(n3166), .Z(n2178) );
  MUX2_X2 U5149 ( .A(n2740), .B(n2933), .S(n3189), .Z(n2179) );
  MUX2_X2 U5150 ( .A(n3906), .B(n2933), .S(n3166), .Z(n2180) );
  MUX2_X2 U5151 ( .A(n2741), .B(n2934), .S(n3189), .Z(n2181) );
  MUX2_X2 U5152 ( .A(n3907), .B(n2934), .S(n3166), .Z(n2182) );
  MUX2_X2 U5153 ( .A(n2742), .B(n2935), .S(n3189), .Z(n2183) );
  MUX2_X2 U5154 ( .A(n3908), .B(n2935), .S(n3166), .Z(n2184) );
  MUX2_X2 U5155 ( .A(n2743), .B(n2936), .S(n3189), .Z(n2185) );
  MUX2_X2 U5156 ( .A(n3909), .B(n2936), .S(n3166), .Z(n2186) );
  MUX2_X2 U5157 ( .A(n2744), .B(n2937), .S(n3189), .Z(n2187) );
  MUX2_X2 U5158 ( .A(n2760), .B(n2937), .S(n3166), .Z(n2188) );
  MUX2_X2 U5159 ( .A(n2745), .B(n2938), .S(n3189), .Z(n2189) );
  MUX2_X2 U5160 ( .A(n3910), .B(n2938), .S(n3166), .Z(n2190) );
  MUX2_X2 U5161 ( .A(n2746), .B(n2939), .S(n3191), .Z(n2191) );
  MUX2_X2 U5162 ( .A(n3911), .B(n2939), .S(n3166), .Z(n2192) );
  MUX2_X2 U5163 ( .A(n2747), .B(n2940), .S(n3189), .Z(n2193) );
  MUX2_X2 U5164 ( .A(n3912), .B(n2940), .S(n3166), .Z(n2194) );
  MUX2_X2 U5165 ( .A(n2899), .B(n2759), .S(n3189), .Z(n2195) );
  MUX2_X2 U5166 ( .A(n2984), .B(n2759), .S(n3166), .Z(n2196) );
  MUX2_X2 U5167 ( .A(n2748), .B(n2941), .S(n3189), .Z(n2197) );
  MUX2_X2 U5168 ( .A(n3913), .B(n2941), .S(n3166), .Z(n2198) );
  MUX2_X2 U5169 ( .A(n2749), .B(n2942), .S(n3189), .Z(n2199) );
  MUX2_X2 U5170 ( .A(n3914), .B(n2942), .S(n3165), .Z(n2200) );
  MUX2_X2 U5171 ( .A(n2750), .B(n2943), .S(n3189), .Z(n2201) );
  MUX2_X2 U5172 ( .A(n3915), .B(n2943), .S(n3166), .Z(n2202) );
  MUX2_X2 U5173 ( .A(n2751), .B(n2944), .S(n3189), .Z(n2203) );
  MUX2_X2 U5174 ( .A(n3916), .B(n2944), .S(n3165), .Z(n2204) );
  MUX2_X2 U5175 ( .A(n2752), .B(n2945), .S(n3189), .Z(n2205) );
  MUX2_X2 U5176 ( .A(n3917), .B(n2945), .S(n3166), .Z(n2206) );
  MUX2_X2 U5177 ( .A(n2753), .B(n2946), .S(n3189), .Z(n2207) );
  MUX2_X2 U5178 ( .A(n3918), .B(n2946), .S(n3165), .Z(n2208) );
  MUX2_X2 U5179 ( .A(n2754), .B(n2947), .S(n3189), .Z(n2209) );
  MUX2_X2 U5180 ( .A(n3919), .B(n2947), .S(n3166), .Z(n2210) );
  MUX2_X2 U5181 ( .A(n2755), .B(n2948), .S(n3188), .Z(n2211) );
  MUX2_X2 U5182 ( .A(n3920), .B(n2948), .S(n3165), .Z(n2212) );
  MUX2_X2 U5183 ( .A(n2756), .B(n2949), .S(n3188), .Z(n2213) );
  MUX2_X2 U5184 ( .A(n3922), .B(n2949), .S(n3166), .Z(n2214) );
  NAND4_X2 U5185 ( .A1(n3055), .A2(n6313), .A3(n3064), .A4(n3235), .ZN(n4073)
         );
  NAND2_X2 U5186 ( .A1(n3924), .A2(n3923), .ZN(n4250) );
  NAND2_X2 U5187 ( .A1(n4524), .A2(memAddr[7]), .ZN(n4252) );
  INV_X4 U5188 ( .A(n4252), .ZN(n4254) );
  INV_X4 U5189 ( .A(n4251), .ZN(n4253) );
  NAND2_X2 U5190 ( .A1(n3927), .A2(n3177), .ZN(n3933) );
  NAND3_X2 U5191 ( .A1(n3928), .A2(n3170), .A3(n3178), .ZN(n3932) );
  NAND2_X2 U5192 ( .A1(reg31Val_0[16]), .A2(n3233), .ZN(n4147) );
  NAND3_X2 U5193 ( .A1(n3933), .A2(n3932), .A3(n3931), .ZN(n4312) );
  INV_X4 U5194 ( .A(n4312), .ZN(n3934) );
  NOR3_X4 U5195 ( .A1(n4390), .A2(n6338), .A3(n3173), .ZN(n3937) );
  NOR3_X4 U5196 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n3940) );
  NAND3_X4 U5197 ( .A1(n3170), .A2(\wb/dsize_reg/z2 [21]), .A3(n4114), .ZN(
        n3939) );
  NAND2_X2 U5198 ( .A1(n3178), .A2(n3233), .ZN(n4391) );
  NAND3_X4 U5199 ( .A1(reg31Val_0[21]), .A2(n3170), .A3(n3969), .ZN(n3938) );
  NAND3_X4 U5200 ( .A1(n3939), .A2(n3940), .A3(n3938), .ZN(n4376) );
  INV_X4 U5201 ( .A(n4376), .ZN(n3941) );
  INV_X4 U5202 ( .A(n4391), .ZN(n3945) );
  INV_X4 U5203 ( .A(n4230), .ZN(n3949) );
  NAND2_X2 U5204 ( .A1(n3950), .A2(n3177), .ZN(n3956) );
  NAND3_X2 U5205 ( .A1(n3951), .A2(n4355), .A3(n3178), .ZN(n3955) );
  NAND3_X2 U5206 ( .A1(n3952), .A2(n3075), .A3(n3178), .ZN(n3954) );
  NAND4_X2 U5207 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n4374)
         );
  INV_X4 U5208 ( .A(n4374), .ZN(n3957) );
  NAND2_X2 U5209 ( .A1(n3958), .A2(n3105), .ZN(n3964) );
  NAND3_X2 U5210 ( .A1(n3959), .A2(n4355), .A3(n3178), .ZN(n3963) );
  NAND3_X2 U5211 ( .A1(n3960), .A2(n3170), .A3(n3178), .ZN(n3962) );
  NAND4_X2 U5212 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n4412)
         );
  INV_X4 U5213 ( .A(n4412), .ZN(n3965) );
  INV_X4 U5214 ( .A(n4391), .ZN(n3969) );
  INV_X4 U5215 ( .A(n4373), .ZN(n3973) );
  INV_X4 U5216 ( .A(n4300), .ZN(n3974) );
  NAND2_X2 U5217 ( .A1(n3974), .A2(n3177), .ZN(n3977) );
  NAND2_X2 U5218 ( .A1(n2887), .A2(n3177), .ZN(n3976) );
  NAND2_X2 U5219 ( .A1(n2891), .A2(n3177), .ZN(n3975) );
  NAND2_X2 U5220 ( .A1(n4524), .A2(memAddr[31]), .ZN(n4303) );
  NAND2_X2 U5221 ( .A1(n4303), .A2(n4304), .ZN(n4302) );
  INV_X4 U5222 ( .A(n4214), .ZN(n4206) );
  NAND2_X2 U5223 ( .A1(n3980), .A2(n3177), .ZN(n4215) );
  AND2_X2 U5224 ( .A1(n4219), .A2(n4213), .ZN(n3981) );
  NAND2_X2 U5225 ( .A1(n4524), .A2(memAddr[4]), .ZN(n4218) );
  INV_X4 U5226 ( .A(n4218), .ZN(n4208) );
  INV_X4 U5227 ( .A(n4220), .ZN(n4209) );
  NAND2_X2 U5228 ( .A1(n3985), .A2(n3167), .ZN(n4275) );
  INV_X4 U5229 ( .A(n4275), .ZN(n3988) );
  INV_X4 U5230 ( .A(n4278), .ZN(n3987) );
  NAND3_X4 U5231 ( .A1(n3989), .A2(n4355), .A3(n3176), .ZN(n4274) );
  INV_X4 U5232 ( .A(n4274), .ZN(n3992) );
  NAND2_X2 U5233 ( .A1(n4626), .A2(n4628), .ZN(n4635) );
  NAND3_X4 U5234 ( .A1(\wb/dsize_reg/z2 [2]), .A2(n4010), .A3(n3176), .ZN(
        n4624) );
  NAND2_X2 U5235 ( .A1(n3996), .A2(n3177), .ZN(n4491) );
  NAND2_X2 U5236 ( .A1(n4491), .A2(n4492), .ZN(n3997) );
  INV_X4 U5237 ( .A(n3997), .ZN(n4623) );
  INV_X4 U5238 ( .A(n4614), .ZN(n4003) );
  INV_X4 U5239 ( .A(n4002), .ZN(n4619) );
  NAND4_X2 U5240 ( .A1(n4611), .A2(n4003), .A3(n4612), .A4(n4619), .ZN(
        regWrData[1]) );
  INV_X4 U5241 ( .A(n4175), .ZN(n4004) );
  NAND2_X2 U5242 ( .A1(n4524), .A2(memAddr[1]), .ZN(n4176) );
  NAND2_X2 U5243 ( .A1(n4524), .A2(memAddr[3]), .ZN(n4198) );
  INV_X4 U5244 ( .A(n4198), .ZN(n4188) );
  INV_X4 U5245 ( .A(n4199), .ZN(n4192) );
  NAND2_X2 U5246 ( .A1(n4009), .A2(n3167), .ZN(n4382) );
  INV_X4 U5247 ( .A(n3145), .ZN(n4010) );
  NAND2_X2 U5248 ( .A1(n4440), .A2(n3167), .ZN(n4528) );
  NAND4_X2 U5249 ( .A1(n4382), .A2(n4380), .A3(n4381), .A4(n4386), .ZN(
        regWrData[6]) );
  INV_X4 U5250 ( .A(n4378), .ZN(n4013) );
  NAND2_X2 U5251 ( .A1(n4524), .A2(memAddr[6]), .ZN(n4379) );
  INV_X4 U5252 ( .A(n4360), .ZN(n4016) );
  AOI211_X2 U5253 ( .C1(n3075), .C2(regWrData[11]), .A(n3070), .B(n4016), .ZN(
        n4017) );
  INV_X4 U5254 ( .A(n4375), .ZN(n4024) );
  NAND2_X2 U5255 ( .A1(n4357), .A2(n3025), .ZN(n4295) );
  INV_X4 U5256 ( .A(n4295), .ZN(n4025) );
  NAND2_X2 U5257 ( .A1(n4025), .A2(n3177), .ZN(n4033) );
  NAND2_X2 U5258 ( .A1(reg31Val_0[8]), .A2(n3233), .ZN(n4293) );
  INV_X4 U5259 ( .A(n4293), .ZN(n4026) );
  NAND2_X2 U5260 ( .A1(n4026), .A2(n3105), .ZN(n4032) );
  NAND4_X2 U5261 ( .A1(\wb/dsize_reg/z2 [24]), .A2(n3055), .A3(n4029), .A4(
        n4028), .ZN(n4030) );
  NAND2_X2 U5262 ( .A1(n4035), .A2(n3177), .ZN(n4511) );
  INV_X4 U5263 ( .A(n4316), .ZN(n4036) );
  NAND2_X2 U5264 ( .A1(n4139), .A2(n3026), .ZN(n4320) );
  INV_X4 U5265 ( .A(n4313), .ZN(n4037) );
  NAND2_X2 U5266 ( .A1(n4524), .A2(memAddr[12]), .ZN(n4314) );
  NAND2_X2 U5267 ( .A1(n4039), .A2(n3167), .ZN(n4339) );
  INV_X4 U5268 ( .A(n4340), .ZN(n4043) );
  NAND2_X2 U5269 ( .A1(n4524), .A2(memAddr[13]), .ZN(n4341) );
  NAND3_X2 U5270 ( .A1(n4355), .A2(n3178), .A3(\wb/dsize_reg/z2 [10]), .ZN(
        n4048) );
  NAND3_X2 U5271 ( .A1(n3178), .A2(n3233), .A3(reg31Val_0[10]), .ZN(n4047) );
  NAND3_X2 U5272 ( .A1(n3178), .A2(n2989), .A3(n4357), .ZN(n4046) );
  NAND4_X2 U5273 ( .A1(n4048), .A2(n4264), .A3(n4047), .A4(n4046), .ZN(
        regWrData[10]) );
  INV_X4 U5274 ( .A(n4263), .ZN(n4049) );
  AOI211_X2 U5275 ( .C1(n3075), .C2(regWrData[10]), .A(n4050), .B(n4049), .ZN(
        n4051) );
  NAND2_X2 U5276 ( .A1(n4052), .A2(n3177), .ZN(n4059) );
  NAND3_X2 U5277 ( .A1(n4053), .A2(n3075), .A3(n3178), .ZN(n4058) );
  NAND2_X2 U5278 ( .A1(reg31Val_0[30]), .A2(n3233), .ZN(n4054) );
  INV_X4 U5279 ( .A(n4246), .ZN(n4060) );
  NAND4_X2 U5280 ( .A1(n3177), .A2(n2991), .A3(n4357), .A4(n3075), .ZN(n4064)
         );
  NAND4_X2 U5281 ( .A1(\wb/dsize_reg/z2 [19]), .A2(n3178), .A3(n4355), .A4(
        n3075), .ZN(n4063) );
  NAND4_X2 U5282 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4372)
         );
  INV_X4 U5283 ( .A(n4372), .ZN(n4067) );
  INV_X4 U5284 ( .A(n6254), .ZN(n4068) );
  NAND2_X2 U5285 ( .A1(n6231), .A2(n4068), .ZN(n4069) );
  NAND2_X2 U5286 ( .A1(n3183), .A2(memAddr[19]), .ZN(n4070) );
  NAND2_X2 U5287 ( .A1(n4074), .A2(n3168), .ZN(n4406) );
  NAND3_X4 U5288 ( .A1(\wb/dsize_reg/z2 [5]), .A2(n4010), .A3(n3168), .ZN(
        n4401) );
  NAND2_X2 U5289 ( .A1(n4081), .A2(n4080), .ZN(regWrData[14]) );
  INV_X4 U5290 ( .A(n4328), .ZN(n4082) );
  INV_X4 U5291 ( .A(n4235), .ZN(n4089) );
  NAND2_X2 U5292 ( .A1(n4139), .A2(n3027), .ZN(n4238) );
  NAND2_X2 U5293 ( .A1(n4085), .A2(n3177), .ZN(n4231) );
  INV_X4 U5294 ( .A(n4231), .ZN(n4087) );
  NAND2_X2 U5295 ( .A1(n4092), .A2(n3177), .ZN(n4097) );
  NAND2_X2 U5296 ( .A1(n4093), .A2(n3177), .ZN(n4096) );
  NAND2_X2 U5297 ( .A1(n4094), .A2(n3177), .ZN(n4095) );
  NAND3_X4 U5298 ( .A1(n4097), .A2(n4096), .A3(n4095), .ZN(regWrData[17]) );
  NAND2_X2 U5299 ( .A1(n4100), .A2(n4099), .ZN(n4395) );
  NAND4_X2 U5300 ( .A1(n4102), .A2(n3234), .A3(n3174), .A4(n3177), .ZN(n4108)
         );
  NAND4_X2 U5301 ( .A1(n4105), .A2(\wb/dsize_reg/z2 [18]), .A3(n3174), .A4(
        n3177), .ZN(n4106) );
  NAND4_X2 U5302 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4272)
         );
  INV_X4 U5303 ( .A(n4272), .ZN(n4110) );
  INV_X4 U5304 ( .A(n4413), .ZN(n4118) );
  NAND4_X2 U5305 ( .A1(n3177), .A2(n3233), .A3(reg31Val_0[26]), .A4(n3170), 
        .ZN(n4123) );
  NAND3_X2 U5306 ( .A1(n4357), .A2(n3178), .A3(n4120), .ZN(n4121) );
  NAND4_X2 U5307 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4229)
         );
  NAND3_X2 U5308 ( .A1(n4126), .A2(n4355), .A3(n3178), .ZN(n4133) );
  NAND2_X2 U5309 ( .A1(n4127), .A2(n3105), .ZN(n4132) );
  NAND3_X2 U5310 ( .A1(n4128), .A2(n3170), .A3(n3178), .ZN(n4131) );
  NAND4_X2 U5311 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4414)
         );
  INV_X4 U5312 ( .A(n4414), .ZN(n4134) );
  NAND4_X2 U5313 ( .A1(n3233), .A2(n3170), .A3(reg31Val_0[28]), .A4(n3177), 
        .ZN(n4141) );
  INV_X4 U5314 ( .A(n4228), .ZN(n4144) );
  INV_X4 U5315 ( .A(regWrData[17]), .ZN(n4146) );
  NAND2_X2 U5316 ( .A1(n3182), .A2(memAddr[17]), .ZN(n4145) );
  INV_X4 U5317 ( .A(n4147), .ZN(n4148) );
  NAND2_X2 U5318 ( .A1(n4148), .A2(n3177), .ZN(n4151) );
  NAND4_X2 U5319 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(
        regWrData[9]) );
  NAND3_X2 U5320 ( .A1(n3178), .A2(n2995), .A3(n4357), .ZN(n4160) );
  NAND3_X2 U5321 ( .A1(\wb/dsize_reg/z2 [30]), .A2(n3178), .A3(n4355), .ZN(
        n4159) );
  OAI211_X2 U5322 ( .C1(n3154), .C2(n2980), .A(n4160), .B(n4159), .ZN(
        regWrData[30]) );
  OAI222_X2 U5323 ( .A1(n6337), .A2(n4162), .B1(n2687), .B2(n3152), .C1(n3154), 
        .C2(n2928), .ZN(regWrData[22]) );
  NAND3_X2 U5324 ( .A1(n4491), .A2(n4628), .A3(n4626), .ZN(n4169) );
  NAND4_X2 U5325 ( .A1(n3243), .A2(n4624), .A3(n4165), .A4(n4492), .ZN(n4168)
         );
  NAND2_X2 U5326 ( .A1(n6601), .A2(n3245), .ZN(n4167) );
  NAND3_X4 U5327 ( .A1(n4173), .A2(n4172), .A3(n2790), .ZN(n4174) );
  NAND2_X2 U5328 ( .A1(n4174), .A2(n3177), .ZN(n4179) );
  NAND2_X2 U5329 ( .A1(n4176), .A2(n4175), .ZN(n4180) );
  NAND2_X2 U5330 ( .A1(n3243), .A2(n4180), .ZN(n4178) );
  NAND3_X2 U5331 ( .A1(n4179), .A2(n4178), .A3(n4177), .ZN(n4182) );
  INV_X4 U5332 ( .A(n4180), .ZN(n4181) );
  NAND2_X2 U5333 ( .A1(n4181), .A2(n3173), .ZN(n4184) );
  NAND2_X2 U5334 ( .A1(n4182), .A2(n4184), .ZN(n4187) );
  NAND2_X2 U5335 ( .A1(n4185), .A2(n4184), .ZN(n4186) );
  NAND3_X4 U5336 ( .A1(n4187), .A2(n2877), .A3(n4186), .ZN(n6040) );
  NAND2_X2 U5337 ( .A1(n6635), .A2(n3097), .ZN(n4202) );
  NAND4_X2 U5338 ( .A1(n3243), .A2(n4199), .A3(n4198), .A4(n3172), .ZN(n4200)
         );
  NAND2_X2 U5339 ( .A1(n4219), .A2(n4215), .ZN(n4207) );
  NAND4_X2 U5340 ( .A1(n4212), .A2(n4213), .A3(n4211), .A4(n4210), .ZN(n4225)
         );
  INV_X4 U5341 ( .A(n4213), .ZN(n4217) );
  NAND2_X2 U5342 ( .A1(n4223), .A2(n4222), .ZN(n4224) );
  MUX2_X2 U5343 ( .A(n2858), .B(n4228), .S(n3243), .Z(n5111) );
  MUX2_X2 U5344 ( .A(n2859), .B(n4229), .S(n3243), .Z(n5003) );
  INV_X4 U5345 ( .A(n5003), .ZN(n4995) );
  NAND3_X2 U5346 ( .A1(n4233), .A2(n4232), .A3(n3172), .ZN(n4240) );
  NAND2_X2 U5347 ( .A1(n4234), .A2(n4240), .ZN(n4237) );
  NAND2_X2 U5348 ( .A1(n4235), .A2(n4240), .ZN(n4236) );
  NAND2_X2 U5349 ( .A1(n4237), .A2(n4236), .ZN(n4245) );
  NAND4_X2 U5350 ( .A1(n4355), .A2(n3178), .A3(\wb/dsize_reg/z2 [15]), .A4(
        n4240), .ZN(n4242) );
  INV_X4 U5351 ( .A(n4238), .ZN(n4239) );
  NAND2_X2 U5352 ( .A1(n4240), .A2(n4239), .ZN(n4241) );
  NAND2_X2 U5353 ( .A1(n6609), .A2(n3245), .ZN(n4243) );
  MUX2_X2 U5354 ( .A(n2713), .B(n4246), .S(n3243), .Z(n5720) );
  NAND2_X2 U5355 ( .A1(reg31Val_0[10]), .A2(n3233), .ZN(n4261) );
  INV_X4 U5356 ( .A(n4264), .ZN(n4265) );
  INV_X4 U5357 ( .A(n4268), .ZN(n4270) );
  NAND2_X2 U5358 ( .A1(n6629), .A2(n3245), .ZN(n4269) );
  NAND3_X4 U5359 ( .A1(n4270), .A2(n4271), .A3(n4269), .ZN(n5346) );
  MUX2_X2 U5360 ( .A(n2860), .B(n4272), .S(n3243), .Z(n4773) );
  NAND2_X2 U5361 ( .A1(n6630), .A2(n3097), .ZN(n4280) );
  OAI21_X4 U5362 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(n5633) );
  NAND2_X2 U5363 ( .A1(n4283), .A2(n3173), .ZN(n4287) );
  INV_X4 U5364 ( .A(n4284), .ZN(n4285) );
  NAND2_X2 U5365 ( .A1(n6631), .A2(n3097), .ZN(n4286) );
  OAI21_X4 U5366 ( .B1(n4287), .B2(n2993), .A(n4286), .ZN(n4288) );
  NAND4_X2 U5367 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), .ZN(n4297)
         );
  NAND3_X2 U5368 ( .A1(n4301), .A2(n4300), .A3(n4299), .ZN(n4311) );
  NAND2_X2 U5369 ( .A1(n6605), .A2(n3245), .ZN(n4310) );
  NAND2_X2 U5370 ( .A1(n4303), .A2(n3173), .ZN(n4306) );
  INV_X4 U5371 ( .A(n4304), .ZN(n4305) );
  MUX2_X2 U5372 ( .A(n2861), .B(n4312), .S(n3243), .Z(n5949) );
  INV_X4 U5373 ( .A(n5949), .ZN(n4675) );
  NAND3_X2 U5374 ( .A1(n4313), .A2(n4511), .A3(n4314), .ZN(n4315) );
  NAND3_X2 U5375 ( .A1(n4314), .A2(n4313), .A3(n3173), .ZN(n4321) );
  NAND2_X2 U5376 ( .A1(n4315), .A2(n4321), .ZN(n4318) );
  NAND2_X2 U5377 ( .A1(n4316), .A2(n4321), .ZN(n4317) );
  NAND2_X2 U5378 ( .A1(n4318), .A2(n4317), .ZN(n4327) );
  INV_X4 U5379 ( .A(n4320), .ZN(n4322) );
  NAND2_X2 U5380 ( .A1(n6607), .A2(n3245), .ZN(n4325) );
  OAI21_X4 U5381 ( .B1(n4326), .B2(n4327), .A(n4325), .ZN(n5392) );
  NAND4_X2 U5382 ( .A1(n4331), .A2(n3233), .A3(n3177), .A4(reg31Val_0[14]), 
        .ZN(n4336) );
  NAND4_X2 U5383 ( .A1(n4337), .A2(n4336), .A3(n4335), .A4(n4334), .ZN(n4338)
         );
  MUX2_X2 U5384 ( .A(n2854), .B(n4338), .S(n3243), .Z(n4883) );
  NAND3_X2 U5385 ( .A1(n4339), .A2(n4340), .A3(n3093), .ZN(n4342) );
  NAND3_X2 U5386 ( .A1(n4341), .A2(n4340), .A3(n3173), .ZN(n4348) );
  NAND2_X2 U5387 ( .A1(n4346), .A2(n4345), .ZN(n4353) );
  NAND3_X2 U5388 ( .A1(n4347), .A2(\wb/dsize_reg/z2 [13]), .A3(n4348), .ZN(
        n4350) );
  NAND2_X2 U5389 ( .A1(n6604), .A2(n3245), .ZN(n4351) );
  NAND3_X2 U5390 ( .A1(n4359), .A2(n4360), .A3(n3173), .ZN(n4361) );
  INV_X4 U5391 ( .A(n4358), .ZN(n4356) );
  NAND3_X4 U5392 ( .A1(n4357), .A2(n2811), .A3(n4356), .ZN(n4365) );
  NAND3_X4 U5393 ( .A1(reg31Val_0[11]), .A2(n3232), .A3(n4356), .ZN(n4364) );
  NAND4_X2 U5394 ( .A1(n4366), .A2(n4365), .A3(n4364), .A4(n4363), .ZN(n4367)
         );
  MUX2_X2 U5395 ( .A(n2855), .B(n4367), .S(n3243), .Z(n5543) );
  NAND4_X2 U5396 ( .A1(n4371), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(n4423)
         );
  MUX2_X2 U5397 ( .A(n2862), .B(n4372), .S(n3243), .Z(n5216) );
  MUX2_X2 U5398 ( .A(n2863), .B(n4373), .S(n3243), .Z(n5790) );
  MUX2_X2 U5399 ( .A(n2716), .B(n4374), .S(n3243), .Z(n5856) );
  INV_X4 U5400 ( .A(n5856), .ZN(n5860) );
  MUX2_X2 U5401 ( .A(n2864), .B(n4375), .S(n3243), .Z(n5463) );
  INV_X4 U5402 ( .A(n5463), .ZN(n5459) );
  MUX2_X2 U5403 ( .A(n2865), .B(n4376), .S(n3243), .Z(n5913) );
  INV_X4 U5404 ( .A(n5913), .ZN(n5019) );
  NAND2_X2 U5405 ( .A1(n5459), .A2(n5019), .ZN(n4431) );
  NAND2_X2 U5406 ( .A1(n4379), .A2(n4378), .ZN(n4384) );
  NAND3_X2 U5407 ( .A1(n4382), .A2(n4381), .A3(n4380), .ZN(n4383) );
  AOI21_X4 U5408 ( .B1(n4387), .B2(n4386), .A(n4385), .ZN(n4389) );
  NAND2_X2 U5409 ( .A1(n6633), .A2(n3245), .ZN(n4388) );
  OAI21_X4 U5410 ( .B1(n4389), .B2(n3245), .A(n4388), .ZN(n5554) );
  NAND2_X2 U5411 ( .A1(n4398), .A2(n4397), .ZN(n4399) );
  MUX2_X2 U5412 ( .A(n2866), .B(n4399), .S(n3243), .Z(n4679) );
  MUX2_X2 U5413 ( .A(n6634), .B(n4411), .S(n3243), .Z(n4916) );
  MUX2_X2 U5414 ( .A(n2867), .B(n4412), .S(n3243), .Z(n5816) );
  INV_X4 U5415 ( .A(n5816), .ZN(n4453) );
  MUX2_X2 U5416 ( .A(n2868), .B(n4413), .S(n3243), .Z(n4836) );
  MUX2_X2 U5417 ( .A(n2869), .B(n4414), .S(n3243), .Z(n5068) );
  NAND2_X2 U5418 ( .A1(n4418), .A2(n4417), .ZN(n4422) );
  NAND2_X2 U5419 ( .A1(n2680), .A2(regWrData[31]), .ZN(n4421) );
  NAND2_X2 U5420 ( .A1(n2723), .A2(n2639), .ZN(n4420) );
  NAND2_X2 U5421 ( .A1(n3182), .A2(memAddr[31]), .ZN(n4419) );
  NAND2_X2 U5422 ( .A1(n5185), .A2(n4445), .ZN(n5699) );
  INV_X4 U5423 ( .A(n5699), .ZN(n5718) );
  NAND2_X2 U5424 ( .A1(n5718), .A2(n2787), .ZN(n6016) );
  INV_X4 U5425 ( .A(n6016), .ZN(n5261) );
  OAI21_X4 U5426 ( .B1(n4423), .B2(n4422), .A(n5261), .ZN(n5688) );
  INV_X4 U5427 ( .A(n4431), .ZN(n4432) );
  NAND4_X2 U5428 ( .A1(n4433), .A2(n5860), .A3(n4880), .A4(n4432), .ZN(n4434)
         );
  INV_X4 U5429 ( .A(n4434), .ZN(n4460) );
  NAND2_X2 U5430 ( .A1(n2723), .A2(n2648), .ZN(n5151) );
  INV_X4 U5431 ( .A(n5146), .ZN(n4438) );
  NAND2_X2 U5432 ( .A1(n3182), .A2(memAddr[0]), .ZN(n5150) );
  INV_X4 U5433 ( .A(n5145), .ZN(n4444) );
  NAND3_X2 U5434 ( .A1(\wb/dsize_reg/z2 [24]), .A2(n3178), .A3(n4440), .ZN(
        n4441) );
  INV_X4 U5435 ( .A(n4443), .ZN(n5149) );
  INV_X4 U5436 ( .A(zeroExt_2), .ZN(n4445) );
  OAI211_X2 U5437 ( .C1(n4448), .C2(n4447), .A(n4446), .B(n4445), .ZN(n6010)
         );
  INV_X4 U5438 ( .A(n6010), .ZN(n6002) );
  NOR4_X2 U5439 ( .A1(n4449), .A2(n5492), .A3(n3061), .A4(n2602), .ZN(n4459)
         );
  NOR3_X4 U5440 ( .A1(n4452), .A2(n4451), .A3(n4450), .ZN(n4458) );
  NAND2_X2 U5441 ( .A1(n4454), .A2(n4453), .ZN(n4456) );
  NAND2_X2 U5442 ( .A1(n5081), .A2(n5718), .ZN(n4461) );
  NAND2_X2 U5443 ( .A1(n5661), .A2(n3157), .ZN(n4975) );
  INV_X4 U5444 ( .A(regWrData[23]), .ZN(n4464) );
  NAND2_X2 U5445 ( .A1(n3182), .A2(memAddr[23]), .ZN(n4463) );
  NAND2_X2 U5446 ( .A1(n5865), .A2(n3041), .ZN(n5701) );
  INV_X4 U5447 ( .A(n5701), .ZN(n5858) );
  NAND2_X2 U5448 ( .A1(n5081), .A2(n5858), .ZN(n4468) );
  NAND2_X2 U5449 ( .A1(n3182), .A2(memAddr[8]), .ZN(n4465) );
  NAND3_X2 U5450 ( .A1(n4468), .A2(n3217), .A3(n4467), .ZN(n4943) );
  NAND2_X2 U5451 ( .A1(n5082), .A2(n4943), .ZN(n4469) );
  NAND2_X2 U5452 ( .A1(n4470), .A2(n4469), .ZN(n5430) );
  INV_X4 U5453 ( .A(n6040), .ZN(n6037) );
  NAND2_X2 U5454 ( .A1(n3182), .A2(memAddr[14]), .ZN(n4877) );
  NAND2_X2 U5455 ( .A1(n2723), .A2(n2641), .ZN(n4878) );
  INV_X4 U5456 ( .A(n4471), .ZN(n4476) );
  INV_X4 U5457 ( .A(n4878), .ZN(n4472) );
  NAND4_X2 U5458 ( .A1(n4080), .A2(n4476), .A3(n4475), .A4(n4877), .ZN(n4477)
         );
  NAND2_X2 U5459 ( .A1(n5080), .A2(n4885), .ZN(n4480) );
  INV_X4 U5460 ( .A(n4735), .ZN(n4765) );
  NAND2_X2 U5461 ( .A1(n5081), .A2(n4765), .ZN(n4479) );
  INV_X4 U5462 ( .A(regWrData[6]), .ZN(n4482) );
  NAND2_X2 U5463 ( .A1(n3183), .A2(memAddr[6]), .ZN(n4481) );
  INV_X4 U5464 ( .A(n5555), .ZN(n5551) );
  NAND2_X2 U5465 ( .A1(n5080), .A2(n5551), .ZN(n4486) );
  INV_X4 U5466 ( .A(regWrData[25]), .ZN(n4484) );
  NAND2_X2 U5467 ( .A1(n3182), .A2(memAddr[25]), .ZN(n4483) );
  NAND2_X2 U5468 ( .A1(n5199), .A2(n4616), .ZN(n5785) );
  INV_X4 U5469 ( .A(n5785), .ZN(n5781) );
  NAND2_X2 U5470 ( .A1(n5081), .A2(n5781), .ZN(n4485) );
  NAND3_X4 U5471 ( .A1(n4486), .A2(n3216), .A3(n4485), .ZN(n4928) );
  NAND2_X2 U5472 ( .A1(n4981), .A2(n4928), .ZN(n4487) );
  NAND2_X2 U5473 ( .A1(n4488), .A2(n4487), .ZN(n4855) );
  AOI22_X2 U5474 ( .A1(n5514), .A2(n5430), .B1(n4867), .B2(n4855), .ZN(n4522)
         );
  INV_X4 U5475 ( .A(regWrData[29]), .ZN(n4490) );
  NAND2_X2 U5476 ( .A1(n3182), .A2(memAddr[29]), .ZN(n4489) );
  OAI221_X2 U5477 ( .B1(n6573), .B2(n3155), .C1(n4490), .C2(n3184), .A(n4489), 
        .ZN(n5187) );
  NAND2_X2 U5478 ( .A1(n5187), .A2(n4445), .ZN(n5462) );
  INV_X4 U5479 ( .A(n5462), .ZN(n5458) );
  NAND2_X2 U5480 ( .A1(n5081), .A2(n5458), .ZN(n4497) );
  NAND2_X2 U5481 ( .A1(n2723), .A2(n2646), .ZN(n5139) );
  NAND2_X2 U5482 ( .A1(n3182), .A2(memAddr[2]), .ZN(n5138) );
  NAND2_X2 U5483 ( .A1(n5139), .A2(n5138), .ZN(n4495) );
  NAND3_X4 U5484 ( .A1(n4491), .A2(n5138), .A3(n4624), .ZN(n4494) );
  NAND3_X4 U5485 ( .A1(n4492), .A2(n5139), .A3(n3998), .ZN(n4493) );
  NAND2_X2 U5486 ( .A1(n5080), .A2(n5611), .ZN(n4496) );
  INV_X4 U5487 ( .A(regWrData[21]), .ZN(n4499) );
  NAND2_X2 U5488 ( .A1(n3183), .A2(memAddr[21]), .ZN(n4498) );
  OAI221_X2 U5489 ( .B1(n6581), .B2(n3155), .C1(n4499), .C2(n3184), .A(n4498), 
        .ZN(n5930) );
  NAND2_X2 U5490 ( .A1(n5930), .A2(n4445), .ZN(n5908) );
  INV_X4 U5491 ( .A(n5908), .ZN(n5903) );
  NAND2_X2 U5492 ( .A1(n5081), .A2(n5903), .ZN(n4501) );
  NAND2_X2 U5493 ( .A1(n2723), .A2(n2645), .ZN(n4589) );
  NAND2_X2 U5494 ( .A1(n3183), .A2(memAddr[10]), .ZN(n4588) );
  NAND2_X2 U5495 ( .A1(n5322), .A2(n4445), .ZN(n5347) );
  INV_X4 U5496 ( .A(n5347), .ZN(n5323) );
  NAND2_X2 U5497 ( .A1(n5080), .A2(n5323), .ZN(n4500) );
  NAND2_X2 U5498 ( .A1(n5082), .A2(n4939), .ZN(n4502) );
  NAND2_X2 U5499 ( .A1(n4503), .A2(n4502), .ZN(n4858) );
  INV_X4 U5500 ( .A(regWrData[4]), .ZN(n4505) );
  NAND2_X2 U5501 ( .A1(n3183), .A2(memAddr[4]), .ZN(n4504) );
  INV_X4 U5502 ( .A(n5672), .ZN(n5662) );
  INV_X4 U5503 ( .A(regWrData[27]), .ZN(n4507) );
  NAND2_X2 U5504 ( .A1(n3183), .A2(memAddr[27]), .ZN(n4506) );
  NAND2_X2 U5505 ( .A1(n5173), .A2(n4616), .ZN(n5053) );
  INV_X4 U5506 ( .A(n5053), .ZN(n5101) );
  NAND2_X2 U5507 ( .A1(n5081), .A2(n5101), .ZN(n4508) );
  NAND2_X2 U5508 ( .A1(n2723), .A2(n2643), .ZN(n5159) );
  NAND2_X2 U5509 ( .A1(n3183), .A2(memAddr[12]), .ZN(n5158) );
  NAND2_X2 U5510 ( .A1(n5159), .A2(n5158), .ZN(n4512) );
  INV_X4 U5511 ( .A(n4512), .ZN(n4510) );
  NAND2_X2 U5512 ( .A1(n4510), .A2(n3185), .ZN(n4516) );
  INV_X4 U5513 ( .A(n4511), .ZN(n4513) );
  NAND2_X2 U5514 ( .A1(n4514), .A2(n2997), .ZN(n4515) );
  INV_X4 U5515 ( .A(n5404), .ZN(n5393) );
  NAND2_X2 U5516 ( .A1(n5080), .A2(n5393), .ZN(n4518) );
  NAND2_X2 U5517 ( .A1(n5226), .A2(n3041), .ZN(n5211) );
  INV_X4 U5518 ( .A(n5211), .ZN(n5207) );
  NAND2_X2 U5519 ( .A1(n5081), .A2(n5207), .ZN(n4517) );
  NAND2_X2 U5520 ( .A1(n4520), .A2(n4519), .ZN(n4782) );
  NAND2_X2 U5521 ( .A1(n4522), .A2(n4521), .ZN(n5939) );
  NAND2_X2 U5522 ( .A1(n6599), .A2(n3215), .ZN(n4544) );
  NAND2_X2 U5523 ( .A1(n4524), .A2(memAddr[0]), .ZN(n4532) );
  NAND2_X2 U5524 ( .A1(n3243), .A2(n4537), .ZN(n4526) );
  INV_X4 U5525 ( .A(n4526), .ZN(n4539) );
  INV_X4 U5526 ( .A(n5148), .ZN(n4527) );
  AOI22_X2 U5527 ( .A1(n4539), .A2(n4527), .B1(n5146), .B2(n4539), .ZN(n4543)
         );
  INV_X4 U5528 ( .A(n4528), .ZN(n4530) );
  NAND2_X2 U5529 ( .A1(n4532), .A2(n4531), .ZN(n5165) );
  NAND2_X2 U5530 ( .A1(n3243), .A2(n5165), .ZN(n4535) );
  NAND2_X2 U5531 ( .A1(n4535), .A2(n4534), .ZN(n4538) );
  NAND2_X2 U5532 ( .A1(n5145), .A2(n4539), .ZN(n4540) );
  INV_X4 U5533 ( .A(n6015), .ZN(n5969) );
  NAND2_X2 U5534 ( .A1(n5939), .A2(n5947), .ZN(n4749) );
  INV_X4 U5535 ( .A(n4544), .ZN(n6100) );
  MUX2_X2 U5536 ( .A(n3229), .B(n3224), .S(n4765), .Z(n4546) );
  INV_X4 U5537 ( .A(n4547), .ZN(n4548) );
  INV_X4 U5538 ( .A(regWrData[15]), .ZN(n4552) );
  NAND2_X2 U5539 ( .A1(n3183), .A2(memAddr[15]), .ZN(n4551) );
  NAND2_X2 U5540 ( .A1(n4790), .A2(n3041), .ZN(n4557) );
  INV_X4 U5541 ( .A(n4557), .ZN(n4818) );
  OAI21_X4 U5542 ( .B1(n6617), .B2(n2602), .A(n6618), .ZN(n5719) );
  XNOR2_X2 U5543 ( .A(n4553), .B(n3221), .ZN(n4558) );
  NAND2_X2 U5544 ( .A1(n4885), .A2(n4554), .ZN(n4801) );
  INV_X4 U5545 ( .A(n4801), .ZN(n4570) );
  NAND2_X2 U5546 ( .A1(n5393), .A2(n4555), .ZN(n5371) );
  NAND2_X2 U5547 ( .A1(n2723), .A2(n2642), .ZN(n4560) );
  NAND2_X2 U5548 ( .A1(n3183), .A2(memAddr[13]), .ZN(n4561) );
  NAND2_X2 U5549 ( .A1(n5386), .A2(n4616), .ZN(n5379) );
  INV_X4 U5550 ( .A(n5379), .ZN(n5369) );
  NAND2_X2 U5551 ( .A1(n5369), .A2(n4556), .ZN(n4791) );
  NAND2_X2 U5552 ( .A1(n5371), .A2(n4791), .ZN(n4803) );
  XNOR2_X2 U5553 ( .A(n4558), .B(n4557), .ZN(n5033) );
  INV_X4 U5554 ( .A(n4559), .ZN(n4563) );
  AOI21_X2 U5555 ( .B1(n4561), .B2(n4560), .A(zeroExt_2), .ZN(n4562) );
  XNOR2_X2 U5556 ( .A(n4565), .B(n3222), .ZN(n5374) );
  INV_X4 U5557 ( .A(n5374), .ZN(n4567) );
  XNOR2_X2 U5558 ( .A(n3134), .B(n3222), .ZN(n4566) );
  INV_X4 U5559 ( .A(n4791), .ZN(n4887) );
  INV_X4 U5560 ( .A(n4571), .ZN(n5886) );
  XNOR2_X2 U5561 ( .A(n5633), .B(n3222), .ZN(n4574) );
  INV_X4 U5562 ( .A(regWrData[9]), .ZN(n4573) );
  AOI22_X2 U5563 ( .A1(n2723), .A2(n2600), .B1(n3182), .B2(memAddr[9]), .ZN(
        n4572) );
  OAI21_X4 U5564 ( .B1(n4573), .B2(n3184), .A(n4572), .ZN(n5656) );
  NAND2_X2 U5565 ( .A1(n5656), .A2(n4445), .ZN(n5634) );
  XNOR2_X2 U5566 ( .A(n4574), .B(n5634), .ZN(n5651) );
  XNOR2_X2 U5567 ( .A(n5422), .B(n3221), .ZN(n4575) );
  INV_X4 U5568 ( .A(n5634), .ZN(n5631) );
  NAND2_X2 U5569 ( .A1(n5631), .A2(n4574), .ZN(n5339) );
  XNOR2_X2 U5570 ( .A(n4575), .B(n5423), .ZN(n5638) );
  NAND2_X2 U5571 ( .A1(n2723), .A2(n2644), .ZN(n5155) );
  NAND2_X2 U5572 ( .A1(n3183), .A2(memAddr[11]), .ZN(n5154) );
  NAND2_X2 U5573 ( .A1(n4579), .A2(n4578), .ZN(n4581) );
  NAND3_X2 U5574 ( .A1(n5154), .A2(n5155), .A3(n3185), .ZN(n4580) );
  OAI211_X2 U5575 ( .C1(n4582), .C2(n4581), .A(n4580), .B(n3041), .ZN(n5538)
         );
  XNOR2_X2 U5576 ( .A(n5538), .B(n3221), .ZN(n4583) );
  XNOR2_X2 U5577 ( .A(n4583), .B(n3061), .ZN(n5535) );
  INV_X4 U5578 ( .A(n4584), .ZN(n4601) );
  NAND2_X2 U5579 ( .A1(n3183), .A2(memAddr[7]), .ZN(n4585) );
  XNOR2_X2 U5580 ( .A(n3223), .B(n5492), .ZN(n4587) );
  NAND2_X2 U5581 ( .A1(n5489), .A2(n4587), .ZN(n5644) );
  XNOR2_X2 U5582 ( .A(n4593), .B(n4592), .ZN(n4594) );
  XNOR2_X2 U5583 ( .A(n4594), .B(n3222), .ZN(n5343) );
  NAND2_X2 U5584 ( .A1(n5323), .A2(n4595), .ZN(n5531) );
  XNOR2_X2 U5585 ( .A(n5554), .B(n3221), .ZN(n4656) );
  NAND2_X2 U5586 ( .A1(n5551), .A2(n4656), .ZN(n5643) );
  NAND2_X2 U5587 ( .A1(n5531), .A2(n5643), .ZN(n4596) );
  INV_X4 U5588 ( .A(n5538), .ZN(n5523) );
  XNOR2_X2 U5589 ( .A(n5392), .B(n5404), .ZN(n4597) );
  XNOR2_X2 U5590 ( .A(n4597), .B(n3221), .ZN(n5400) );
  INV_X4 U5591 ( .A(n5326), .ZN(n4600) );
  OAI21_X4 U5592 ( .B1(n4600), .B2(n4601), .A(n4599), .ZN(n4604) );
  XNOR2_X2 U5593 ( .A(n4602), .B(n3221), .ZN(n5639) );
  OAI21_X4 U5594 ( .B1(n4606), .B2(n5528), .A(n5530), .ZN(n4607) );
  NAND3_X4 U5595 ( .A1(n4661), .A2(n5032), .A3(n5531), .ZN(n5038) );
  INV_X4 U5596 ( .A(regWrData[16]), .ZN(n4609) );
  AOI22_X2 U5597 ( .A1(n2723), .A2(n2599), .B1(n3182), .B2(memAddr[16]), .ZN(
        n4608) );
  NAND2_X2 U5598 ( .A1(n2723), .A2(n2647), .ZN(n5143) );
  NAND2_X2 U5599 ( .A1(n3183), .A2(memAddr[1]), .ZN(n5142) );
  INV_X4 U5600 ( .A(n4612), .ZN(n4613) );
  INV_X4 U5601 ( .A(zeroExt_2), .ZN(n4616) );
  NAND2_X2 U5602 ( .A1(n4617), .A2(n4616), .ZN(n4618) );
  AOI21_X4 U5603 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n5600) );
  INV_X4 U5604 ( .A(n5600), .ZN(n4645) );
  XNOR2_X2 U5605 ( .A(n6040), .B(n3221), .ZN(n4646) );
  NAND2_X2 U5606 ( .A1(n5600), .A2(n4621), .ZN(n5572) );
  NAND2_X2 U5607 ( .A1(n3223), .A2(n3243), .ZN(n4629) );
  INV_X4 U5608 ( .A(n4629), .ZN(n4627) );
  NAND3_X4 U5609 ( .A1(n4624), .A2(n4165), .A3(n4623), .ZN(n4637) );
  INV_X4 U5610 ( .A(n4637), .ZN(n4625) );
  NAND4_X2 U5611 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4642)
         );
  NAND2_X2 U5612 ( .A1(n3243), .A2(n3222), .ZN(n4636) );
  XNOR2_X2 U5613 ( .A(n3222), .B(n2833), .ZN(n4634) );
  INV_X4 U5614 ( .A(n4636), .ZN(n4638) );
  INV_X4 U5615 ( .A(n4644), .ZN(n4798) );
  XNOR2_X2 U5616 ( .A(n4646), .B(n4645), .ZN(n5593) );
  INV_X4 U5617 ( .A(n5593), .ZN(n4649) );
  NAND2_X2 U5618 ( .A1(n6002), .A2(n6015), .ZN(n4648) );
  NAND2_X2 U5619 ( .A1(n5969), .A2(n3222), .ZN(n4647) );
  NAND2_X2 U5620 ( .A1(n4649), .A2(n5592), .ZN(n5573) );
  NAND2_X2 U5621 ( .A1(n4798), .A2(n5573), .ZN(n5664) );
  INV_X4 U5622 ( .A(regWrData[3]), .ZN(n4651) );
  NAND2_X2 U5623 ( .A1(n3183), .A2(memAddr[3]), .ZN(n4650) );
  OAI221_X2 U5624 ( .B1(n6572), .B2(n3155), .C1(n4651), .C2(n3184), .A(n4650), 
        .ZN(n5586) );
  INV_X4 U5625 ( .A(n5581), .ZN(n5569) );
  XNOR2_X2 U5626 ( .A(n3223), .B(n3156), .ZN(n4662) );
  NAND2_X2 U5627 ( .A1(n5569), .A2(n4662), .ZN(n5665) );
  XNOR2_X2 U5628 ( .A(n5661), .B(n3221), .ZN(n4652) );
  NAND2_X2 U5629 ( .A1(n5665), .A2(n5334), .ZN(n4667) );
  NAND2_X2 U5630 ( .A1(n3183), .A2(memAddr[5]), .ZN(n4653) );
  XNOR2_X2 U5631 ( .A(n2577), .B(n3221), .ZN(n4914) );
  INV_X4 U5632 ( .A(n5395), .ZN(n4655) );
  XNOR2_X2 U5633 ( .A(n4656), .B(n5555), .ZN(n5642) );
  FA_X1 U5634 ( .A(n3223), .B(n4935), .CI(n2577), .S(n4657) );
  INV_X4 U5635 ( .A(n4662), .ZN(n4663) );
  XNOR2_X2 U5636 ( .A(n4663), .B(n5569), .ZN(n5571) );
  XNOR2_X2 U5637 ( .A(n5611), .B(n5610), .ZN(n4664) );
  XNOR2_X2 U5638 ( .A(n4664), .B(n3221), .ZN(n4665) );
  NOR3_X4 U5639 ( .A1(n4668), .A2(n4667), .A3(n4655), .ZN(n4671) );
  XNOR2_X2 U5640 ( .A(n5672), .B(n3221), .ZN(n4669) );
  XNOR2_X2 U5641 ( .A(n4669), .B(n5661), .ZN(n5668) );
  INV_X4 U5642 ( .A(n5334), .ZN(n5329) );
  NOR3_X4 U5643 ( .A1(n5668), .A2(n4655), .A3(n5329), .ZN(n4670) );
  XNOR2_X2 U5644 ( .A(n2620), .B(n3221), .ZN(n4676) );
  XNOR2_X2 U5645 ( .A(n4676), .B(n4675), .ZN(n5942) );
  INV_X4 U5646 ( .A(n4770), .ZN(n4677) );
  AOI21_X4 U5647 ( .B1(n2895), .B2(n4678), .A(n4677), .ZN(n4681) );
  XNOR2_X2 U5648 ( .A(n4765), .B(n3221), .ZN(n4680) );
  XNOR2_X2 U5649 ( .A(n4681), .B(n4771), .ZN(n5961) );
  INV_X4 U5650 ( .A(n5961), .ZN(n4682) );
  NAND2_X2 U5651 ( .A1(n6005), .A2(n4682), .ZN(n4747) );
  NAND2_X2 U5652 ( .A1(n5505), .A2(n4855), .ZN(n4690) );
  NAND2_X2 U5653 ( .A1(n4929), .A2(n2620), .ZN(n4944) );
  NAND2_X2 U5654 ( .A1(n4966), .A2(n4818), .ZN(n4946) );
  NAND2_X2 U5655 ( .A1(n4683), .A2(n3157), .ZN(n4686) );
  NAND2_X2 U5656 ( .A1(n2836), .A2(n3156), .ZN(n4984) );
  INV_X4 U5657 ( .A(n4984), .ZN(n4684) );
  AOI21_X2 U5658 ( .B1(n4981), .B2(n4943), .A(n4684), .ZN(n4685) );
  NAND2_X2 U5659 ( .A1(n4867), .A2(n5451), .ZN(n4689) );
  AOI22_X2 U5660 ( .A1(n5514), .A2(n4858), .B1(n5695), .B2(n4782), .ZN(n4688)
         );
  NAND3_X2 U5661 ( .A1(n4690), .A2(n4689), .A3(n4688), .ZN(n5937) );
  INV_X4 U5662 ( .A(n6022), .ZN(n4961) );
  NAND2_X2 U5663 ( .A1(n5080), .A2(n5489), .ZN(n4694) );
  INV_X4 U5664 ( .A(regWrData[24]), .ZN(n4692) );
  NAND2_X2 U5665 ( .A1(n3182), .A2(memAddr[24]), .ZN(n4691) );
  NAND2_X2 U5666 ( .A1(n5825), .A2(n3041), .ZN(n5811) );
  INV_X4 U5667 ( .A(n5811), .ZN(n5807) );
  NAND2_X2 U5668 ( .A1(n5081), .A2(n5807), .ZN(n4693) );
  NAND3_X4 U5669 ( .A1(n4694), .A2(n3216), .A3(n4693), .ZN(n5706) );
  INV_X4 U5670 ( .A(n5706), .ZN(n4695) );
  NAND2_X2 U5671 ( .A1(n2680), .A2(regWrData[30]), .ZN(n4698) );
  NAND2_X2 U5672 ( .A1(n2723), .A2(n2640), .ZN(n4697) );
  NAND2_X2 U5673 ( .A1(n3183), .A2(memAddr[30]), .ZN(n4696) );
  NAND2_X2 U5674 ( .A1(n5262), .A2(n3041), .ZN(n5729) );
  INV_X4 U5675 ( .A(n5729), .ZN(n5722) );
  NAND2_X2 U5676 ( .A1(n5081), .A2(n5722), .ZN(n4700) );
  NAND2_X2 U5677 ( .A1(n5080), .A2(n5600), .ZN(n4699) );
  INV_X4 U5678 ( .A(regWrData[22]), .ZN(n4702) );
  NAND2_X2 U5679 ( .A1(n3183), .A2(memAddr[22]), .ZN(n4701) );
  OAI221_X2 U5680 ( .B1(n6580), .B2(n3155), .C1(n4702), .C2(n3184), .A(n4701), 
        .ZN(n5897) );
  NAND2_X2 U5681 ( .A1(n5897), .A2(n3041), .ZN(n5879) );
  INV_X4 U5682 ( .A(n5879), .ZN(n5875) );
  NAND2_X2 U5683 ( .A1(n5081), .A2(n5875), .ZN(n4704) );
  NAND3_X2 U5684 ( .A1(n4704), .A2(n3216), .A3(n4703), .ZN(n4973) );
  NAND2_X2 U5685 ( .A1(n5082), .A2(n4973), .ZN(n4705) );
  NAND2_X2 U5686 ( .A1(n4706), .A2(n4705), .ZN(n5353) );
  AOI22_X2 U5687 ( .A1(n4985), .A2(n5448), .B1(n5695), .B2(n5353), .ZN(n4729)
         );
  NAND2_X2 U5688 ( .A1(n3183), .A2(memAddr[26]), .ZN(n4707) );
  OAI221_X2 U5689 ( .B1(n6576), .B2(n3155), .C1(n4708), .C2(n3185), .A(n4707), 
        .ZN(n5190) );
  NAND2_X2 U5690 ( .A1(n5190), .A2(n3041), .ZN(n5004) );
  INV_X4 U5691 ( .A(n5004), .ZN(n5056) );
  NAND2_X2 U5692 ( .A1(n5081), .A2(n5056), .ZN(n4710) );
  NAND3_X2 U5693 ( .A1(n4710), .A2(n3216), .A3(n4709), .ZN(n4965) );
  AOI21_X2 U5694 ( .B1(n4981), .B2(n4965), .A(n2836), .ZN(n4716) );
  INV_X4 U5695 ( .A(regWrData[18]), .ZN(n4712) );
  NAND2_X2 U5696 ( .A1(n3183), .A2(memAddr[18]), .ZN(n4711) );
  OAI221_X2 U5697 ( .B1(n6584), .B2(n3155), .C1(n4712), .C2(n3184), .A(n4711), 
        .ZN(n5188) );
  NAND2_X2 U5698 ( .A1(n5081), .A2(n4837), .ZN(n4714) );
  NAND2_X2 U5699 ( .A1(n5082), .A2(n5281), .ZN(n4715) );
  NAND2_X2 U5700 ( .A1(n4716), .A2(n4715), .ZN(n4864) );
  NAND2_X2 U5701 ( .A1(n4867), .A2(n4864), .ZN(n4728) );
  INV_X4 U5702 ( .A(regWrData[28]), .ZN(n4718) );
  NAND2_X2 U5703 ( .A1(n3183), .A2(memAddr[28]), .ZN(n4717) );
  OAI221_X2 U5704 ( .B1(n6574), .B2(n3155), .C1(n4718), .C2(n3184), .A(n4717), 
        .ZN(n5174) );
  NAND2_X2 U5705 ( .A1(n5174), .A2(n3041), .ZN(n5099) );
  INV_X4 U5706 ( .A(n5099), .ZN(n5236) );
  NAND2_X2 U5707 ( .A1(n5081), .A2(n5236), .ZN(n4720) );
  NAND2_X2 U5708 ( .A1(n5080), .A2(n5569), .ZN(n4719) );
  NAND3_X2 U5709 ( .A1(n4720), .A2(n3216), .A3(n4719), .ZN(n4922) );
  AOI21_X2 U5710 ( .B1(n4981), .B2(n4922), .A(n2836), .ZN(n4726) );
  INV_X4 U5711 ( .A(regWrData[20]), .ZN(n4722) );
  NAND2_X2 U5712 ( .A1(n3182), .A2(memAddr[20]), .ZN(n4721) );
  NAND2_X2 U5713 ( .A1(n5172), .A2(n4445), .ZN(n4847) );
  INV_X4 U5714 ( .A(n4847), .ZN(n5017) );
  NAND2_X2 U5715 ( .A1(n5081), .A2(n5017), .ZN(n4724) );
  NAND2_X2 U5716 ( .A1(n5080), .A2(n5523), .ZN(n4723) );
  NAND2_X2 U5717 ( .A1(n5505), .A2(n4828), .ZN(n4727) );
  INV_X4 U5718 ( .A(n5387), .ZN(n4899) );
  OAI22_X2 U5719 ( .A1(n2626), .A2(n4898), .B1(n4899), .B2(n2778), .ZN(n4745)
         );
  NAND2_X2 U5720 ( .A1(n5081), .A2(n2620), .ZN(n4731) );
  INV_X4 U5721 ( .A(n4811), .ZN(n5357) );
  INV_X4 U5722 ( .A(n5277), .ZN(n4736) );
  NAND3_X4 U5723 ( .A1(n4737), .A2(n3216), .A3(n4738), .ZN(n4972) );
  NAND2_X2 U5724 ( .A1(n4972), .A2(n3157), .ZN(n4740) );
  NAND2_X2 U5725 ( .A1(n4981), .A2(n4973), .ZN(n4739) );
  NAND4_X2 U5726 ( .A1(n4746), .A2(n4748), .A3(n4747), .A4(n4749), .ZN(
        \ex_mem/N213 ) );
  MUX2_X2 U5727 ( .A(n3229), .B(n3224), .S(n4837), .Z(n4751) );
  NAND2_X2 U5728 ( .A1(n4751), .A2(n3226), .ZN(n4762) );
  INV_X4 U5729 ( .A(n4858), .ZN(n4752) );
  INV_X4 U5730 ( .A(n5430), .ZN(n4754) );
  INV_X4 U5731 ( .A(n6018), .ZN(n4960) );
  OAI22_X2 U5732 ( .A1(n4754), .A2(n2625), .B1(n2777), .B2(n4860), .ZN(n4755)
         );
  NOR3_X4 U5733 ( .A1(n4757), .A2(n4756), .A3(n4755), .ZN(n5412) );
  INV_X4 U5734 ( .A(n4758), .ZN(n4759) );
  XNOR2_X2 U5735 ( .A(n4763), .B(n3221), .ZN(n4764) );
  NAND2_X2 U5736 ( .A1(n4765), .A2(n4764), .ZN(n5013) );
  NAND2_X2 U5737 ( .A1(n4771), .A2(n4770), .ZN(n5015) );
  NAND2_X2 U5738 ( .A1(n4772), .A2(n4840), .ZN(n4775) );
  XNOR2_X2 U5739 ( .A(n4775), .B(n5011), .ZN(n5963) );
  NAND2_X2 U5740 ( .A1(n6005), .A2(n4776), .ZN(n4788) );
  NAND2_X2 U5741 ( .A1(n5505), .A2(n5451), .ZN(n4785) );
  NAND2_X2 U5742 ( .A1(n4966), .A2(n5369), .ZN(n4777) );
  NAND2_X2 U5743 ( .A1(n4778), .A2(n4777), .ZN(n4938) );
  NAND2_X2 U5744 ( .A1(n4981), .A2(n4939), .ZN(n4780) );
  NAND4_X2 U5745 ( .A1(n4781), .A2(n4984), .A3(n4780), .A4(n4779), .ZN(n5513)
         );
  NAND2_X2 U5746 ( .A1(n4867), .A2(n5513), .ZN(n4784) );
  NAND3_X2 U5747 ( .A1(n4785), .A2(n4784), .A3(n4783), .ZN(n5409) );
  AOI22_X2 U5748 ( .A1(n5947), .A2(n5387), .B1(n5938), .B2(n5409), .ZN(n4786)
         );
  NAND4_X2 U5749 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(
        \ex_mem/N214 ) );
  NAND2_X2 U5750 ( .A1(n4791), .A2(n5374), .ZN(n5034) );
  INV_X4 U5751 ( .A(n5034), .ZN(n4892) );
  INV_X4 U5752 ( .A(n4804), .ZN(n4807) );
  INV_X4 U5753 ( .A(n4792), .ZN(n4793) );
  INV_X4 U5754 ( .A(n5642), .ZN(n5338) );
  NAND2_X2 U5755 ( .A1(n5665), .A2(n5666), .ZN(n5333) );
  XNOR2_X2 U5756 ( .A(n5600), .B(n6040), .ZN(n4796) );
  XNOR2_X2 U5757 ( .A(n4796), .B(n3221), .ZN(n4797) );
  NAND2_X2 U5758 ( .A1(n4797), .A2(n5592), .ZN(n4799) );
  NAND3_X2 U5759 ( .A1(n4799), .A2(n5665), .A3(n4798), .ZN(n5330) );
  NAND2_X2 U5760 ( .A1(n4800), .A2(n4890), .ZN(n5373) );
  INV_X4 U5761 ( .A(n5372), .ZN(n4886) );
  NAND2_X2 U5762 ( .A1(n4804), .A2(n4803), .ZN(n4805) );
  MUX2_X2 U5763 ( .A(n3231), .B(n2844), .S(n4818), .Z(n4809) );
  NAND2_X2 U5764 ( .A1(n5505), .A2(n4864), .ZN(n4815) );
  NAND2_X2 U5765 ( .A1(n5514), .A2(n5353), .ZN(n4814) );
  NAND2_X2 U5766 ( .A1(n5695), .A2(n4828), .ZN(n4812) );
  NAND2_X2 U5767 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  AOI221_X2 U5768 ( .B1(n5948), .B2(n5939), .C1(n5947), .C2(n5937), .A(n4823), 
        .ZN(n4824) );
  NAND2_X2 U5769 ( .A1(n4825), .A2(n4824), .ZN(\ex_mem/N211 ) );
  MUX2_X2 U5770 ( .A(n3230), .B(n3224), .S(n5017), .Z(n4827) );
  NAND2_X2 U5771 ( .A1(n5127), .A2(n4828), .ZN(n4833) );
  NAND2_X2 U5772 ( .A1(n5505), .A2(n5353), .ZN(n4832) );
  INV_X4 U5773 ( .A(n5448), .ZN(n5354) );
  INV_X4 U5774 ( .A(n5544), .ZN(n5209) );
  INV_X4 U5775 ( .A(n4834), .ZN(n4835) );
  INV_X4 U5776 ( .A(n5916), .ZN(n5837) );
  OAI21_X4 U5777 ( .B1(n2849), .B2(n3112), .A(n5032), .ZN(n5838) );
  INV_X4 U5778 ( .A(n5219), .ZN(n5887) );
  NAND2_X2 U5779 ( .A1(n4837), .A2(n2724), .ZN(n5885) );
  INV_X4 U5780 ( .A(n5042), .ZN(n5218) );
  XNOR2_X2 U5781 ( .A(n3223), .B(n4838), .ZN(n4842) );
  INV_X4 U5782 ( .A(n5922), .ZN(n5832) );
  INV_X4 U5783 ( .A(n4840), .ZN(n4841) );
  XNOR2_X2 U5784 ( .A(n4842), .B(n5211), .ZN(n5223) );
  INV_X4 U5785 ( .A(n5223), .ZN(n5918) );
  XNOR2_X2 U5786 ( .A(n3223), .B(n4846), .ZN(n5016) );
  XNOR2_X2 U5787 ( .A(n5016), .B(n4847), .ZN(n5020) );
  INV_X4 U5788 ( .A(n5020), .ZN(n5831) );
  XNOR2_X2 U5789 ( .A(n4848), .B(n5831), .ZN(n5962) );
  INV_X4 U5790 ( .A(n5962), .ZN(n4849) );
  NAND2_X2 U5791 ( .A1(n6005), .A2(n4849), .ZN(n4875) );
  NAND2_X2 U5792 ( .A1(n4966), .A2(n5523), .ZN(n4850) );
  NAND4_X2 U5793 ( .A1(n4854), .A2(n4984), .A3(n4853), .A4(n4852), .ZN(n5512)
         );
  AOI22_X2 U5794 ( .A1(n4867), .A2(n5512), .B1(n5505), .B2(n5513), .ZN(n4857)
         );
  AOI22_X2 U5795 ( .A1(n5695), .A2(n5451), .B1(n5514), .B2(n4855), .ZN(n4856)
         );
  NAND2_X2 U5796 ( .A1(n4857), .A2(n4856), .ZN(n5929) );
  AOI22_X2 U5797 ( .A1(n3225), .A2(n5172), .B1(n5938), .B2(n5929), .ZN(n4874)
         );
  NAND2_X2 U5798 ( .A1(n5127), .A2(n4858), .ZN(n4863) );
  NAND2_X2 U5799 ( .A1(n5505), .A2(n5430), .ZN(n4862) );
  INV_X4 U5800 ( .A(n4860), .ZN(n5503) );
  NAND3_X2 U5801 ( .A1(n4863), .A2(n4862), .A3(n4861), .ZN(n5932) );
  NAND2_X2 U5802 ( .A1(n4864), .A2(n4985), .ZN(n4872) );
  INV_X4 U5803 ( .A(n6036), .ZN(n4867) );
  NAND2_X2 U5804 ( .A1(n4966), .A2(n5393), .ZN(n5686) );
  NAND2_X2 U5805 ( .A1(n5670), .A2(n4922), .ZN(n5689) );
  NAND2_X2 U5806 ( .A1(n4929), .A2(n5207), .ZN(n5687) );
  NAND4_X2 U5807 ( .A1(n5686), .A2(n3216), .A3(n5689), .A4(n5687), .ZN(n5078)
         );
  NAND2_X2 U5808 ( .A1(n5078), .A2(n3157), .ZN(n4866) );
  NAND3_X4 U5809 ( .A1(n4866), .A2(n4984), .A3(n4865), .ZN(n5435) );
  NAND2_X2 U5810 ( .A1(n4867), .A2(n5435), .ZN(n4871) );
  NOR2_X4 U5811 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  NAND3_X4 U5812 ( .A1(n4872), .A2(n4871), .A3(n4870), .ZN(n5546) );
  NAND4_X2 U5813 ( .A1(n4876), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(
        \ex_mem/N216 ) );
  INV_X4 U5814 ( .A(regWrData[14]), .ZN(n4879) );
  OAI211_X2 U5815 ( .C1(n4879), .C2(n3185), .A(n4878), .B(n4877), .ZN(n5197)
         );
  INV_X4 U5816 ( .A(n5197), .ZN(n4897) );
  MUX2_X2 U5817 ( .A(n3230), .B(n3224), .S(n4885), .Z(n4881) );
  INV_X4 U5818 ( .A(n4882), .ZN(n4906) );
  NAND2_X2 U5819 ( .A1(n4885), .A2(n4884), .ZN(n4905) );
  NOR2_X4 U5820 ( .A1(n4887), .A2(n4886), .ZN(n4894) );
  INV_X4 U5821 ( .A(n5371), .ZN(n4891) );
  NAND2_X2 U5822 ( .A1(n5371), .A2(n4888), .ZN(n4889) );
  OAI21_X4 U5823 ( .B1(n4891), .B2(n4890), .A(n4889), .ZN(n4893) );
  AOI21_X4 U5824 ( .B1(n4894), .B2(n4893), .A(n4892), .ZN(n4896) );
  AOI22_X2 U5825 ( .A1(n5938), .A2(n5939), .B1(n6005), .B2(n5989), .ZN(n4904)
         );
  OAI22_X2 U5826 ( .A1(n4898), .A2(n2778), .B1(n4897), .B2(n2592), .ZN(n4902)
         );
  INV_X4 U5827 ( .A(n5385), .ZN(n4900) );
  OAI22_X2 U5828 ( .A1(n4900), .A2(n2779), .B1(n4899), .B2(n2626), .ZN(n4901)
         );
  NAND4_X2 U5829 ( .A1(n4903), .A2(n4905), .A3(n4904), .A4(n4906), .ZN(
        \ex_mem/N210 ) );
  INV_X4 U5830 ( .A(n5940), .ZN(n5178) );
  INV_X4 U5831 ( .A(n5930), .ZN(n4907) );
  INV_X4 U5832 ( .A(n5897), .ZN(n4908) );
  INV_X4 U5833 ( .A(n5865), .ZN(n4909) );
  INV_X4 U5834 ( .A(n5825), .ZN(n5181) );
  INV_X4 U5835 ( .A(n5199), .ZN(n5799) );
  MUX2_X2 U5836 ( .A(n3230), .B(n3224), .S(n4911), .Z(n4912) );
  NAND2_X2 U5837 ( .A1(n4912), .A2(n3226), .ZN(n4920) );
  NAND2_X2 U5838 ( .A1(n4913), .A2(n5334), .ZN(n4915) );
  XNOR2_X2 U5839 ( .A(n4915), .B(n5328), .ZN(n5972) );
  INV_X4 U5840 ( .A(n5257), .ZN(n5446) );
  NAND2_X2 U5841 ( .A1(n5446), .A2(n5695), .ZN(n4927) );
  INV_X4 U5842 ( .A(n4923), .ZN(n5445) );
  NAND2_X2 U5843 ( .A1(n5445), .A2(n5505), .ZN(n4926) );
  INV_X4 U5844 ( .A(n4924), .ZN(n5447) );
  NAND2_X2 U5845 ( .A1(n5938), .A2(n5802), .ZN(n4992) );
  NAND2_X2 U5846 ( .A1(n5514), .A2(n5512), .ZN(n4958) );
  NAND2_X2 U5847 ( .A1(n5670), .A2(n4928), .ZN(n4931) );
  AOI22_X2 U5848 ( .A1(n4929), .A2(n5875), .B1(n4966), .B2(n5631), .ZN(n4930)
         );
  NAND3_X2 U5849 ( .A1(n4931), .A2(n3217), .A3(n4930), .ZN(n5310) );
  NAND2_X2 U5850 ( .A1(n5310), .A2(n3157), .ZN(n4933) );
  INV_X4 U5851 ( .A(n5511), .ZN(n4934) );
  NAND2_X2 U5852 ( .A1(n3156), .A2(n4938), .ZN(n4941) );
  NAND3_X4 U5853 ( .A1(n4942), .A2(n4941), .A3(n4940), .ZN(n5314) );
  INV_X4 U5854 ( .A(n4944), .ZN(n4945) );
  NAND2_X2 U5855 ( .A1(n4945), .A2(n3156), .ZN(n4955) );
  INV_X4 U5856 ( .A(n4946), .ZN(n4947) );
  NAND2_X2 U5857 ( .A1(n5082), .A2(n5807), .ZN(n4948) );
  NAND2_X2 U5858 ( .A1(n5082), .A2(n5489), .ZN(n4949) );
  NOR3_X4 U5859 ( .A1(n4952), .A2(n2853), .A3(n4951), .ZN(n4953) );
  NAND2_X2 U5860 ( .A1(n5429), .A2(n5505), .ZN(n4963) );
  NAND2_X2 U5861 ( .A1(n5695), .A2(n5260), .ZN(n4962) );
  INV_X4 U5862 ( .A(n2626), .ZN(n4989) );
  INV_X4 U5863 ( .A(n4965), .ZN(n5289) );
  NOR2_X4 U5864 ( .A1(n5289), .A2(n5661), .ZN(n4969) );
  NAND2_X2 U5865 ( .A1(n4966), .A2(n5323), .ZN(n5283) );
  NAND2_X2 U5866 ( .A1(n4967), .A2(n5283), .ZN(n4968) );
  NAND2_X2 U5867 ( .A1(n4981), .A2(n5281), .ZN(n4970) );
  INV_X4 U5868 ( .A(n4972), .ZN(n4978) );
  NAND2_X2 U5869 ( .A1(n2605), .A2(n4973), .ZN(n5266) );
  INV_X4 U5870 ( .A(n5265), .ZN(n5270) );
  NAND2_X2 U5871 ( .A1(n4976), .A2(n5081), .ZN(n5264) );
  INV_X4 U5872 ( .A(n5264), .ZN(n5269) );
  AOI22_X2 U5873 ( .A1(n5695), .A2(n5436), .B1(n4867), .B2(n5087), .ZN(n4988)
         );
  AOI22_X2 U5874 ( .A1(n4981), .A2(n5712), .B1(n2605), .B2(n5706), .ZN(n4982)
         );
  NAND2_X2 U5875 ( .A1(n5505), .A2(n5438), .ZN(n4987) );
  INV_X4 U5876 ( .A(n2777), .ZN(n4985) );
  NAND3_X4 U5877 ( .A1(n4988), .A2(n4987), .A3(n4986), .ZN(n4999) );
  AOI22_X2 U5878 ( .A1(n5681), .A2(n4989), .B1(n6029), .B2(n4999), .ZN(n4990)
         );
  NAND4_X2 U5879 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(
        \ex_mem/N200 ) );
  INV_X4 U5880 ( .A(n5190), .ZN(n4994) );
  MUX2_X2 U5881 ( .A(n3230), .B(n3224), .S(n5056), .Z(n4996) );
  INV_X4 U5882 ( .A(n4997), .ZN(n5052) );
  NAND2_X2 U5883 ( .A1(n5056), .A2(n4998), .ZN(n5051) );
  OAI22_X2 U5884 ( .A1(n4994), .A2(n2592), .B1(n5091), .B2(n2627), .ZN(n5002)
         );
  INV_X4 U5885 ( .A(n5681), .ZN(n5000) );
  XNOR2_X2 U5886 ( .A(n5003), .B(n3221), .ZN(n5054) );
  XNOR2_X2 U5887 ( .A(n5054), .B(n5004), .ZN(n5740) );
  XNOR2_X2 U5888 ( .A(n3223), .B(n5005), .ZN(n5007) );
  INV_X4 U5889 ( .A(n5007), .ZN(n5006) );
  XNOR2_X2 U5890 ( .A(n5007), .B(n5785), .ZN(n5030) );
  XNOR2_X2 U5891 ( .A(n5816), .B(n3221), .ZN(n5010) );
  INV_X4 U5892 ( .A(n5010), .ZN(n5008) );
  NAND2_X2 U5893 ( .A1(n5807), .A2(n5008), .ZN(n5060) );
  XNOR2_X2 U5894 ( .A(n5856), .B(n3221), .ZN(n5029) );
  INV_X4 U5895 ( .A(n5029), .ZN(n5009) );
  XNOR2_X2 U5896 ( .A(n5010), .B(n5811), .ZN(n5748) );
  INV_X4 U5897 ( .A(n5748), .ZN(n5823) );
  NAND2_X2 U5898 ( .A1(n2714), .A2(n5823), .ZN(n5059) );
  OAI22_X2 U5899 ( .A1(n5030), .A2(n5060), .B1(n5030), .B2(n5059), .ZN(n5241)
         );
  INV_X4 U5900 ( .A(n5920), .ZN(n5012) );
  NOR2_X4 U5901 ( .A1(n5223), .A2(n5012), .ZN(n5018) );
  INV_X4 U5902 ( .A(n5014), .ZN(n5040) );
  XNOR2_X2 U5903 ( .A(n3223), .B(n5019), .ZN(n5021) );
  XNOR2_X2 U5904 ( .A(n3223), .B(n3096), .ZN(n5023) );
  XNOR2_X2 U5905 ( .A(n5023), .B(n5879), .ZN(n5895) );
  INV_X4 U5906 ( .A(n5895), .ZN(n5846) );
  NAND2_X2 U5907 ( .A1(n5020), .A2(n5921), .ZN(n5925) );
  INV_X4 U5908 ( .A(n5021), .ZN(n5022) );
  INV_X4 U5909 ( .A(n5023), .ZN(n5024) );
  NAND2_X2 U5910 ( .A1(n5875), .A2(n5024), .ZN(n5836) );
  INV_X4 U5911 ( .A(n5836), .ZN(n5844) );
  OAI21_X4 U5912 ( .B1(n5028), .B2(n5027), .A(n5026), .ZN(n5817) );
  XNOR2_X2 U5913 ( .A(n5029), .B(n5701), .ZN(n5853) );
  INV_X4 U5914 ( .A(n5853), .ZN(n5818) );
  NAND2_X2 U5915 ( .A1(n5823), .A2(n5818), .ZN(n5057) );
  INV_X4 U5916 ( .A(n5057), .ZN(n5792) );
  INV_X4 U5917 ( .A(n5030), .ZN(n5796) );
  NAND2_X2 U5918 ( .A1(n5792), .A2(n5796), .ZN(n5031) );
  NOR2_X4 U5919 ( .A1(n5046), .A2(n5749), .ZN(n5820) );
  XNOR2_X2 U5920 ( .A(n5740), .B(n5048), .ZN(n6063) );
  NAND4_X2 U5921 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(
        \ex_mem/N222 ) );
  INV_X4 U5922 ( .A(n5173), .ZN(n5092) );
  XNOR2_X2 U5923 ( .A(n5100), .B(n5053), .ZN(n5103) );
  INV_X4 U5924 ( .A(n5103), .ZN(n5243) );
  INV_X4 U5925 ( .A(n5054), .ZN(n5055) );
  NAND2_X2 U5926 ( .A1(n5056), .A2(n5055), .ZN(n5102) );
  NAND2_X2 U5927 ( .A1(n5102), .A2(n5755), .ZN(n5469) );
  AOI21_X4 U5928 ( .B1(n5244), .B2(n5796), .A(n5061), .ZN(n5063) );
  INV_X4 U5929 ( .A(n5058), .ZN(n5061) );
  NAND2_X2 U5930 ( .A1(n5060), .A2(n5059), .ZN(n5791) );
  XNOR2_X2 U5931 ( .A(n5243), .B(n5066), .ZN(n6064) );
  MUX2_X2 U5932 ( .A(n3231), .B(n2844), .S(n5101), .Z(n5067) );
  NAND2_X2 U5933 ( .A1(n5101), .A2(n5069), .ZN(n5070) );
  NAND2_X2 U5934 ( .A1(n5446), .A2(n5505), .ZN(n5074) );
  NAND2_X2 U5935 ( .A1(n5445), .A2(n5127), .ZN(n5073) );
  NAND2_X2 U5936 ( .A1(n5616), .A2(n5261), .ZN(n5116) );
  NAND3_X2 U5937 ( .A1(n5074), .A2(n5073), .A3(n5116), .ZN(n5677) );
  INV_X4 U5938 ( .A(n5677), .ZN(n5075) );
  INV_X4 U5939 ( .A(n5078), .ZN(n5086) );
  NAND2_X2 U5940 ( .A1(n2605), .A2(n5079), .ZN(n5692) );
  NAND2_X2 U5941 ( .A1(n5082), .A2(n5080), .ZN(n5698) );
  INV_X4 U5942 ( .A(n5698), .ZN(n5304) );
  NAND2_X2 U5943 ( .A1(n5304), .A2(n5101), .ZN(n5691) );
  INV_X4 U5944 ( .A(n5691), .ZN(n5084) );
  NAND2_X2 U5945 ( .A1(n5082), .A2(n5081), .ZN(n5709) );
  INV_X4 U5946 ( .A(n5709), .ZN(n5303) );
  NAND2_X2 U5947 ( .A1(n5303), .A2(n5662), .ZN(n5693) );
  NAND2_X2 U5948 ( .A1(n5693), .A2(n5306), .ZN(n5083) );
  AOI22_X2 U5949 ( .A1(n4985), .A2(n5436), .B1(n5298), .B2(n4867), .ZN(n5089)
         );
  NAND2_X2 U5950 ( .A1(n5089), .A2(n5088), .ZN(n5680) );
  INV_X4 U5951 ( .A(n5680), .ZN(n5120) );
  NAND2_X2 U5952 ( .A1(n5947), .A2(n5681), .ZN(n5090) );
  NAND2_X2 U5953 ( .A1(n5097), .A2(n5096), .ZN(\ex_mem/N223 ) );
  INV_X4 U5954 ( .A(n5174), .ZN(n5098) );
  XNOR2_X2 U5955 ( .A(n3223), .B(n5114), .ZN(n5234) );
  XNOR2_X2 U5956 ( .A(n5234), .B(n5099), .ZN(n5737) );
  NAND2_X2 U5957 ( .A1(n5101), .A2(n3071), .ZN(n5237) );
  NAND2_X2 U5958 ( .A1(n5102), .A2(n5237), .ZN(n5104) );
  NAND2_X2 U5959 ( .A1(n5103), .A2(n5237), .ZN(n5741) );
  NAND2_X2 U5960 ( .A1(n5104), .A2(n5741), .ZN(n5754) );
  INV_X4 U5961 ( .A(n5241), .ZN(n5105) );
  INV_X4 U5962 ( .A(n5741), .ZN(n5106) );
  XNOR2_X2 U5963 ( .A(n5109), .B(n3057), .ZN(n6061) );
  INV_X4 U5964 ( .A(n6061), .ZN(n6048) );
  MUX2_X2 U5965 ( .A(n3231), .B(n2844), .S(n5236), .Z(n5110) );
  NAND2_X2 U5966 ( .A1(n5236), .A2(n5112), .ZN(n5113) );
  INV_X4 U5967 ( .A(n5260), .ZN(n5500) );
  OAI221_X2 U5968 ( .B1(n6036), .B2(n5499), .C1(n5500), .C2(n5510), .A(n5116), 
        .ZN(n5626) );
  INV_X4 U5969 ( .A(n5626), .ZN(n5482) );
  NAND2_X2 U5970 ( .A1(n3225), .A2(n5174), .ZN(n5119) );
  NAND2_X2 U5971 ( .A1(n5314), .A2(n5505), .ZN(n5130) );
  AOI22_X2 U5972 ( .A1(n2685), .A2(n5122), .B1(n2605), .B2(n5121), .ZN(n5126)
         );
  AOI221_X2 U5973 ( .B1(n5303), .B2(n5569), .C1(n5304), .C2(n5236), .A(n5711), 
        .ZN(n5125) );
  NAND2_X2 U5974 ( .A1(n3156), .A2(n5123), .ZN(n5124) );
  INV_X4 U5975 ( .A(n6036), .ZN(n5127) );
  NAND2_X2 U5976 ( .A1(n5947), .A2(n5677), .ZN(n5131) );
  INV_X4 U5977 ( .A(regWrData[2]), .ZN(n5140) );
  OAI211_X2 U5978 ( .C1(n5140), .C2(n3185), .A(n5139), .B(n5138), .ZN(n5624)
         );
  INV_X4 U5979 ( .A(n5624), .ZN(n5141) );
  INV_X4 U5980 ( .A(regWrData[1]), .ZN(n5144) );
  OAI211_X2 U5981 ( .C1(n5144), .C2(n3185), .A(n5143), .B(n5142), .ZN(n5195)
         );
  INV_X4 U5982 ( .A(n5195), .ZN(n5603) );
  INV_X4 U5983 ( .A(regWrData[0]), .ZN(n5152) );
  OAI211_X2 U5984 ( .C1(n5152), .C2(n3185), .A(n5151), .B(n5150), .ZN(n5186)
         );
  INV_X4 U5985 ( .A(n5186), .ZN(n6007) );
  INV_X4 U5986 ( .A(n5198), .ZN(n5561) );
  INV_X4 U5987 ( .A(n5656), .ZN(n5153) );
  INV_X4 U5988 ( .A(regWrData[11]), .ZN(n5156) );
  OAI211_X2 U5989 ( .C1(n5156), .C2(n3185), .A(n5155), .B(n5154), .ZN(n5545)
         );
  INV_X4 U5990 ( .A(n5545), .ZN(n5157) );
  INV_X4 U5991 ( .A(regWrData[12]), .ZN(n5160) );
  OAI211_X2 U5992 ( .C1(n5160), .C2(n3185), .A(n5159), .B(n5158), .ZN(n5410)
         );
  INV_X4 U5993 ( .A(n5410), .ZN(n5161) );
  INV_X4 U5994 ( .A(n5386), .ZN(n5162) );
  INV_X4 U5995 ( .A(n5187), .ZN(n5480) );
  INV_X4 U5996 ( .A(n5262), .ZN(n5163) );
  INV_X4 U5997 ( .A(n5185), .ZN(n5773) );
  NAND2_X2 U5998 ( .A1(n3194), .A2(n3028), .ZN(n5168) );
  NAND4_X2 U5999 ( .A1(n5169), .A2(n5168), .A3(n6433), .A4(n5167), .ZN(
        \id_ex/N37 ) );
  INV_X4 U6000 ( .A(n5170), .ZN(\id_ex/N30 ) );
  NAND4_X2 U6001 ( .A1(n5177), .A2(n5136), .A3(n5176), .A4(n5175), .ZN(n5206)
         );
  NAND4_X2 U6002 ( .A1(n5180), .A2(n4909), .A3(n5179), .A4(n5178), .ZN(n5184)
         );
  NAND2_X2 U6003 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  NAND4_X2 U6004 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n5205)
         );
  NAND4_X2 U6005 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n5204)
         );
  MUX2_X2 U6006 ( .A(n3230), .B(n3224), .S(n5207), .Z(n5208) );
  NAND2_X2 U6007 ( .A1(n5208), .A2(n3226), .ZN(n5215) );
  INV_X4 U6008 ( .A(n5210), .ZN(n5212) );
  XNOR2_X2 U6009 ( .A(n5224), .B(n5223), .ZN(n5964) );
  NAND2_X2 U6010 ( .A1(n6005), .A2(n5225), .ZN(n5231) );
  AOI22_X2 U6011 ( .A1(n3225), .A2(n5226), .B1(n5948), .B2(n5409), .ZN(n5230)
         );
  INV_X4 U6012 ( .A(n5546), .ZN(n5411) );
  NOR2_X4 U6013 ( .A1(n5411), .A2(n2627), .ZN(n5228) );
  NOR2_X4 U6014 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND4_X2 U6015 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(
        \ex_mem/N215 ) );
  XNOR2_X2 U6016 ( .A(n3223), .B(n5459), .ZN(n5238) );
  INV_X4 U6017 ( .A(n5238), .ZN(n5233) );
  NAND2_X2 U6018 ( .A1(n5236), .A2(n5235), .ZN(n5727) );
  XNOR2_X2 U6019 ( .A(n5238), .B(n5462), .ZN(n5731) );
  INV_X4 U6020 ( .A(n5240), .ZN(n5247) );
  INV_X4 U6021 ( .A(n5242), .ZN(n5245) );
  XOR2_X2 U6022 ( .A(n5729), .B(n3221), .Z(n5251) );
  XNOR2_X2 U6023 ( .A(n5251), .B(n5720), .ZN(n5723) );
  XNOR2_X2 U6024 ( .A(n5252), .B(n5723), .ZN(n6062) );
  INV_X4 U6025 ( .A(n6062), .ZN(n6047) );
  MUX2_X2 U6026 ( .A(n3231), .B(n2844), .S(n5722), .Z(n5253) );
  NAND2_X2 U6027 ( .A1(n5722), .A2(n5254), .ZN(n5255) );
  MUX2_X2 U6028 ( .A(n6016), .B(n5257), .S(n4867), .Z(n5601) );
  MUX2_X2 U6029 ( .A(n5261), .B(n5260), .S(n4867), .Z(n5772) );
  INV_X4 U6030 ( .A(n5772), .ZN(n5602) );
  NAND2_X2 U6031 ( .A1(n3225), .A2(n5262), .ZN(n5263) );
  NAND2_X2 U6032 ( .A1(n5265), .A2(n5264), .ZN(n5268) );
  INV_X4 U6033 ( .A(n5266), .ZN(n5267) );
  NAND2_X2 U6034 ( .A1(n5271), .A2(n5616), .ZN(n5272) );
  NAND2_X2 U6035 ( .A1(n5616), .A2(n2605), .ZN(n5276) );
  INV_X4 U6036 ( .A(n5283), .ZN(n5284) );
  NAND2_X2 U6037 ( .A1(n2908), .A2(n5284), .ZN(n5285) );
  NAND3_X2 U6038 ( .A1(n5287), .A2(n5286), .A3(n5285), .ZN(n5293) );
  NAND2_X2 U6039 ( .A1(n2908), .A2(n5670), .ZN(n5288) );
  AOI22_X2 U6040 ( .A1(n5304), .A2(n5458), .B1(n5303), .B2(n5611), .ZN(n5290)
         );
  OAI21_X4 U6041 ( .B1(n5296), .B2(n5295), .A(n5294), .ZN(n5297) );
  INV_X4 U6042 ( .A(n5297), .ZN(n6044) );
  NAND2_X2 U6043 ( .A1(n5514), .A2(n5438), .ZN(n5299) );
  NAND2_X2 U6044 ( .A1(n5303), .A2(n5600), .ZN(n5308) );
  NAND2_X2 U6045 ( .A1(n5304), .A2(n5722), .ZN(n5309) );
  NAND2_X2 U6046 ( .A1(n5695), .A2(n5314), .ZN(n6023) );
  INV_X4 U6047 ( .A(n5771), .ZN(n5315) );
  NAND2_X2 U6048 ( .A1(n5320), .A2(n5319), .ZN(\ex_mem/N226 ) );
  MUX2_X2 U6049 ( .A(n3230), .B(n3224), .S(n5323), .Z(n5324) );
  NAND2_X2 U6050 ( .A1(n5324), .A2(n3226), .ZN(n5351) );
  NAND2_X2 U6051 ( .A1(n2923), .A2(n5639), .ZN(n5342) );
  INV_X4 U6052 ( .A(n5328), .ZN(n5332) );
  AOI21_X4 U6053 ( .B1(n5330), .B2(n5668), .A(n5329), .ZN(n5331) );
  NOR2_X4 U6054 ( .A1(n5332), .A2(n5331), .ZN(n5337) );
  NAND2_X2 U6055 ( .A1(n5335), .A2(n5334), .ZN(n5336) );
  NAND3_X4 U6056 ( .A1(n5643), .A2(n5395), .A3(n5396), .ZN(n5533) );
  NAND2_X2 U6057 ( .A1(n5338), .A2(n5643), .ZN(n5525) );
  NAND2_X2 U6058 ( .A1(n5533), .A2(n5525), .ZN(n5498) );
  NAND2_X2 U6059 ( .A1(n2923), .A2(n5340), .ZN(n5341) );
  NAND2_X2 U6060 ( .A1(n4867), .A2(n5353), .ZN(n5356) );
  AOI22_X2 U6061 ( .A1(n5445), .A2(n5514), .B1(n5447), .B2(n5695), .ZN(n5355)
         );
  NAND3_X2 U6062 ( .A1(n5356), .A2(n2875), .A3(n5355), .ZN(n5905) );
  NAND2_X2 U6063 ( .A1(n5564), .A2(n5905), .ZN(n5366) );
  AOI22_X2 U6064 ( .A1(n2761), .A2(n2872), .B1(n6029), .B2(n5929), .ZN(n5365)
         );
  INV_X4 U6065 ( .A(n2627), .ZN(n5363) );
  NAND2_X2 U6066 ( .A1(n4867), .A2(n5436), .ZN(n5361) );
  NAND2_X2 U6067 ( .A1(n5505), .A2(n5435), .ZN(n5360) );
  NAND3_X4 U6068 ( .A1(n5362), .A2(n5361), .A3(n5360), .ZN(n5931) );
  AOI22_X2 U6069 ( .A1(n5363), .A2(n5932), .B1(n5947), .B2(n5931), .ZN(n5364)
         );
  NAND4_X2 U6070 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(
        \ex_mem/N206 ) );
  MUX2_X2 U6071 ( .A(n3230), .B(n3224), .S(n5369), .Z(n5370) );
  NAND2_X2 U6072 ( .A1(n5370), .A2(n3226), .ZN(n5383) );
  NAND3_X2 U6073 ( .A1(n5373), .A2(n5372), .A3(n5371), .ZN(n5375) );
  INV_X4 U6074 ( .A(n5378), .ZN(n5380) );
  NAND2_X2 U6075 ( .A1(n5564), .A2(n5384), .ZN(n5390) );
  AOI22_X2 U6076 ( .A1(n5938), .A2(n5387), .B1(n5947), .B2(n5409), .ZN(n5388)
         );
  NAND4_X2 U6077 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(
        \ex_mem/N209 ) );
  MUX2_X2 U6078 ( .A(n3230), .B(n3224), .S(n5393), .Z(n5394) );
  NAND2_X2 U6079 ( .A1(n5394), .A2(n3227), .ZN(n5408) );
  INV_X4 U6080 ( .A(n5553), .ZN(n5650) );
  INV_X4 U6081 ( .A(n5403), .ZN(n5405) );
  AOI22_X2 U6082 ( .A1(n3225), .A2(n5410), .B1(n6029), .B2(n5409), .ZN(n5416)
         );
  INV_X4 U6083 ( .A(n3092), .ZN(n5428) );
  MUX2_X2 U6084 ( .A(n3230), .B(n3224), .S(n5707), .Z(n5419) );
  NAND2_X2 U6085 ( .A1(n5419), .A2(n3227), .ZN(n5427) );
  NAND2_X2 U6086 ( .A1(n3092), .A2(n3231), .ZN(n5424) );
  INV_X4 U6087 ( .A(n5499), .ZN(n5429) );
  NAND2_X2 U6088 ( .A1(n5429), .A2(n4985), .ZN(n5433) );
  NAND2_X2 U6089 ( .A1(n5503), .A2(n5505), .ZN(n5432) );
  NAND2_X2 U6090 ( .A1(n5127), .A2(n5430), .ZN(n5431) );
  NAND4_X2 U6091 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n5653)
         );
  NAND2_X2 U6092 ( .A1(n5938), .A2(n5653), .ZN(n5456) );
  INV_X4 U6093 ( .A(n5435), .ZN(n5443) );
  INV_X4 U6094 ( .A(n5436), .ZN(n5437) );
  INV_X4 U6095 ( .A(n5438), .ZN(n5439) );
  NOR2_X4 U6096 ( .A1(n5439), .A2(n6036), .ZN(n5440) );
  NOR2_X4 U6097 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  AOI22_X2 U6098 ( .A1(n5446), .A2(n5514), .B1(n5445), .B2(n5695), .ZN(n5450)
         );
  AOI22_X2 U6099 ( .A1(n4867), .A2(n5448), .B1(n5447), .B2(n5505), .ZN(n5449)
         );
  NAND2_X2 U6100 ( .A1(n5450), .A2(n5449), .ZN(n5868) );
  AOI22_X2 U6101 ( .A1(n4867), .A2(n5511), .B1(n5505), .B2(n5512), .ZN(n5453)
         );
  AOI22_X2 U6102 ( .A1(n5695), .A2(n5513), .B1(n5514), .B2(n5451), .ZN(n5452)
         );
  NAND2_X2 U6103 ( .A1(n5453), .A2(n5452), .ZN(n5898) );
  AOI22_X2 U6104 ( .A1(n5868), .A2(n4989), .B1(n6029), .B2(n5898), .ZN(n5454)
         );
  NAND4_X2 U6105 ( .A1(n5455), .A2(n5456), .A3(n5457), .A4(n5454), .ZN(
        \ex_mem/N204 ) );
  MUX2_X2 U6106 ( .A(n3230), .B(n3224), .S(n5458), .Z(n5460) );
  INV_X4 U6107 ( .A(n5461), .ZN(n5488) );
  NAND2_X2 U6108 ( .A1(n5458), .A2(n5464), .ZN(n5487) );
  INV_X4 U6109 ( .A(n5601), .ZN(n5479) );
  NAND2_X2 U6110 ( .A1(n3089), .A2(n5796), .ZN(n5471) );
  NAND2_X2 U6111 ( .A1(n5471), .A2(n5472), .ZN(n5473) );
  NAND3_X2 U6112 ( .A1(n5473), .A2(n5817), .A3(n5792), .ZN(n5476) );
  INV_X4 U6113 ( .A(n5791), .ZN(n5763) );
  NAND2_X2 U6114 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  XNOR2_X2 U6115 ( .A(n5478), .B(n5731), .ZN(n6068) );
  INV_X4 U6116 ( .A(n5623), .ZN(n5481) );
  OAI22_X2 U6117 ( .A1(n5301), .A2(n2627), .B1(n5482), .B2(n2779), .ZN(n5483)
         );
  NAND4_X2 U6118 ( .A1(n5485), .A2(n5487), .A3(n5486), .A4(n5488), .ZN(
        \ex_mem/N225 ) );
  MUX2_X2 U6119 ( .A(n3230), .B(n3224), .S(n5489), .Z(n5491) );
  INV_X4 U6120 ( .A(n5493), .ZN(n5495) );
  XNOR2_X2 U6121 ( .A(n5498), .B(n5639), .ZN(n5978) );
  AOI22_X2 U6122 ( .A1(n5505), .A2(n5504), .B1(n5503), .B2(n5127), .ZN(n5506)
         );
  NAND2_X2 U6123 ( .A1(n5507), .A2(n5506), .ZN(n5783) );
  AOI22_X2 U6124 ( .A1(n5978), .A2(n6005), .B1(n5564), .B2(n5783), .ZN(n5521)
         );
  NAND2_X2 U6125 ( .A1(n5695), .A2(n5512), .ZN(n5516) );
  NAND2_X2 U6126 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  NAND4_X2 U6127 ( .A1(n5518), .A2(n5517), .A3(n5516), .A4(n5515), .ZN(n5826)
         );
  AOI22_X2 U6128 ( .A1(n5363), .A2(n5868), .B1(n5947), .B2(n5826), .ZN(n5519)
         );
  NAND4_X2 U6129 ( .A1(n5520), .A2(n5521), .A3(n5522), .A4(n5519), .ZN(
        \ex_mem/N203 ) );
  MUX2_X2 U6130 ( .A(n3230), .B(n3224), .S(n5523), .Z(n5524) );
  NAND2_X2 U6131 ( .A1(n5524), .A2(n3226), .ZN(n5542) );
  INV_X4 U6132 ( .A(n5525), .ZN(n5529) );
  AOI21_X4 U6133 ( .B1(n5534), .B2(n5533), .A(n5532), .ZN(n5536) );
  XNOR2_X2 U6134 ( .A(n5536), .B(n2591), .ZN(n5977) );
  INV_X4 U6135 ( .A(n5537), .ZN(n5539) );
  NAND2_X2 U6136 ( .A1(n5938), .A2(n5544), .ZN(n5549) );
  AOI22_X2 U6137 ( .A1(n3225), .A2(n5545), .B1(n5947), .B2(n5929), .ZN(n5548)
         );
  AOI22_X2 U6138 ( .A1(n6029), .A2(n5546), .B1(n5948), .B2(n5932), .ZN(n5547)
         );
  NAND4_X2 U6139 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(
        \ex_mem/N207 ) );
  INV_X4 U6140 ( .A(n5554), .ZN(n5560) );
  MUX2_X2 U6141 ( .A(n3230), .B(n3224), .S(n5551), .Z(n5552) );
  NAND2_X2 U6142 ( .A1(n5552), .A2(n3227), .ZN(n5559) );
  NAND2_X2 U6143 ( .A1(n5554), .A2(n3231), .ZN(n5556) );
  NAND2_X2 U6144 ( .A1(n5938), .A2(n5783), .ZN(n5567) );
  INV_X4 U6145 ( .A(n2626), .ZN(n5564) );
  AOI22_X2 U6146 ( .A1(n5802), .A2(n5564), .B1(n6029), .B2(n5826), .ZN(n5565)
         );
  NAND4_X2 U6147 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(
        \ex_mem/N202 ) );
  MUX2_X2 U6148 ( .A(n3230), .B(n3224), .S(n5569), .Z(n5570) );
  NAND2_X2 U6149 ( .A1(n5570), .A2(n3227), .ZN(n5585) );
  NAND2_X2 U6150 ( .A1(n5573), .A2(n5572), .ZN(n5614) );
  INV_X4 U6151 ( .A(n5613), .ZN(n5577) );
  AOI21_X2 U6152 ( .B1(n5614), .B2(n5577), .A(n5576), .ZN(n5578) );
  XNOR2_X2 U6153 ( .A(n5579), .B(n5578), .ZN(n5973) );
  INV_X4 U6154 ( .A(n5580), .ZN(n5582) );
  NAND2_X2 U6155 ( .A1(n5948), .A2(n5626), .ZN(n5589) );
  AOI22_X2 U6156 ( .A1(n5363), .A2(n5677), .B1(n5947), .B2(n5623), .ZN(n5587)
         );
  NAND4_X2 U6157 ( .A1(n5587), .A2(n5589), .A3(n5588), .A4(n5590), .ZN(
        \ex_mem/N198 ) );
  MUX2_X2 U6158 ( .A(n3224), .B(n3229), .S(n6037), .Z(n5591) );
  NAND2_X2 U6159 ( .A1(n5591), .A2(n3226), .ZN(n5599) );
  INV_X4 U6160 ( .A(n5970), .ZN(n5594) );
  INV_X4 U6161 ( .A(n5596), .ZN(n5597) );
  NAND2_X2 U6162 ( .A1(n5938), .A2(n5479), .ZN(n5608) );
  NAND4_X2 U6163 ( .A1(n5606), .A2(n5608), .A3(n5607), .A4(n5609), .ZN(
        \ex_mem/N196 ) );
  MUX2_X2 U6164 ( .A(n3230), .B(n3224), .S(n5611), .Z(n5612) );
  NAND2_X2 U6165 ( .A1(n5612), .A2(n3226), .ZN(n5622) );
  XNOR2_X2 U6166 ( .A(n5614), .B(n5613), .ZN(n5971) );
  INV_X4 U6167 ( .A(n5971), .ZN(n5615) );
  INV_X4 U6168 ( .A(n5617), .ZN(n5619) );
  NAND2_X2 U6169 ( .A1(n5948), .A2(n5479), .ZN(n5629) );
  AOI22_X2 U6170 ( .A1(n3225), .A2(n5624), .B1(n6029), .B2(n5623), .ZN(n5628)
         );
  NAND4_X2 U6171 ( .A1(n5628), .A2(n5629), .A3(n5630), .A4(n5627), .ZN(
        \ex_mem/N197 ) );
  MUX2_X2 U6172 ( .A(n3229), .B(n3224), .S(n5631), .Z(n5632) );
  INV_X4 U6173 ( .A(n5641), .ZN(n5646) );
  NAND2_X2 U6174 ( .A1(n5646), .A2(n5642), .ZN(n5649) );
  NAND2_X2 U6175 ( .A1(n5646), .A2(n5645), .ZN(n5648) );
  XNOR2_X2 U6176 ( .A(n5652), .B(n5651), .ZN(n5982) );
  INV_X4 U6177 ( .A(n5653), .ZN(n5877) );
  AOI22_X2 U6178 ( .A1(n3225), .A2(n5656), .B1(n6029), .B2(n5931), .ZN(n5658)
         );
  AOI22_X2 U6179 ( .A1(n5363), .A2(n5905), .B1(n5947), .B2(n5898), .ZN(n5657)
         );
  NAND4_X2 U6180 ( .A1(n5660), .A2(n5659), .A3(n5658), .A4(n5657), .ZN(
        \ex_mem/N205 ) );
  MUX2_X2 U6181 ( .A(n3230), .B(n3224), .S(n5662), .Z(n5663) );
  NAND2_X2 U6182 ( .A1(n5663), .A2(n3226), .ZN(n5676) );
  INV_X4 U6183 ( .A(n5664), .ZN(n5667) );
  INV_X4 U6184 ( .A(n5671), .ZN(n5673) );
  NAND2_X2 U6185 ( .A1(n5948), .A2(n5677), .ZN(n5684) );
  AOI22_X2 U6186 ( .A1(n5363), .A2(n5681), .B1(n5947), .B2(n5680), .ZN(n5682)
         );
  NAND4_X2 U6187 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(
        \ex_mem/N199 ) );
  NAND4_X2 U6188 ( .A1(n5687), .A2(n5686), .A3(n5691), .A4(n5693), .ZN(n5697)
         );
  NAND3_X2 U6189 ( .A1(n5689), .A2(n3217), .A3(n5692), .ZN(n5696) );
  NAND4_X2 U6190 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n5694)
         );
  OAI211_X2 U6191 ( .C1(n5697), .C2(n5696), .A(n5695), .B(n5694), .ZN(n6042)
         );
  NAND3_X2 U6192 ( .A1(n5715), .A2(n5714), .A3(n5713), .ZN(n6039) );
  NAND2_X2 U6193 ( .A1(n5127), .A2(n6039), .ZN(n6043) );
  AOI22_X2 U6194 ( .A1(n5717), .A2(n2844), .B1(n5938), .B2(n5716), .ZN(n5780)
         );
  INV_X4 U6195 ( .A(n6091), .ZN(n6088) );
  XNOR2_X2 U6196 ( .A(n2622), .B(n3221), .ZN(n5764) );
  INV_X4 U6197 ( .A(n5754), .ZN(n5733) );
  XNOR2_X2 U6198 ( .A(n5720), .B(n3221), .ZN(n5730) );
  INV_X4 U6199 ( .A(n5730), .ZN(n5721) );
  NAND2_X2 U6200 ( .A1(n5722), .A2(n5721), .ZN(n5726) );
  INV_X4 U6201 ( .A(n5726), .ZN(n5724) );
  OAI21_X4 U6202 ( .B1(n5728), .B2(n2990), .A(n5727), .ZN(n5732) );
  NAND2_X2 U6203 ( .A1(n5730), .A2(n5729), .ZN(n5735) );
  NAND3_X4 U6204 ( .A1(n5732), .A2(n5735), .A3(n5734), .ZN(n5756) );
  INV_X4 U6205 ( .A(n5756), .ZN(n5739) );
  NOR2_X4 U6206 ( .A1(n5733), .A2(n5739), .ZN(n5746) );
  INV_X4 U6207 ( .A(n5735), .ZN(n5736) );
  NOR2_X4 U6208 ( .A1(n5739), .A2(n5743), .ZN(n5745) );
  OAI21_X4 U6209 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(n5757) );
  NAND2_X2 U6210 ( .A1(n5757), .A2(n5796), .ZN(n5765) );
  NAND2_X2 U6211 ( .A1(n5753), .A2(n5752), .ZN(n5762) );
  NAND2_X2 U6212 ( .A1(n5758), .A2(n5757), .ZN(n5769) );
  AOI21_X4 U6213 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n6050) );
  NAND2_X2 U6214 ( .A1(n5763), .A2(n5764), .ZN(n5767) );
  NAND2_X2 U6215 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NAND2_X2 U6216 ( .A1(n6050), .A2(n6049), .ZN(n6084) );
  AOI22_X2 U6217 ( .A1(n3231), .A2(n6075), .B1(n5948), .B2(n5771), .ZN(n5778)
         );
  NAND4_X2 U6218 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(
        \ex_mem/N227 ) );
  MUX2_X2 U6219 ( .A(n3230), .B(n3224), .S(n5781), .Z(n5782) );
  NAND2_X2 U6220 ( .A1(n5782), .A2(n3226), .ZN(n5789) );
  INV_X4 U6221 ( .A(n5783), .ZN(n5809) );
  INV_X4 U6222 ( .A(n5784), .ZN(n5786) );
  XNOR2_X2 U6223 ( .A(n5795), .B(n5796), .ZN(n5996) );
  NAND2_X2 U6224 ( .A1(n6005), .A2(n5797), .ZN(n5805) );
  AOI22_X2 U6225 ( .A1(n6029), .A2(n5802), .B1(n5948), .B2(n5826), .ZN(n5803)
         );
  NAND4_X2 U6226 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(
        \ex_mem/N221 ) );
  MUX2_X2 U6227 ( .A(n3229), .B(n3224), .S(n5807), .Z(n5808) );
  NAND2_X2 U6228 ( .A1(n5808), .A2(n3226), .ZN(n5815) );
  NOR2_X4 U6229 ( .A1(n5809), .A2(n2778), .ZN(n5814) );
  INV_X4 U6230 ( .A(n5810), .ZN(n5812) );
  AOI21_X4 U6231 ( .B1(n5821), .B2(n5820), .A(n5819), .ZN(n5822) );
  XNOR2_X2 U6232 ( .A(n5823), .B(n5822), .ZN(n5997) );
  NAND2_X2 U6233 ( .A1(n6005), .A2(n5824), .ZN(n5829) );
  AOI22_X2 U6234 ( .A1(n5947), .A2(n5868), .B1(n5938), .B2(n5826), .ZN(n5827)
         );
  NAND4_X2 U6235 ( .A1(n5828), .A2(n5829), .A3(n5830), .A4(n5827), .ZN(
        \ex_mem/N220 ) );
  NAND2_X2 U6236 ( .A1(n5835), .A2(n5928), .ZN(n5890) );
  INV_X4 U6237 ( .A(n5841), .ZN(n5842) );
  NAND3_X2 U6238 ( .A1(n5850), .A2(n5849), .A3(n5848), .ZN(n5851) );
  XNOR2_X2 U6239 ( .A(n5854), .B(n5853), .ZN(n6065) );
  MUX2_X2 U6240 ( .A(n3231), .B(n2844), .S(n5858), .Z(n5855) );
  NAND2_X2 U6241 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  NAND2_X2 U6242 ( .A1(n3225), .A2(n5865), .ZN(n5866) );
  INV_X4 U6243 ( .A(n5898), .ZN(n5870) );
  NAND2_X2 U6244 ( .A1(n6029), .A2(n5868), .ZN(n5869) );
  MUX2_X2 U6245 ( .A(n3229), .B(n3224), .S(n5875), .Z(n5876) );
  NAND2_X2 U6246 ( .A1(n5876), .A2(n3226), .ZN(n5883) );
  INV_X4 U6247 ( .A(n5878), .ZN(n5880) );
  XNOR2_X2 U6248 ( .A(n5895), .B(n5894), .ZN(n5990) );
  NAND2_X2 U6249 ( .A1(n6005), .A2(n5896), .ZN(n5901) );
  AOI22_X2 U6250 ( .A1(n3225), .A2(n5897), .B1(n5948), .B2(n5931), .ZN(n5900)
         );
  AOI22_X2 U6251 ( .A1(n5947), .A2(n5905), .B1(n5938), .B2(n5898), .ZN(n5899)
         );
  NAND4_X2 U6252 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(
        \ex_mem/N218 ) );
  MUX2_X2 U6253 ( .A(n3229), .B(n3224), .S(n5903), .Z(n5904) );
  NAND2_X2 U6254 ( .A1(n5904), .A2(n3226), .ZN(n5912) );
  INV_X4 U6255 ( .A(n5905), .ZN(n5906) );
  INV_X4 U6256 ( .A(n5907), .ZN(n5909) );
  OAI211_X2 U6257 ( .C1(n5926), .C2(n5892), .A(n5925), .B(n5924), .ZN(n5927)
         );
  XNOR2_X2 U6258 ( .A(n5927), .B(n5928), .ZN(n5958) );
  AOI22_X2 U6259 ( .A1(n3225), .A2(n5930), .B1(n5948), .B2(n5929), .ZN(n5934)
         );
  AOI22_X2 U6260 ( .A1(n5947), .A2(n5932), .B1(n5938), .B2(n5931), .ZN(n5933)
         );
  NAND4_X2 U6261 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(
        \ex_mem/N217 ) );
  NAND2_X2 U6262 ( .A1(n3225), .A2(n5940), .ZN(n5956) );
  XNOR2_X2 U6263 ( .A(n5943), .B(n5942), .ZN(n5968) );
  INV_X4 U6264 ( .A(n5968), .ZN(n5946) );
  MUX2_X2 U6265 ( .A(n3231), .B(n2844), .S(n2620), .Z(n5944) );
  NAND2_X2 U6266 ( .A1(n2620), .A2(n5950), .ZN(n5951) );
  NAND3_X2 U6267 ( .A1(n5957), .A2(n5956), .A3(n5955), .ZN(\ex_mem/N212 ) );
  NOR3_X4 U6268 ( .A1(n5965), .A2(n5966), .A3(n5967), .ZN(n6060) );
  XNOR2_X2 U6269 ( .A(n5969), .B(n6002), .ZN(n6004) );
  NAND4_X2 U6270 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n5981)
         );
  INV_X4 U6271 ( .A(n5976), .ZN(n5980) );
  INV_X4 U6272 ( .A(n5977), .ZN(n5979) );
  INV_X4 U6273 ( .A(n5982), .ZN(n5983) );
  NAND4_X2 U6274 ( .A1(n5946), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n5994)
         );
  NOR2_X4 U6275 ( .A1(n5994), .A2(n5993), .ZN(n6059) );
  NAND2_X2 U6276 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  INV_X4 U6277 ( .A(n5998), .ZN(n6070) );
  NAND2_X2 U6278 ( .A1(n6617), .A2(setInv_2), .ZN(n6087) );
  NAND3_X4 U6279 ( .A1(setInv_2), .A2(n2622), .A3(n6049), .ZN(n6000) );
  NAND3_X4 U6280 ( .A1(n6001), .A2(n6087), .A3(n6000), .ZN(n6057) );
  MUX2_X2 U6281 ( .A(n2776), .B(n3224), .S(n6002), .Z(n6003) );
  NAND2_X2 U6282 ( .A1(n6003), .A2(n3227), .ZN(n6014) );
  NAND2_X2 U6283 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  OAI221_X2 U6284 ( .B1(n6007), .B2(n2592), .C1(n6016), .C2(n2626), .A(n6006), 
        .ZN(n6013) );
  INV_X4 U6285 ( .A(n6009), .ZN(n6011) );
  INV_X4 U6286 ( .A(n6023), .ZN(n6026) );
  OAI21_X4 U6287 ( .B1(n6026), .B2(n6025), .A(n6029), .ZN(n6033) );
  INV_X4 U6288 ( .A(n6027), .ZN(n6031) );
  INV_X4 U6289 ( .A(n6028), .ZN(n6030) );
  INV_X4 U6290 ( .A(n2584), .ZN(n6103) );
  NAND2_X2 U6291 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  OAI21_X4 U6292 ( .B1(n6040), .B2(n6039), .A(n6038), .ZN(n6041) );
  AOI21_X2 U6293 ( .B1(n6041), .B2(n6042), .A(n2779), .ZN(n6046) );
  NAND3_X2 U6294 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n6045) );
  NOR2_X4 U6295 ( .A1(n6048), .A2(n6047), .ZN(n6054) );
  AOI21_X4 U6296 ( .B1(n6054), .B2(n6053), .A(n6052), .ZN(n6055) );
  AOI211_X4 U6297 ( .C1(n6058), .C2(n6057), .A(n6056), .B(n6055), .ZN(n6108)
         );
  NAND2_X2 U6298 ( .A1(n6062), .A2(n6061), .ZN(n6073) );
  INV_X4 U6299 ( .A(n6068), .ZN(n6069) );
  NAND2_X2 U6300 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND3_X2 U6301 ( .A1(n6086), .A2(n6603), .A3(n2622), .ZN(n6082) );
  NAND2_X2 U6302 ( .A1(setInv_2), .A2(n6603), .ZN(n6078) );
  NAND2_X2 U6303 ( .A1(n6091), .A2(n2787), .ZN(n6076) );
  INV_X4 U6304 ( .A(n2622), .ZN(n6075) );
  NAND2_X2 U6305 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  OAI21_X4 U6306 ( .B1(n6083), .B2(n6082), .A(n6081), .ZN(n6107) );
  INV_X4 U6307 ( .A(n6087), .ZN(n6085) );
  NAND3_X2 U6308 ( .A1(n6086), .A2(n2622), .A3(n6089), .ZN(n6098) );
  INV_X4 U6309 ( .A(n6089), .ZN(n6090) );
  NAND3_X2 U6310 ( .A1(n6099), .A2(n6098), .A3(n6097), .ZN(n6105) );
  NAND3_X2 U6311 ( .A1(n6103), .A2(n6102), .A3(n6101), .ZN(n6104) );
  NAND2_X2 U6312 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  OAI222_X2 U6313 ( .A1(n6140), .A2(n3239), .B1(n3242), .B2(n2668), .C1(n3237), 
        .C2(n6299), .ZN(memWrData[16]) );
  OAI222_X2 U6314 ( .A1(n6166), .A2(n3239), .B1(n3241), .B2(n2670), .C1(n3237), 
        .C2(n6172), .ZN(memWrData[17]) );
  OAI222_X2 U6315 ( .A1(n6167), .A2(n3239), .B1(n3242), .B2(n2701), .C1(n3237), 
        .C2(n6173), .ZN(memWrData[18]) );
  OAI222_X2 U6316 ( .A1(n6161), .A2(n3239), .B1(n3241), .B2(n3124), .C1(n3237), 
        .C2(n6258), .ZN(memWrData[19]) );
  OAI222_X2 U6317 ( .A1(n6168), .A2(n3239), .B1(n3242), .B2(n2699), .C1(n3237), 
        .C2(n6175), .ZN(memWrData[20]) );
  OAI222_X2 U6318 ( .A1(n6141), .A2(n3239), .B1(n3241), .B2(n2719), .C1(n3237), 
        .C2(n6298), .ZN(memWrData[21]) );
  OAI222_X2 U6319 ( .A1(n6142), .A2(n3239), .B1(n3242), .B2(n2687), .C1(n3237), 
        .C2(n6297), .ZN(memWrData[22]) );
  OAI222_X2 U6320 ( .A1(n6143), .A2(n3239), .B1(n3242), .B2(n2707), .C1(n3237), 
        .C2(n6296), .ZN(memWrData[23]) );
  OAI222_X2 U6321 ( .A1(n6144), .A2(n3239), .B1(n3242), .B2(n2667), .C1(n3237), 
        .C2(n6295), .ZN(memWrData[24]) );
  OAI222_X2 U6322 ( .A1(n6145), .A2(n3239), .B1(n3242), .B2(n2703), .C1(n3237), 
        .C2(n6294), .ZN(memWrData[25]) );
  OAI222_X2 U6323 ( .A1(n6169), .A2(n3239), .B1(n3242), .B2(n2665), .C1(n3237), 
        .C2(n6180), .ZN(memWrData[26]) );
  OAI222_X2 U6324 ( .A1(n6170), .A2(n3240), .B1(n3241), .B2(n2666), .C1(n3238), 
        .C2(n6181), .ZN(memWrData[27]) );
  OAI222_X2 U6325 ( .A1(n6171), .A2(n3240), .B1(n3241), .B2(n2686), .C1(n3238), 
        .C2(n6182), .ZN(memWrData[28]) );
  OAI222_X2 U6326 ( .A1(n6154), .A2(n3240), .B1(n3241), .B2(n2673), .C1(n3238), 
        .C2(n6284), .ZN(memWrData[29]) );
  OAI222_X2 U6327 ( .A1(n6160), .A2(n3240), .B1(n3241), .B2(n2783), .C1(n3238), 
        .C2(n6259), .ZN(memWrData[30]) );
  OAI222_X2 U6328 ( .A1(n6146), .A2(n3240), .B1(n3241), .B2(n2845), .C1(n3238), 
        .C2(n6293), .ZN(memWrData[31]) );
  MUX2_X1 U6329 ( .A(reg31Val_3[1]), .B(reg31Val_0[1]), .S(n3297), .Z(n6637)
         );
  MUX2_X1 U6330 ( .A(reg31Val_3[0]), .B(reg31Val_0[0]), .S(n3294), .Z(n6638)
         );
  MUX2_X1 U6331 ( .A(rd_3[4]), .B(rd[4]), .S(n3294), .Z(n6639) );
  MUX2_X1 U6332 ( .A(rd_3[3]), .B(rd[3]), .S(n3294), .Z(n6640) );
  MUX2_X1 U6333 ( .A(rd_3[2]), .B(rd[2]), .S(n3294), .Z(n6641) );
  MUX2_X1 U6334 ( .A(rd_3[1]), .B(rd[1]), .S(n3294), .Z(n6642) );
  MUX2_X1 U6335 ( .A(rd_3[0]), .B(rd[0]), .S(n3294), .Z(n6643) );
  INV_X1 U6336 ( .A(n6342), .ZN(n6645) );
  MUX2_X1 U6337 ( .A(n6291), .B(n6331), .S(n3295), .Z(n6342) );
  INV_X1 U6338 ( .A(n6343), .ZN(n6646) );
  MUX2_X1 U6339 ( .A(n6283), .B(n6323), .S(n3295), .Z(n6343) );
  INV_X1 U6340 ( .A(n6344), .ZN(n6647) );
  MUX2_X1 U6341 ( .A(n6293), .B(n6333), .S(n3295), .Z(n6344) );
  INV_X1 U6342 ( .A(n6345), .ZN(n6648) );
  MUX2_X1 U6343 ( .A(n6259), .B(n6319), .S(n3295), .Z(n6345) );
  INV_X1 U6344 ( .A(n6346), .ZN(n6649) );
  MUX2_X1 U6345 ( .A(n6284), .B(n6324), .S(n3295), .Z(n6346) );
  INV_X1 U6346 ( .A(n6347), .ZN(n6650) );
  MUX2_X1 U6347 ( .A(n6182), .B(n6309), .S(n3295), .Z(n6347) );
  INV_X1 U6348 ( .A(n6348), .ZN(n6651) );
  MUX2_X1 U6349 ( .A(n6181), .B(n6308), .S(n3295), .Z(n6348) );
  INV_X1 U6350 ( .A(n6349), .ZN(n6652) );
  MUX2_X1 U6351 ( .A(n6180), .B(n6307), .S(n3295), .Z(n6349) );
  INV_X1 U6352 ( .A(n6350), .ZN(n6653) );
  MUX2_X1 U6353 ( .A(n6294), .B(n6334), .S(n3295), .Z(n6350) );
  INV_X1 U6354 ( .A(n6351), .ZN(n6654) );
  MUX2_X1 U6355 ( .A(n6295), .B(n6335), .S(n3295), .Z(n6351) );
  INV_X1 U6356 ( .A(n6352), .ZN(n6655) );
  MUX2_X1 U6357 ( .A(n6296), .B(n6336), .S(n3295), .Z(n6352) );
  INV_X1 U6358 ( .A(n6353), .ZN(n6656) );
  MUX2_X1 U6359 ( .A(n6297), .B(n6337), .S(n3295), .Z(n6353) );
  INV_X1 U6360 ( .A(n6354), .ZN(n6657) );
  MUX2_X1 U6361 ( .A(n6298), .B(n6338), .S(n3295), .Z(n6354) );
  INV_X1 U6362 ( .A(n6355), .ZN(n6658) );
  MUX2_X1 U6363 ( .A(n6175), .B(n6304), .S(n3295), .Z(n6355) );
  INV_X1 U6364 ( .A(n6356), .ZN(n6659) );
  MUX2_X1 U6365 ( .A(n6258), .B(n6318), .S(n3295), .Z(n6356) );
  INV_X1 U6366 ( .A(n6357), .ZN(n6660) );
  MUX2_X1 U6367 ( .A(n6173), .B(n6302), .S(n3295), .Z(n6357) );
  INV_X1 U6368 ( .A(n6358), .ZN(n6661) );
  MUX2_X1 U6369 ( .A(n6172), .B(n6301), .S(n3295), .Z(n6358) );
  INV_X1 U6370 ( .A(n6359), .ZN(n6662) );
  MUX2_X1 U6371 ( .A(n6299), .B(n6339), .S(n3295), .Z(n6359) );
  INV_X1 U6372 ( .A(n6360), .ZN(n6663) );
  MUX2_X1 U6373 ( .A(n6174), .B(n6303), .S(n3296), .Z(n6360) );
  INV_X1 U6374 ( .A(n6361), .ZN(n6664) );
  MUX2_X1 U6375 ( .A(n6176), .B(n6305), .S(n3296), .Z(n6361) );
  INV_X1 U6376 ( .A(n6362), .ZN(n6665) );
  MUX2_X1 U6377 ( .A(n6281), .B(n6321), .S(n3296), .Z(n6362) );
  INV_X1 U6378 ( .A(n6363), .ZN(n6666) );
  MUX2_X1 U6379 ( .A(n6282), .B(n6322), .S(n3296), .Z(n6363) );
  INV_X1 U6380 ( .A(n6364), .ZN(n6667) );
  MUX2_X1 U6381 ( .A(n6286), .B(n6326), .S(n3296), .Z(n6364) );
  INV_X1 U6382 ( .A(n6365), .ZN(n6668) );
  MUX2_X1 U6383 ( .A(n6280), .B(n6320), .S(n3296), .Z(n6365) );
  INV_X1 U6384 ( .A(n6565), .ZN(n6366) );
  INV_X1 U6385 ( .A(n6566), .ZN(n6367) );
  MUX2_X1 U6386 ( .A(memRdData[0]), .B(\wb/dsize_reg/z2 [0]), .S(n3296), .Z(
        n2267) );
  MUX2_X1 U6387 ( .A(memRdData[1]), .B(\wb/dsize_reg/z2 [1]), .S(n3296), .Z(
        n2266) );
  MUX2_X1 U6388 ( .A(memRdData[2]), .B(\wb/dsize_reg/z2 [2]), .S(n3296), .Z(
        n2265) );
  MUX2_X1 U6389 ( .A(memRdData[3]), .B(\wb/dsize_reg/z2 [3]), .S(n3296), .Z(
        n2264) );
  MUX2_X1 U6390 ( .A(memRdData[4]), .B(\wb/dsize_reg/z2 [4]), .S(n3296), .Z(
        n2263) );
  MUX2_X1 U6391 ( .A(memRdData[5]), .B(\wb/dsize_reg/z2 [5]), .S(n3296), .Z(
        n2262) );
  MUX2_X1 U6392 ( .A(memRdData[6]), .B(\wb/dsize_reg/z2 [6]), .S(n3296), .Z(
        n2261) );
  MUX2_X1 U6393 ( .A(memRdData[7]), .B(\wb/dsize_reg/z2 [7]), .S(n3296), .Z(
        n2260) );
  MUX2_X1 U6394 ( .A(memRdData[8]), .B(\wb/dsize_reg/z2 [8]), .S(n3296), .Z(
        n2259) );
  MUX2_X1 U6395 ( .A(memRdData[9]), .B(\wb/dsize_reg/z2 [9]), .S(n3296), .Z(
        n2258) );
  MUX2_X1 U6396 ( .A(memRdData[10]), .B(\wb/dsize_reg/z2 [10]), .S(n3296), .Z(
        n2257) );
  MUX2_X1 U6397 ( .A(memRdData[11]), .B(\wb/dsize_reg/z2 [11]), .S(n3296), .Z(
        n2256) );
  MUX2_X1 U6398 ( .A(memRdData[12]), .B(\wb/dsize_reg/z2 [12]), .S(n3297), .Z(
        n2255) );
  MUX2_X1 U6399 ( .A(memRdData[13]), .B(\wb/dsize_reg/z2 [13]), .S(n3297), .Z(
        n2254) );
  MUX2_X1 U6400 ( .A(memRdData[14]), .B(\wb/dsize_reg/z2 [14]), .S(n3297), .Z(
        n2253) );
  MUX2_X1 U6401 ( .A(memRdData[15]), .B(\wb/dsize_reg/z2 [15]), .S(n3297), .Z(
        n2252) );
  MUX2_X1 U6402 ( .A(memRdData[16]), .B(\wb/dsize_reg/z2 [16]), .S(n3297), .Z(
        n2251) );
  MUX2_X1 U6403 ( .A(memRdData[17]), .B(\wb/dsize_reg/z2 [17]), .S(n3297), .Z(
        n2250) );
  MUX2_X1 U6404 ( .A(memRdData[18]), .B(\wb/dsize_reg/z2 [18]), .S(n3297), .Z(
        n2249) );
  MUX2_X1 U6405 ( .A(memRdData[19]), .B(\wb/dsize_reg/z2 [19]), .S(n3297), .Z(
        n2248) );
  MUX2_X1 U6406 ( .A(memRdData[20]), .B(\wb/dsize_reg/z2 [20]), .S(n3297), .Z(
        n2247) );
  MUX2_X1 U6407 ( .A(memRdData[21]), .B(\wb/dsize_reg/z2 [21]), .S(n3297), .Z(
        n2246) );
  MUX2_X1 U6408 ( .A(memRdData[22]), .B(\wb/dsize_reg/z2 [22]), .S(n3297), .Z(
        n2245) );
  MUX2_X1 U6409 ( .A(memRdData[23]), .B(\wb/dsize_reg/z2 [23]), .S(n3297), .Z(
        n2244) );
  MUX2_X1 U6410 ( .A(memRdData[24]), .B(\wb/dsize_reg/z2 [24]), .S(n3297), .Z(
        n2243) );
  MUX2_X1 U6411 ( .A(memRdData[25]), .B(\wb/dsize_reg/z2 [25]), .S(n3297), .Z(
        n2242) );
  MUX2_X1 U6412 ( .A(memRdData[26]), .B(\wb/dsize_reg/z2 [26]), .S(n3297), .Z(
        n2241) );
  MUX2_X1 U6413 ( .A(memRdData[27]), .B(\wb/dsize_reg/z2 [27]), .S(n3297), .Z(
        n2240) );
  MUX2_X1 U6414 ( .A(memRdData[28]), .B(\wb/dsize_reg/z2 [28]), .S(n3297), .Z(
        n2239) );
  MUX2_X1 U6415 ( .A(memRdData[29]), .B(\wb/dsize_reg/z2 [29]), .S(n3298), .Z(
        n2238) );
  MUX2_X1 U6416 ( .A(memRdData[30]), .B(\wb/dsize_reg/z2 [30]), .S(n3298), .Z(
        n2237) );
  MUX2_X1 U6417 ( .A(memRdData[31]), .B(\wb/dsize_reg/z2 [31]), .S(n3298), .Z(
        n2236) );
  INV_X1 U6418 ( .A(n6373), .ZN(n2235) );
  MUX2_X1 U6419 ( .A(n6300), .B(n6340), .S(n3298), .Z(n6373) );
  INV_X1 U6420 ( .A(n6374), .ZN(n2227) );
  MUX2_X1 U6421 ( .A(n6292), .B(n6332), .S(n3298), .Z(n6374) );
  INV_X1 U6422 ( .A(n6375), .ZN(n2225) );
  MUX2_X1 U6423 ( .A(n6290), .B(n6330), .S(n3298), .Z(n6375) );
  INV_X1 U6424 ( .A(n6376), .ZN(n2224) );
  MUX2_X1 U6425 ( .A(n6289), .B(n6329), .S(n3298), .Z(n6376) );
  INV_X1 U6426 ( .A(n6377), .ZN(n2223) );
  MUX2_X1 U6427 ( .A(n6288), .B(n6328), .S(n3298), .Z(n6377) );
  INV_X1 U6428 ( .A(n6378), .ZN(n2222) );
  MUX2_X1 U6429 ( .A(n6287), .B(n6327), .S(n3298), .Z(n6378) );
  INV_X1 U6430 ( .A(n6379), .ZN(n2220) );
  MUX2_X1 U6431 ( .A(n6285), .B(n6325), .S(n3298), .Z(n6379) );
  NOR2_X1 U6432 ( .A1(n6385), .A2(n6386), .ZN(n6384) );
  NAND4_X1 U6433 ( .A1(n6387), .A2(n6388), .A3(n6389), .A4(n6390), .ZN(n2135)
         );
  NAND3_X1 U6434 ( .A1(n6589), .A2(n6392), .A3(n6136), .ZN(n6389) );
  OAI21_X1 U6435 ( .B1(n2597), .B2(n2630), .A(n2603), .ZN(n6392) );
  NAND4_X1 U6436 ( .A1(n6592), .A2(n6393), .A3(n6135), .A4(n2837), .ZN(n6387)
         );
  INV_X1 U6437 ( .A(n6399), .ZN(n6369) );
  INV_X1 U6438 ( .A(n6405), .ZN(n6404) );
  AOI21_X1 U6439 ( .B1(n6394), .B2(n6406), .A(n6315), .ZN(n6405) );
  NAND2_X1 U6440 ( .A1(n6407), .A2(n6587), .ZN(n6403) );
  NAND3_X1 U6441 ( .A1(n6593), .A2(n6317), .A3(n6591), .ZN(n6413) );
  NAND2_X1 U6442 ( .A1(n6419), .A2(n6133), .ZN(n6388) );
  OAI21_X1 U6443 ( .B1(n6420), .B2(n6421), .A(n6382), .ZN(n6415) );
  NAND2_X1 U6444 ( .A1(n6422), .A2(n6132), .ZN(n6382) );
  OAI221_X1 U6445 ( .B1(n2604), .B2(n6425), .C1(n6316), .C2(n6418), .A(n6426), 
        .ZN(n6424) );
  NAND3_X1 U6446 ( .A1(n6427), .A2(n6428), .A3(n6429), .ZN(n2017) );
  OAI33_X1 U6447 ( .A1(n2603), .A2(n6589), .A3(n6433), .B1(n6421), .B2(n2630), 
        .B3(n6397), .ZN(n6432) );
  INV_X1 U6448 ( .A(n6425), .ZN(n6431) );
  NAND3_X1 U6449 ( .A1(n6593), .A2(n6434), .A3(n6386), .ZN(n6425) );
  MUX2_X1 U6450 ( .A(n6435), .B(n6592), .S(n6591), .Z(n6430) );
  NOR2_X1 U6451 ( .A1(n6592), .A2(n6316), .ZN(n6435) );
  INV_X1 U6452 ( .A(n6391), .ZN(n6428) );
  NAND2_X1 U6453 ( .A1(n6423), .A2(n2630), .ZN(n6436) );
  INV_X1 U6454 ( .A(n6420), .ZN(n6423) );
  NAND3_X1 U6455 ( .A1(n6135), .A2(n2636), .A3(n6393), .ZN(n6426) );
  INV_X1 U6456 ( .A(n6437), .ZN(n6393) );
  NAND2_X1 U6457 ( .A1(n6419), .A2(n2837), .ZN(n6438) );
  NOR3_X1 U6458 ( .A1(n6437), .A2(n6316), .A3(n2636), .ZN(n6419) );
  NAND3_X1 U6459 ( .A1(n6439), .A2(n6440), .A3(n6441), .ZN(n2016) );
  AOI211_X1 U6460 ( .C1(n6138), .C2(n6316), .A(n6131), .B(n6442), .ZN(n6441)
         );
  INV_X1 U6461 ( .A(n6371), .ZN(n6442) );
  AOI21_X1 U6462 ( .B1(n6444), .B2(n6587), .A(n6400), .ZN(n6443) );
  AOI21_X1 U6463 ( .B1(n6128), .B2(n6445), .A(n6383), .ZN(n6439) );
  NOR2_X1 U6464 ( .A1(op0_1), .A2(n6397), .ZN(n6446) );
  INV_X1 U6465 ( .A(n6422), .ZN(n6397) );
  NOR2_X1 U6466 ( .A1(n2594), .A2(n6587), .ZN(n6422) );
  NAND4_X1 U6467 ( .A1(n6386), .A2(n6317), .A3(n2649), .A4(n2604), .ZN(n6437)
         );
  MUX2_X1 U6468 ( .A(n2583), .B(reg31Val_0[2]), .S(n3298), .Z(n1979) );
  INV_X1 U6469 ( .A(n6447), .ZN(n1948) );
  MUX2_X1 U6470 ( .A(n6178), .B(n6306), .S(n3298), .Z(n6447) );
  OR2_X1 U6471 ( .A1(n3282), .A2(initPC[30]), .ZN(n1914) );
  NAND2_X1 U6472 ( .A1(initPC[30]), .A2(n3298), .ZN(n1913) );
  OR2_X1 U6473 ( .A1(n3282), .A2(initPC[29]), .ZN(n1912) );
  NAND2_X1 U6474 ( .A1(initPC[29]), .A2(n3298), .ZN(n1911) );
  OR2_X1 U6475 ( .A1(n3282), .A2(initPC[28]), .ZN(n1910) );
  NAND2_X1 U6476 ( .A1(initPC[28]), .A2(n3298), .ZN(n1909) );
  OR2_X1 U6477 ( .A1(n3282), .A2(initPC[27]), .ZN(n1908) );
  NAND2_X1 U6478 ( .A1(initPC[27]), .A2(n3298), .ZN(n1907) );
  OR2_X1 U6479 ( .A1(n3282), .A2(initPC[26]), .ZN(n1906) );
  NAND2_X1 U6480 ( .A1(initPC[26]), .A2(n3298), .ZN(n1905) );
  OR2_X1 U6481 ( .A1(n3283), .A2(initPC[25]), .ZN(n1904) );
  NAND2_X1 U6482 ( .A1(initPC[25]), .A2(n3298), .ZN(n1903) );
  OR2_X1 U6483 ( .A1(n3283), .A2(initPC[24]), .ZN(n1902) );
  NAND2_X1 U6484 ( .A1(initPC[24]), .A2(n3298), .ZN(n1901) );
  OR2_X1 U6485 ( .A1(n3283), .A2(initPC[23]), .ZN(n1900) );
  NAND2_X1 U6486 ( .A1(initPC[23]), .A2(n3298), .ZN(n1899) );
  OR2_X1 U6487 ( .A1(n3283), .A2(initPC[22]), .ZN(n1898) );
  NAND2_X1 U6488 ( .A1(initPC[22]), .A2(n3298), .ZN(n1897) );
  OR2_X1 U6489 ( .A1(n3283), .A2(initPC[21]), .ZN(n1896) );
  NAND2_X1 U6490 ( .A1(initPC[21]), .A2(n3299), .ZN(n1895) );
  OR2_X1 U6491 ( .A1(n3283), .A2(initPC[20]), .ZN(n1894) );
  NAND2_X1 U6492 ( .A1(initPC[20]), .A2(n3299), .ZN(n1893) );
  OR2_X1 U6493 ( .A1(n3283), .A2(initPC[19]), .ZN(n1892) );
  NAND2_X1 U6494 ( .A1(initPC[19]), .A2(n3299), .ZN(n1891) );
  OR2_X1 U6495 ( .A1(n3283), .A2(initPC[18]), .ZN(n1890) );
  NAND2_X1 U6496 ( .A1(initPC[18]), .A2(n3299), .ZN(n1889) );
  OR2_X1 U6497 ( .A1(n3283), .A2(initPC[17]), .ZN(n1888) );
  NAND2_X1 U6498 ( .A1(initPC[17]), .A2(n3299), .ZN(n1887) );
  OR2_X1 U6499 ( .A1(n3283), .A2(initPC[16]), .ZN(n1886) );
  NAND2_X1 U6500 ( .A1(initPC[16]), .A2(n3299), .ZN(n1885) );
  OR2_X1 U6501 ( .A1(n3283), .A2(initPC[15]), .ZN(n1884) );
  NAND2_X1 U6502 ( .A1(initPC[15]), .A2(n3299), .ZN(n1883) );
  OR2_X1 U6503 ( .A1(n3283), .A2(initPC[14]), .ZN(n1882) );
  NAND2_X1 U6504 ( .A1(initPC[14]), .A2(n3299), .ZN(n1881) );
  OR2_X1 U6505 ( .A1(n3283), .A2(initPC[13]), .ZN(n1880) );
  NAND2_X1 U6506 ( .A1(initPC[13]), .A2(n3299), .ZN(n1879) );
  OR2_X1 U6507 ( .A1(n3283), .A2(initPC[11]), .ZN(n1878) );
  NAND2_X1 U6508 ( .A1(initPC[11]), .A2(n3299), .ZN(n1877) );
  OR2_X1 U6509 ( .A1(n3283), .A2(initPC[10]), .ZN(n1876) );
  NAND2_X1 U6510 ( .A1(initPC[10]), .A2(n3299), .ZN(n1875) );
  OR2_X1 U6511 ( .A1(n3283), .A2(initPC[0]), .ZN(n1874) );
  NAND2_X1 U6512 ( .A1(initPC[0]), .A2(n3299), .ZN(n1873) );
  OR2_X1 U6513 ( .A1(n3283), .A2(initPC[1]), .ZN(n1872) );
  NAND2_X1 U6514 ( .A1(initPC[1]), .A2(n3299), .ZN(n1871) );
  OR2_X1 U6515 ( .A1(n3283), .A2(initPC[2]), .ZN(n1870) );
  NAND2_X1 U6516 ( .A1(initPC[2]), .A2(n3299), .ZN(n1869) );
  OR2_X1 U6517 ( .A1(n3283), .A2(initPC[3]), .ZN(n1868) );
  NAND2_X1 U6518 ( .A1(initPC[3]), .A2(n3299), .ZN(n1867) );
  OR2_X1 U6519 ( .A1(n3283), .A2(initPC[4]), .ZN(n1866) );
  NAND2_X1 U6520 ( .A1(initPC[4]), .A2(n3299), .ZN(n1865) );
  OR2_X1 U6521 ( .A1(n3247), .A2(initPC[6]), .ZN(n1864) );
  NAND2_X1 U6522 ( .A1(initPC[6]), .A2(n3299), .ZN(n1863) );
  OR2_X1 U6523 ( .A1(n3246), .A2(initPC[7]), .ZN(n1862) );
  NAND2_X1 U6524 ( .A1(initPC[7]), .A2(n3299), .ZN(n1861) );
  OR2_X1 U6525 ( .A1(n3283), .A2(initPC[8]), .ZN(n1860) );
  NAND2_X1 U6526 ( .A1(initPC[8]), .A2(n3299), .ZN(n1859) );
  OR2_X1 U6527 ( .A1(n3279), .A2(initPC[9]), .ZN(n1858) );
  NAND2_X1 U6528 ( .A1(initPC[9]), .A2(n3299), .ZN(n1857) );
  OR2_X1 U6529 ( .A1(n3283), .A2(initPC[12]), .ZN(n1856) );
  NAND2_X1 U6530 ( .A1(initPC[12]), .A2(n3299), .ZN(n1855) );
  OR2_X1 U6531 ( .A1(n3279), .A2(initPC[5]), .ZN(n1854) );
  NAND2_X1 U6532 ( .A1(initPC[5]), .A2(n3299), .ZN(n1853) );
  OR2_X1 U6533 ( .A1(n3279), .A2(initPC[31]), .ZN(n1852) );
  NAND2_X1 U6534 ( .A1(initPC[31]), .A2(n3299), .ZN(n1851) );
  OAI222_X1 U6535 ( .A1(n6291), .A2(n3238), .B1(n6148), .B2(n3240), .C1(n2898), 
        .C2(n3242), .ZN(memWrData[9]) );
  OAI222_X1 U6536 ( .A1(n6283), .A2(n3237), .B1(n6155), .B2(n3239), .C1(n2702), 
        .C2(n3242), .ZN(memWrData[8]) );
  OAI222_X1 U6537 ( .A1(n6285), .A2(n3238), .B1(n6139), .B2(n3240), .C1(n2704), 
        .C2(n3242), .ZN(memWrData[7]) );
  OAI222_X1 U6538 ( .A1(n6287), .A2(n3237), .B1(n6152), .B2(n3239), .C1(n2693), 
        .C2(n3242), .ZN(memWrData[6]) );
  OAI222_X1 U6539 ( .A1(n6178), .A2(n3238), .B1(n6163), .B2(n3240), .C1(n2694), 
        .C2(n3242), .ZN(memWrData[5]) );
  OAI222_X1 U6540 ( .A1(n6292), .A2(n3237), .B1(n6147), .B2(n3239), .C1(n2705), 
        .C2(n3242), .ZN(memWrData[4]) );
  OAI222_X1 U6541 ( .A1(n6288), .A2(n3238), .B1(n6151), .B2(n3240), .C1(n2992), 
        .C2(n3242), .ZN(memWrData[3]) );
  OAI222_X1 U6542 ( .A1(n6290), .A2(n3238), .B1(n6149), .B2(n3240), .C1(n2830), 
        .C2(n3241), .ZN(memWrData[2]) );
  OAI222_X1 U6543 ( .A1(n6289), .A2(n3238), .B1(n6150), .B2(n3240), .C1(n2828), 
        .C2(n3241), .ZN(memWrData[1]) );
  OAI222_X1 U6544 ( .A1(n6174), .A2(n3238), .B1(n6165), .B2(n3240), .C1(n2893), 
        .C2(n3241), .ZN(memWrData[15]) );
  OAI222_X1 U6545 ( .A1(n6176), .A2(n3238), .B1(n6164), .B2(n3240), .C1(n2892), 
        .C2(n3241), .ZN(memWrData[14]) );
  OAI222_X1 U6546 ( .A1(n6281), .A2(n3238), .B1(n6157), .B2(n3240), .C1(n2829), 
        .C2(n3241), .ZN(memWrData[13]) );
  OAI222_X1 U6547 ( .A1(n6282), .A2(n3238), .B1(n6156), .B2(n3240), .C1(n3086), 
        .C2(n3241), .ZN(memWrData[12]) );
  OAI222_X1 U6548 ( .A1(n6286), .A2(n3238), .B1(n6153), .B2(n3240), .C1(n2827), 
        .C2(n3241), .ZN(memWrData[11]) );
  OAI222_X1 U6549 ( .A1(n6280), .A2(n3238), .B1(n6158), .B2(n3240), .C1(n2959), 
        .C2(n3241), .ZN(memWrData[10]) );
  OAI222_X1 U6550 ( .A1(n6300), .A2(n3237), .B1(n6234), .B2(n3239), .C1(n2695), 
        .C2(n3242), .ZN(memWrData[0]) );
  NAND3_X1 U6551 ( .A1(n2594), .A2(n2597), .A3(n6407), .ZN(n6399) );
  NOR3_X1 U6552 ( .A1(n2630), .A2(n2662), .A3(n6412), .ZN(n6407) );
  AND2_X1 U6553 ( .A1(n6370), .A2(n6450), .ZN(n6406) );
  NAND4_X1 U6554 ( .A1(n6451), .A2(n6452), .A3(n6453), .A4(n6454), .ZN(n6368)
         );
  NOR4_X1 U6555 ( .A1(n6455), .A2(n6456), .A3(n6253), .A4(n2797), .ZN(n6454)
         );
  NAND3_X1 U6556 ( .A1(instr_2[2]), .A2(instr_2[4]), .A3(instr_2[0]), .ZN(
        n6456) );
  NAND4_X1 U6557 ( .A1(n6457), .A2(n6252), .A3(n6236), .A4(n6458), .ZN(n6455)
         );
  NOR2_X1 U6558 ( .A1(instr_2[6]), .A2(instr_2[7]), .ZN(n6458) );
  NOR4_X1 U6559 ( .A1(n6459), .A2(n6460), .A3(instr_2[16]), .A4(instr_2[17]), 
        .ZN(n6453) );
  NAND3_X1 U6560 ( .A1(n6242), .A2(n6241), .A3(n6243), .ZN(n6460) );
  NAND4_X1 U6561 ( .A1(n6240), .A2(n6239), .A3(n6461), .A4(n6238), .ZN(n6459)
         );
  NOR2_X1 U6562 ( .A1(instr_2[8]), .A2(instr_2[9]), .ZN(n6461) );
  NOR4_X1 U6563 ( .A1(n6462), .A2(n6463), .A3(instr_2[26]), .A4(instr_2[27]), 
        .ZN(n6452) );
  NAND3_X1 U6564 ( .A1(n6248), .A2(n6247), .A3(n6249), .ZN(n6463) );
  NAND4_X1 U6565 ( .A1(n6246), .A2(n6245), .A3(n6464), .A4(n6244), .ZN(n6462)
         );
  NOR2_X1 U6566 ( .A1(instr_2[18]), .A2(instr_2[19]), .ZN(n6464) );
  NOR4_X1 U6567 ( .A1(n6465), .A2(n6466), .A3(instr_2[5]), .A4(n6467), .ZN(
        n6451) );
  XNOR2_X1 U6568 ( .A(n2633), .B(rd_2[0]), .ZN(n6467) );
  NAND3_X1 U6569 ( .A1(n6255), .A2(n6250), .A3(n6256), .ZN(n6466) );
  NAND4_X1 U6570 ( .A1(n6468), .A2(n6469), .A3(n6470), .A4(n6471), .ZN(n6465)
         );
  XNOR2_X1 U6571 ( .A(n2785), .B(n2628), .ZN(n6471) );
  XOR2_X1 U6572 ( .A(n2784), .B(rd_2[2]), .Z(n6470) );
  XOR2_X1 U6573 ( .A(n2598), .B(rd_2[3]), .Z(n6469) );
  XNOR2_X1 U6574 ( .A(rd_3[4]), .B(rd_2[4]), .ZN(n6468) );
  NOR4_X1 U6575 ( .A1(n6472), .A2(n3052), .A3(n6473), .A4(n6474), .ZN(
        \id_ex/N41 ) );
  XOR2_X1 U6576 ( .A(n2632), .B(n6411), .Z(n6474) );
  XNOR2_X1 U6577 ( .A(n2784), .B(\hazard_detect/eq_83/A[2] ), .ZN(n6473) );
  NAND4_X1 U6578 ( .A1(n6475), .A2(n6476), .A3(n6477), .A4(n6478), .ZN(n6472)
         );
  XOR2_X1 U6579 ( .A(n2598), .B(\hazard_detect/eq_83/A[3] ), .Z(n6477) );
  XNOR2_X1 U6580 ( .A(rd_3[0]), .B(\hazard_detect/eq_83/A[0] ), .ZN(n6476) );
  XOR2_X1 U6581 ( .A(n2785), .B(\hazard_detect/eq_83/A[1] ), .Z(n6475) );
  NOR4_X1 U6582 ( .A1(n6479), .A2(n6480), .A3(n6481), .A4(n6482), .ZN(
        \id_ex/N39 ) );
  XOR2_X1 U6583 ( .A(rs1[2]), .B(rd_3[2]), .Z(n6482) );
  XOR2_X1 U6584 ( .A(rs1[1]), .B(rd_3[1]), .Z(n6481) );
  MUX2_X1 U6585 ( .A(n3043), .B(n6483), .S(rd_3[3]), .Z(n6480) );
  NAND4_X1 U6586 ( .A1(n6484), .A2(n6485), .A3(n6457), .A4(n6486), .ZN(n6479)
         );
  INV_X1 U6587 ( .A(n6487), .ZN(n6457) );
  OAI21_X1 U6588 ( .B1(n6488), .B2(n6489), .A(valid_3), .ZN(n6487) );
  NAND2_X1 U6589 ( .A1(n2633), .A2(n2785), .ZN(n6489) );
  NAND3_X1 U6590 ( .A1(n2598), .A2(n2632), .A3(n2784), .ZN(n6488) );
  XOR2_X1 U6591 ( .A(n2633), .B(rs1[0]), .Z(n6485) );
  XOR2_X1 U6592 ( .A(n2632), .B(rs1[4]), .Z(n6484) );
  NOR2_X1 U6593 ( .A1(n6394), .A2(n2597), .ZN(n6386) );
  NAND2_X1 U6594 ( .A1(n6445), .A2(n6588), .ZN(n6394) );
  NAND2_X1 U6595 ( .A1(n6395), .A2(n6449), .ZN(n6450) );
  AOI221_X1 U6596 ( .B1(n6587), .B2(n6444), .C1(n2662), .C2(n6594), .A(n6445), 
        .ZN(n6449) );
  NOR3_X1 U6597 ( .A1(n2650), .A2(n2780), .A3(n2594), .ZN(n6445) );
  INV_X1 U6598 ( .A(n6400), .ZN(n6395) );
  INV_X1 U6599 ( .A(n6385), .ZN(n6370) );
  NAND4_X1 U6600 ( .A1(op0_1), .A2(n6588), .A3(n6494), .A4(n6590), .ZN(n6493)
         );
  NOR2_X1 U6601 ( .A1(n6594), .A2(n2597), .ZN(n6494) );
  INV_X1 U6602 ( .A(n6398), .ZN(\id_ex/N36 ) );
  INV_X1 U6603 ( .A(n6412), .ZN(n6444) );
  NAND2_X1 U6604 ( .A1(n6594), .A2(n2780), .ZN(n6412) );
  XNOR2_X1 U6605 ( .A(rd_2[4]), .B(n6411), .ZN(n6502) );
  XNOR2_X1 U6606 ( .A(rd_2[0]), .B(n6381), .ZN(n6500) );
  XOR2_X1 U6607 ( .A(n2629), .B(\hazard_detect/eq_83/A[2] ), .Z(n6497) );
  XNOR2_X1 U6608 ( .A(rd_2[3]), .B(\hazard_detect/eq_83/A[3] ), .ZN(n6496) );
  NAND4_X1 U6609 ( .A1(n6503), .A2(n6504), .A3(n6505), .A4(n6506), .ZN(n6486)
         );
  NOR4_X1 U6610 ( .A1(n6499), .A2(n2786), .A3(n6507), .A4(n6508), .ZN(n6506)
         );
  XNOR2_X1 U6611 ( .A(rs1[1]), .B(n2628), .ZN(n6508) );
  XNOR2_X1 U6612 ( .A(rs1[0]), .B(n2781), .ZN(n6507) );
  AND4_X1 U6613 ( .A1(n2593), .A2(n2782), .A3(n2629), .A4(n6509), .ZN(n6499)
         );
  NOR2_X1 U6614 ( .A1(rd_2[1]), .A2(rd_2[0]), .ZN(n6509) );
  XNOR2_X1 U6615 ( .A(n2709), .B(n2593), .ZN(n6505) );
  XNOR2_X1 U6616 ( .A(rs1[4]), .B(rd_2[4]), .ZN(n6504) );
  XNOR2_X1 U6617 ( .A(rs1[2]), .B(rd_2[2]), .ZN(n6503) );
  INV_X1 U6618 ( .A(n6410), .ZN(\hazard_detect/eq_83/A[3] ) );
  NOR2_X1 U6619 ( .A1(n2972), .A2(n6396), .ZN(n6410) );
  INV_X1 U6620 ( .A(n6409), .ZN(\hazard_detect/eq_83/A[2] ) );
  NOR2_X1 U6621 ( .A1(n2973), .A2(n6396), .ZN(n6409) );
  INV_X1 U6622 ( .A(n2579), .ZN(\hazard_detect/eq_83/A[1] ) );
  NOR2_X1 U6623 ( .A1(n2974), .A2(n6396), .ZN(n6408) );
  INV_X1 U6624 ( .A(n6381), .ZN(\hazard_detect/eq_83/A[0] ) );
endmodule

