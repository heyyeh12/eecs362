
// NOT GATE



module not_gate (a, z);

// Ports

input a;
output z;

// Implementation

    begin
        assign z = ~a;
    end
endmodule
