
module ex_mem ( clk, rst, ctrl, valid_d, instr_d, incPC_d, busA_d, busB_d, 
        imm32_d, busFP_d, aluRes_d, regDst_d, memRd_d, memWr_d, regWr_d, 
        branch_d, jr_d, jump_d, link_d, op0_d, fp_d, dSize_d, rd_d, 
        memWrData_sel_d, isZero_d, not_trap_d, instr_q, incPC_q, busA_q, 
        busB_q, imm32_q, busFP_q, aluRes_q, regDst_q, memRd_q, memWr_q, 
        regWr_q, branch_q, jr_q, jump_q, link_q, op0_q, fp_q, dSize_q, rd_q, 
        memWrData_sel_q, valid_q, isZero_q, not_trap_q );
  input [1:0] ctrl;
  input [31:0] instr_d;
  input [31:0] incPC_d;
  input [31:0] busA_d;
  input [31:0] busB_d;
  input [31:0] imm32_d;
  input [31:0] busFP_d;
  input [31:0] aluRes_d;
  input [1:0] dSize_d;
  input [4:0] rd_d;
  input [1:0] memWrData_sel_d;
  output [31:0] instr_q;
  output [31:0] incPC_q;
  output [31:0] busA_q;
  output [31:0] busB_q;
  output [31:0] imm32_q;
  output [31:0] busFP_q;
  output [31:0] aluRes_q;
  output [1:0] dSize_q;
  output [4:0] rd_q;
  output [1:0] memWrData_sel_q;
  input clk, rst, valid_d, regDst_d, memRd_d, memWr_d, regWr_d, branch_d, jr_d,
         jump_d, link_d, op0_d, fp_d, isZero_d, not_trap_d;
  output regDst_q, memRd_q, memWr_q, regWr_q, branch_q, jr_q, jump_q, link_q,
         op0_q, fp_q, valid_q, isZero_q, not_trap_q;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561;

  DFFR_X1 valid_q_reg ( .D(n499), .CK(clk), .RN(n560), .Q(valid_q) );
  DFFS_X1 not_trap_q_reg ( .D(n498), .CK(clk), .SN(n561), .Q(not_trap_q) );
  DFFR_X1 rd_q_reg_4_ ( .D(n497), .CK(clk), .RN(n559), .Q(rd_q[4]) );
  DFFR_X1 rd_q_reg_3_ ( .D(n496), .CK(clk), .RN(n554), .Q(rd_q[3]) );
  DFFR_X1 rd_q_reg_2_ ( .D(n495), .CK(clk), .RN(n559), .Q(rd_q[2]) );
  DFFR_X1 rd_q_reg_1_ ( .D(n494), .CK(clk), .RN(n553), .Q(rd_q[1]) );
  DFFR_X1 rd_q_reg_0_ ( .D(n493), .CK(clk), .RN(n558), .Q(rd_q[0]) );
  DFF_X1 dSize_q_reg_1_ ( .D(n492), .CK(clk), .Q(dSize_q[1]) );
  DFF_X1 dSize_q_reg_0_ ( .D(n491), .CK(clk), .Q(dSize_q[0]) );
  DFFR_X1 instr_q_reg_31_ ( .D(n490), .CK(clk), .RN(n557), .Q(instr_q[31]) );
  DFFR_X1 instr_q_reg_30_ ( .D(n489), .CK(clk), .RN(n555), .Q(instr_q[30]) );
  DFFR_X1 instr_q_reg_29_ ( .D(n488), .CK(clk), .RN(n558), .Q(instr_q[29]) );
  DFFR_X1 instr_q_reg_28_ ( .D(n487), .CK(clk), .RN(n553), .Q(instr_q[28]) );
  DFFR_X1 instr_q_reg_27_ ( .D(n486), .CK(clk), .RN(n559), .Q(instr_q[27]) );
  DFFR_X1 instr_q_reg_26_ ( .D(n485), .CK(clk), .RN(n553), .Q(instr_q[26]) );
  DFFR_X1 instr_q_reg_25_ ( .D(n484), .CK(clk), .RN(n560), .Q(instr_q[25]) );
  DFFR_X1 instr_q_reg_24_ ( .D(n483), .CK(clk), .RN(n553), .Q(instr_q[24]) );
  DFFR_X1 instr_q_reg_23_ ( .D(n482), .CK(clk), .RN(n556), .Q(instr_q[23]) );
  DFFR_X1 instr_q_reg_22_ ( .D(n481), .CK(clk), .RN(n553), .Q(instr_q[22]) );
  DFFR_X1 instr_q_reg_21_ ( .D(n480), .CK(clk), .RN(n553), .Q(instr_q[21]) );
  DFFR_X1 instr_q_reg_20_ ( .D(n479), .CK(clk), .RN(n553), .Q(instr_q[20]) );
  DFFR_X1 instr_q_reg_19_ ( .D(n478), .CK(clk), .RN(n553), .Q(instr_q[19]) );
  DFFR_X1 instr_q_reg_18_ ( .D(n477), .CK(clk), .RN(n552), .Q(instr_q[18]) );
  DFFR_X1 instr_q_reg_17_ ( .D(n476), .CK(clk), .RN(n553), .Q(instr_q[17]) );
  DFFR_X1 instr_q_reg_16_ ( .D(n475), .CK(clk), .RN(n551), .Q(instr_q[16]) );
  DFFR_X1 instr_q_reg_15_ ( .D(n474), .CK(clk), .RN(n553), .Q(instr_q[15]) );
  DFFR_X1 instr_q_reg_14_ ( .D(n473), .CK(clk), .RN(n550), .Q(instr_q[14]) );
  DFFR_X1 instr_q_reg_13_ ( .D(n472), .CK(clk), .RN(n553), .Q(instr_q[13]) );
  DFFR_X1 instr_q_reg_12_ ( .D(n471), .CK(clk), .RN(n549), .Q(instr_q[12]) );
  DFFR_X1 instr_q_reg_11_ ( .D(n470), .CK(clk), .RN(n553), .Q(instr_q[11]) );
  DFFR_X1 instr_q_reg_10_ ( .D(n469), .CK(clk), .RN(n548), .Q(instr_q[10]) );
  DFFR_X1 instr_q_reg_9_ ( .D(n468), .CK(clk), .RN(n552), .Q(instr_q[9]) );
  DFFR_X1 instr_q_reg_8_ ( .D(n467), .CK(clk), .RN(n555), .Q(instr_q[8]) );
  DFFR_X1 instr_q_reg_7_ ( .D(n466), .CK(clk), .RN(n551), .Q(instr_q[7]) );
  DFFR_X1 instr_q_reg_6_ ( .D(n465), .CK(clk), .RN(n556), .Q(instr_q[6]) );
  DFFR_X1 instr_q_reg_5_ ( .D(n464), .CK(clk), .RN(n550), .Q(instr_q[5]) );
  DFFS_X1 instr_q_reg_4_ ( .D(n463), .CK(clk), .SN(n561), .Q(instr_q[4]) );
  DFFR_X1 instr_q_reg_3_ ( .D(n462), .CK(clk), .RN(n549), .Q(instr_q[3]) );
  DFFS_X1 instr_q_reg_2_ ( .D(n461), .CK(clk), .SN(n561), .Q(instr_q[2]) );
  DFFR_X1 instr_q_reg_1_ ( .D(n460), .CK(clk), .RN(n547), .Q(instr_q[1]) );
  DFFS_X1 instr_q_reg_0_ ( .D(n459), .CK(clk), .SN(n561), .Q(instr_q[0]) );
  DFFR_X1 incPC_q_reg_31_ ( .D(n458), .CK(clk), .RN(n554), .Q(incPC_q[31]) );
  DFFR_X1 incPC_q_reg_30_ ( .D(n457), .CK(clk), .RN(n552), .Q(incPC_q[30]) );
  DFFR_X1 incPC_q_reg_29_ ( .D(n456), .CK(clk), .RN(n552), .Q(incPC_q[29]) );
  DFFR_X1 incPC_q_reg_28_ ( .D(n455), .CK(clk), .RN(n554), .Q(incPC_q[28]) );
  DFFR_X1 incPC_q_reg_27_ ( .D(n454), .CK(clk), .RN(n552), .Q(incPC_q[27]) );
  DFFR_X1 incPC_q_reg_26_ ( .D(n453), .CK(clk), .RN(n554), .Q(incPC_q[26]) );
  DFFR_X1 incPC_q_reg_25_ ( .D(n452), .CK(clk), .RN(n552), .Q(incPC_q[25]) );
  DFFR_X1 incPC_q_reg_24_ ( .D(n451), .CK(clk), .RN(n554), .Q(incPC_q[24]) );
  DFFR_X1 incPC_q_reg_23_ ( .D(n450), .CK(clk), .RN(n552), .Q(incPC_q[23]) );
  DFFR_X1 incPC_q_reg_22_ ( .D(n449), .CK(clk), .RN(n554), .Q(incPC_q[22]) );
  DFFR_X1 incPC_q_reg_21_ ( .D(n448), .CK(clk), .RN(n552), .Q(incPC_q[21]) );
  DFFR_X1 incPC_q_reg_20_ ( .D(n447), .CK(clk), .RN(n554), .Q(incPC_q[20]) );
  DFFR_X1 incPC_q_reg_19_ ( .D(n446), .CK(clk), .RN(n554), .Q(incPC_q[19]) );
  DFFR_X1 incPC_q_reg_18_ ( .D(n445), .CK(clk), .RN(n552), .Q(incPC_q[18]) );
  DFFR_X1 incPC_q_reg_17_ ( .D(n444), .CK(clk), .RN(n554), .Q(incPC_q[17]) );
  DFFR_X1 incPC_q_reg_16_ ( .D(n443), .CK(clk), .RN(n552), .Q(incPC_q[16]) );
  DFFR_X1 incPC_q_reg_15_ ( .D(n442), .CK(clk), .RN(n554), .Q(incPC_q[15]) );
  DFFR_X1 incPC_q_reg_14_ ( .D(n441), .CK(clk), .RN(n551), .Q(incPC_q[14]) );
  DFFR_X1 incPC_q_reg_13_ ( .D(n440), .CK(clk), .RN(n554), .Q(incPC_q[13]) );
  DFFR_X1 incPC_q_reg_12_ ( .D(n439), .CK(clk), .RN(n550), .Q(incPC_q[12]) );
  DFFR_X1 incPC_q_reg_11_ ( .D(n438), .CK(clk), .RN(n555), .Q(incPC_q[11]) );
  DFFR_X1 incPC_q_reg_10_ ( .D(n437), .CK(clk), .RN(n549), .Q(incPC_q[10]) );
  DFFR_X1 incPC_q_reg_9_ ( .D(n436), .CK(clk), .RN(n546), .Q(incPC_q[9]) );
  DFFR_X1 incPC_q_reg_8_ ( .D(n435), .CK(clk), .RN(n553), .Q(incPC_q[8]) );
  DFFR_X1 incPC_q_reg_7_ ( .D(n434), .CK(clk), .RN(n552), .Q(incPC_q[7]) );
  DFFR_X1 incPC_q_reg_6_ ( .D(n433), .CK(clk), .RN(n553), .Q(incPC_q[6]) );
  DFFR_X1 incPC_q_reg_5_ ( .D(n432), .CK(clk), .RN(n552), .Q(incPC_q[5]) );
  DFFR_X1 incPC_q_reg_4_ ( .D(n431), .CK(clk), .RN(n554), .Q(incPC_q[4]) );
  DFFR_X1 incPC_q_reg_3_ ( .D(n430), .CK(clk), .RN(n552), .Q(incPC_q[3]) );
  DFFR_X1 incPC_q_reg_2_ ( .D(n429), .CK(clk), .RN(n554), .Q(incPC_q[2]) );
  DFFR_X1 incPC_q_reg_1_ ( .D(n428), .CK(clk), .RN(n552), .Q(incPC_q[1]) );
  DFFR_X1 incPC_q_reg_0_ ( .D(n427), .CK(clk), .RN(n555), .Q(incPC_q[0]) );
  DFFR_X1 busA_q_reg_31_ ( .D(n426), .CK(clk), .RN(n548), .Q(busA_q[31]) );
  DFFR_X1 busA_q_reg_30_ ( .D(n425), .CK(clk), .RN(n558), .Q(busA_q[30]) );
  DFFR_X1 busA_q_reg_29_ ( .D(n424), .CK(clk), .RN(n558), .Q(busA_q[29]) );
  DFFR_X1 busA_q_reg_28_ ( .D(n423), .CK(clk), .RN(n548), .Q(busA_q[28]) );
  DFFR_X1 busA_q_reg_27_ ( .D(n422), .CK(clk), .RN(n558), .Q(busA_q[27]) );
  DFFR_X1 busA_q_reg_26_ ( .D(n421), .CK(clk), .RN(n548), .Q(busA_q[26]) );
  DFFR_X1 busA_q_reg_25_ ( .D(n420), .CK(clk), .RN(n558), .Q(busA_q[25]) );
  DFFR_X1 busA_q_reg_24_ ( .D(n419), .CK(clk), .RN(n548), .Q(busA_q[24]) );
  DFFR_X1 busA_q_reg_23_ ( .D(n418), .CK(clk), .RN(n559), .Q(busA_q[23]) );
  DFFR_X1 busA_q_reg_22_ ( .D(n417), .CK(clk), .RN(n547), .Q(busA_q[22]) );
  DFFR_X1 busA_q_reg_21_ ( .D(n416), .CK(clk), .RN(n559), .Q(busA_q[21]) );
  DFFR_X1 busA_q_reg_20_ ( .D(n415), .CK(clk), .RN(n547), .Q(busA_q[20]) );
  DFFR_X1 busA_q_reg_19_ ( .D(n414), .CK(clk), .RN(n547), .Q(busA_q[19]) );
  DFFR_X1 busA_q_reg_18_ ( .D(n413), .CK(clk), .RN(n559), .Q(busA_q[18]) );
  DFFR_X1 busA_q_reg_17_ ( .D(n412), .CK(clk), .RN(n547), .Q(busA_q[17]) );
  DFFR_X1 busA_q_reg_16_ ( .D(n411), .CK(clk), .RN(n558), .Q(busA_q[16]) );
  DFFR_X1 busA_q_reg_15_ ( .D(n410), .CK(clk), .RN(n547), .Q(busA_q[15]) );
  DFFR_X1 busA_q_reg_14_ ( .D(n409), .CK(clk), .RN(n559), .Q(busA_q[14]) );
  DFFR_X1 busA_q_reg_13_ ( .D(n408), .CK(clk), .RN(n547), .Q(busA_q[13]) );
  DFFR_X1 busA_q_reg_12_ ( .D(n407), .CK(clk), .RN(n559), .Q(busA_q[12]) );
  DFFR_X1 busA_q_reg_11_ ( .D(n406), .CK(clk), .RN(n547), .Q(busA_q[11]) );
  DFFR_X1 busA_q_reg_10_ ( .D(n405), .CK(clk), .RN(n559), .Q(busA_q[10]) );
  DFFR_X1 busA_q_reg_9_ ( .D(n404), .CK(clk), .RN(n557), .Q(busA_q[9]) );
  DFFR_X1 busA_q_reg_8_ ( .D(n403), .CK(clk), .RN(n548), .Q(busA_q[8]) );
  DFFR_X1 busA_q_reg_7_ ( .D(n402), .CK(clk), .RN(n558), .Q(busA_q[7]) );
  DFFR_X1 busA_q_reg_6_ ( .D(n401), .CK(clk), .RN(n548), .Q(busA_q[6]) );
  DFFR_X1 busA_q_reg_5_ ( .D(n400), .CK(clk), .RN(n558), .Q(busA_q[5]) );
  DFFR_X1 busA_q_reg_4_ ( .D(n399), .CK(clk), .RN(n548), .Q(busA_q[4]) );
  DFFR_X1 busA_q_reg_3_ ( .D(n398), .CK(clk), .RN(n558), .Q(busA_q[3]) );
  DFFR_X1 busA_q_reg_2_ ( .D(n397), .CK(clk), .RN(n548), .Q(busA_q[2]) );
  DFFR_X1 busA_q_reg_1_ ( .D(n396), .CK(clk), .RN(n559), .Q(busA_q[1]) );
  DFFR_X1 busA_q_reg_0_ ( .D(n395), .CK(clk), .RN(n547), .Q(busA_q[0]) );
  DFFR_X1 busB_q_reg_31_ ( .D(n394), .CK(clk), .RN(n549), .Q(busB_q[31]) );
  DFFR_X1 busB_q_reg_30_ ( .D(n393), .CK(clk), .RN(n560), .Q(busB_q[30]) );
  DFFR_X1 busB_q_reg_29_ ( .D(n392), .CK(clk), .RN(n557), .Q(busB_q[29]) );
  DFFR_X1 busB_q_reg_28_ ( .D(n391), .CK(clk), .RN(n549), .Q(busB_q[28]) );
  DFFR_X1 busB_q_reg_27_ ( .D(n390), .CK(clk), .RN(n557), .Q(busB_q[27]) );
  DFFR_X1 busB_q_reg_26_ ( .D(n389), .CK(clk), .RN(n549), .Q(busB_q[26]) );
  DFFR_X1 busB_q_reg_25_ ( .D(n388), .CK(clk), .RN(n557), .Q(busB_q[25]) );
  DFFR_X1 busB_q_reg_24_ ( .D(n387), .CK(clk), .RN(n549), .Q(busB_q[24]) );
  DFFR_X1 busB_q_reg_23_ ( .D(n386), .CK(clk), .RN(n557), .Q(busB_q[23]) );
  DFFR_X1 busB_q_reg_22_ ( .D(n385), .CK(clk), .RN(n549), .Q(busB_q[22]) );
  DFFR_X1 busB_q_reg_21_ ( .D(n384), .CK(clk), .RN(n557), .Q(busB_q[21]) );
  DFFR_X1 busB_q_reg_20_ ( .D(n383), .CK(clk), .RN(n549), .Q(busB_q[20]) );
  DFFR_X1 busB_q_reg_19_ ( .D(n382), .CK(clk), .RN(n549), .Q(busB_q[19]) );
  DFFR_X1 busB_q_reg_18_ ( .D(n381), .CK(clk), .RN(n557), .Q(busB_q[18]) );
  DFFR_X1 busB_q_reg_17_ ( .D(n380), .CK(clk), .RN(n549), .Q(busB_q[17]) );
  DFFR_X1 busB_q_reg_16_ ( .D(n379), .CK(clk), .RN(n558), .Q(busB_q[16]) );
  DFFR_X1 busB_q_reg_15_ ( .D(n378), .CK(clk), .RN(n548), .Q(busB_q[15]) );
  DFFR_X1 busB_q_reg_14_ ( .D(n377), .CK(clk), .RN(n558), .Q(busB_q[14]) );
  DFFR_X1 busB_q_reg_13_ ( .D(n376), .CK(clk), .RN(n548), .Q(busB_q[13]) );
  DFFR_X1 busB_q_reg_12_ ( .D(n375), .CK(clk), .RN(n558), .Q(busB_q[12]) );
  DFFR_X1 busB_q_reg_11_ ( .D(n374), .CK(clk), .RN(n548), .Q(busB_q[11]) );
  DFFR_X1 busB_q_reg_10_ ( .D(n373), .CK(clk), .RN(n558), .Q(busB_q[10]) );
  DFFR_X1 busB_q_reg_9_ ( .D(n372), .CK(clk), .RN(n557), .Q(busB_q[9]) );
  DFFR_X1 busB_q_reg_8_ ( .D(n371), .CK(clk), .RN(n549), .Q(busB_q[8]) );
  DFFR_X1 busB_q_reg_7_ ( .D(n370), .CK(clk), .RN(n557), .Q(busB_q[7]) );
  DFFR_X1 busB_q_reg_6_ ( .D(n369), .CK(clk), .RN(n549), .Q(busB_q[6]) );
  DFFR_X1 busB_q_reg_5_ ( .D(n368), .CK(clk), .RN(n557), .Q(busB_q[5]) );
  DFFR_X1 busB_q_reg_4_ ( .D(n367), .CK(clk), .RN(n549), .Q(busB_q[4]) );
  DFFR_X1 busB_q_reg_3_ ( .D(n366), .CK(clk), .RN(n557), .Q(busB_q[3]) );
  DFFR_X1 busB_q_reg_2_ ( .D(n365), .CK(clk), .RN(n549), .Q(busB_q[2]) );
  DFFR_X1 busB_q_reg_1_ ( .D(n364), .CK(clk), .RN(n557), .Q(busB_q[1]) );
  DFFR_X1 busB_q_reg_0_ ( .D(n363), .CK(clk), .RN(n548), .Q(busB_q[0]) );
  DFFR_X1 imm32_q_reg_31_ ( .D(n362), .CK(clk), .RN(n555), .Q(imm32_q[31]) );
  DFFR_X1 imm32_q_reg_30_ ( .D(n361), .CK(clk), .RN(n548), .Q(imm32_q[30]) );
  DFFR_X1 imm32_q_reg_29_ ( .D(n360), .CK(clk), .RN(n547), .Q(imm32_q[29]) );
  DFFR_X1 imm32_q_reg_28_ ( .D(n359), .CK(clk), .RN(n555), .Q(imm32_q[28]) );
  DFFR_X1 imm32_q_reg_27_ ( .D(n358), .CK(clk), .RN(n546), .Q(imm32_q[27]) );
  DFFR_X1 imm32_q_reg_26_ ( .D(n357), .CK(clk), .RN(n555), .Q(imm32_q[26]) );
  DFFR_X1 imm32_q_reg_25_ ( .D(n356), .CK(clk), .RN(n557), .Q(imm32_q[25]) );
  DFFR_X1 imm32_q_reg_24_ ( .D(n355), .CK(clk), .RN(n555), .Q(imm32_q[24]) );
  DFFR_X1 imm32_q_reg_23_ ( .D(n354), .CK(clk), .RN(n558), .Q(imm32_q[23]) );
  DFFR_X1 imm32_q_reg_22_ ( .D(n353), .CK(clk), .RN(n555), .Q(imm32_q[22]) );
  DFFR_X1 imm32_q_reg_21_ ( .D(n352), .CK(clk), .RN(n551), .Q(imm32_q[21]) );
  DFFR_X1 imm32_q_reg_20_ ( .D(n351), .CK(clk), .RN(n555), .Q(imm32_q[20]) );
  DFFR_X1 imm32_q_reg_19_ ( .D(n350), .CK(clk), .RN(n556), .Q(imm32_q[19]) );
  DFFR_X1 imm32_q_reg_18_ ( .D(n349), .CK(clk), .RN(n551), .Q(imm32_q[18]) );
  DFFR_X1 imm32_q_reg_17_ ( .D(n348), .CK(clk), .RN(n556), .Q(imm32_q[17]) );
  DFFR_X1 imm32_q_reg_16_ ( .D(n347), .CK(clk), .RN(n551), .Q(imm32_q[16]) );
  DFFR_X1 imm32_q_reg_15_ ( .D(n346), .CK(clk), .RN(n556), .Q(imm32_q[15]) );
  DFFR_X1 imm32_q_reg_14_ ( .D(n345), .CK(clk), .RN(n551), .Q(imm32_q[14]) );
  DFFR_X1 imm32_q_reg_13_ ( .D(n344), .CK(clk), .RN(n556), .Q(imm32_q[13]) );
  DFFR_X1 imm32_q_reg_12_ ( .D(n343), .CK(clk), .RN(n551), .Q(imm32_q[12]) );
  DFFR_X1 imm32_q_reg_11_ ( .D(n342), .CK(clk), .RN(n556), .Q(imm32_q[11]) );
  DFFR_X1 imm32_q_reg_10_ ( .D(n341), .CK(clk), .RN(n551), .Q(imm32_q[10]) );
  DFFR_X1 imm32_q_reg_9_ ( .D(n340), .CK(clk), .RN(n559), .Q(imm32_q[9]) );
  DFFR_X1 imm32_q_reg_8_ ( .D(n339), .CK(clk), .RN(n555), .Q(imm32_q[8]) );
  DFFR_X1 imm32_q_reg_7_ ( .D(n338), .CK(clk), .RN(n560), .Q(imm32_q[7]) );
  DFFR_X1 imm32_q_reg_6_ ( .D(n337), .CK(clk), .RN(n555), .Q(imm32_q[6]) );
  DFFR_X1 imm32_q_reg_5_ ( .D(n336), .CK(clk), .RN(n554), .Q(imm32_q[5]) );
  DFFR_X1 imm32_q_reg_4_ ( .D(n335), .CK(clk), .RN(n555), .Q(imm32_q[4]) );
  DFFR_X1 imm32_q_reg_3_ ( .D(n334), .CK(clk), .RN(n556), .Q(imm32_q[3]) );
  DFFR_X1 imm32_q_reg_2_ ( .D(n333), .CK(clk), .RN(n555), .Q(imm32_q[2]) );
  DFFR_X1 imm32_q_reg_1_ ( .D(n332), .CK(clk), .RN(n551), .Q(imm32_q[1]) );
  DFFR_X1 imm32_q_reg_0_ ( .D(n331), .CK(clk), .RN(n556), .Q(imm32_q[0]) );
  DFFR_X1 busFP_q_reg_31_ ( .D(n330), .CK(clk), .RN(n551), .Q(busFP_q[31]) );
  DFFR_X1 busFP_q_reg_30_ ( .D(n329), .CK(clk), .RN(n556), .Q(busFP_q[30]) );
  DFFR_X1 busFP_q_reg_29_ ( .D(n328), .CK(clk), .RN(n556), .Q(busFP_q[29]) );
  DFFR_X1 busFP_q_reg_28_ ( .D(n327), .CK(clk), .RN(n550), .Q(busFP_q[28]) );
  DFFR_X1 busFP_q_reg_27_ ( .D(n326), .CK(clk), .RN(n556), .Q(busFP_q[27]) );
  DFFR_X1 busFP_q_reg_26_ ( .D(n325), .CK(clk), .RN(n550), .Q(busFP_q[26]) );
  DFFR_X1 busFP_q_reg_25_ ( .D(n324), .CK(clk), .RN(n553), .Q(busFP_q[25]) );
  DFFR_X1 busFP_q_reg_24_ ( .D(n323), .CK(clk), .RN(n550), .Q(busFP_q[24]) );
  DFFR_X1 busFP_q_reg_23_ ( .D(n322), .CK(clk), .RN(n554), .Q(busFP_q[23]) );
  DFFR_X1 busFP_q_reg_22_ ( .D(n321), .CK(clk), .RN(n550), .Q(busFP_q[22]) );
  DFFR_X1 busFP_q_reg_21_ ( .D(n320), .CK(clk), .RN(n552), .Q(busFP_q[21]) );
  DFFR_X1 busFP_q_reg_20_ ( .D(n319), .CK(clk), .RN(n550), .Q(busFP_q[20]) );
  DFFR_X1 busFP_q_reg_19_ ( .D(n318), .CK(clk), .RN(n550), .Q(busFP_q[19]) );
  DFFR_X1 busFP_q_reg_18_ ( .D(n317), .CK(clk), .RN(n551), .Q(busFP_q[18]) );
  DFFR_X1 busFP_q_reg_17_ ( .D(n316), .CK(clk), .RN(n550), .Q(busFP_q[17]) );
  DFFR_X1 busFP_q_reg_16_ ( .D(n315), .CK(clk), .RN(n550), .Q(busFP_q[16]) );
  DFFR_X1 busFP_q_reg_15_ ( .D(n314), .CK(clk), .RN(n550), .Q(busFP_q[15]) );
  DFFR_X1 busFP_q_reg_14_ ( .D(n313), .CK(clk), .RN(n549), .Q(busFP_q[14]) );
  DFFR_X1 busFP_q_reg_13_ ( .D(n312), .CK(clk), .RN(n550), .Q(busFP_q[13]) );
  DFFR_X1 busFP_q_reg_12_ ( .D(n311), .CK(clk), .RN(n548), .Q(busFP_q[12]) );
  DFFR_X1 busFP_q_reg_11_ ( .D(n310), .CK(clk), .RN(n550), .Q(busFP_q[11]) );
  DFFR_X1 busFP_q_reg_10_ ( .D(n309), .CK(clk), .RN(n547), .Q(busFP_q[10]) );
  DFFR_X1 busFP_q_reg_9_ ( .D(n308), .CK(clk), .RN(n556), .Q(busFP_q[9]) );
  DFFR_X1 busFP_q_reg_8_ ( .D(n307), .CK(clk), .RN(n551), .Q(busFP_q[8]) );
  DFFR_X1 busFP_q_reg_7_ ( .D(n306), .CK(clk), .RN(n556), .Q(busFP_q[7]) );
  DFFR_X1 busFP_q_reg_6_ ( .D(n305), .CK(clk), .RN(n555), .Q(busFP_q[6]) );
  DFFR_X1 busFP_q_reg_5_ ( .D(n304), .CK(clk), .RN(n556), .Q(busFP_q[5]) );
  DFFR_X1 busFP_q_reg_4_ ( .D(n303), .CK(clk), .RN(n551), .Q(busFP_q[4]) );
  DFFR_X1 busFP_q_reg_3_ ( .D(n302), .CK(clk), .RN(n556), .Q(busFP_q[3]) );
  DFFR_X1 busFP_q_reg_2_ ( .D(n301), .CK(clk), .RN(n550), .Q(busFP_q[2]) );
  DFFR_X1 busFP_q_reg_1_ ( .D(n300), .CK(clk), .RN(n546), .Q(busFP_q[1]) );
  DFFR_X1 busFP_q_reg_0_ ( .D(n299), .CK(clk), .RN(n550), .Q(busFP_q[0]) );
  DFFR_X1 aluRes_q_reg_31_ ( .D(n298), .CK(clk), .RN(n560), .Q(aluRes_q[31])
         );
  DFFR_X1 aluRes_q_reg_30_ ( .D(n297), .CK(clk), .RN(n546), .Q(aluRes_q[30])
         );
  DFFR_X1 aluRes_q_reg_29_ ( .D(n296), .CK(clk), .RN(n546), .Q(aluRes_q[29])
         );
  DFFR_X1 aluRes_q_reg_28_ ( .D(n295), .CK(clk), .RN(n560), .Q(aluRes_q[28])
         );
  DFFR_X1 aluRes_q_reg_27_ ( .D(n294), .CK(clk), .RN(n546), .Q(aluRes_q[27])
         );
  DFFR_X1 aluRes_q_reg_26_ ( .D(n293), .CK(clk), .RN(n560), .Q(aluRes_q[26])
         );
  DFFR_X1 aluRes_q_reg_25_ ( .D(n292), .CK(clk), .RN(n546), .Q(aluRes_q[25])
         );
  DFFR_X1 aluRes_q_reg_24_ ( .D(n291), .CK(clk), .RN(n560), .Q(aluRes_q[24])
         );
  DFFR_X1 aluRes_q_reg_23_ ( .D(n290), .CK(clk), .RN(n546), .Q(aluRes_q[23])
         );
  DFFR_X1 aluRes_q_reg_22_ ( .D(n289), .CK(clk), .RN(n560), .Q(aluRes_q[22])
         );
  DFFR_X1 aluRes_q_reg_21_ ( .D(n288), .CK(clk), .RN(n546), .Q(aluRes_q[21])
         );
  DFFR_X1 aluRes_q_reg_20_ ( .D(n287), .CK(clk), .RN(n560), .Q(aluRes_q[20])
         );
  DFFR_X1 aluRes_q_reg_19_ ( .D(n286), .CK(clk), .RN(n560), .Q(aluRes_q[19])
         );
  DFFR_X1 aluRes_q_reg_18_ ( .D(n285), .CK(clk), .RN(n546), .Q(aluRes_q[18])
         );
  DFFR_X1 aluRes_q_reg_17_ ( .D(n284), .CK(clk), .RN(n560), .Q(aluRes_q[17])
         );
  DFFR_X1 aluRes_q_reg_16_ ( .D(n283), .CK(clk), .RN(n546), .Q(aluRes_q[16])
         );
  DFFR_X1 aluRes_q_reg_15_ ( .D(n282), .CK(clk), .RN(n560), .Q(aluRes_q[15])
         );
  DFFR_X1 aluRes_q_reg_14_ ( .D(n281), .CK(clk), .RN(n546), .Q(aluRes_q[14])
         );
  DFFR_X1 aluRes_q_reg_13_ ( .D(n280), .CK(clk), .RN(n560), .Q(aluRes_q[13])
         );
  DFFR_X1 aluRes_q_reg_12_ ( .D(n279), .CK(clk), .RN(n546), .Q(aluRes_q[12])
         );
  DFFR_X1 aluRes_q_reg_11_ ( .D(n278), .CK(clk), .RN(n560), .Q(aluRes_q[11])
         );
  DFFR_X1 aluRes_q_reg_10_ ( .D(n277), .CK(clk), .RN(n551), .Q(aluRes_q[10])
         );
  DFFR_X1 aluRes_q_reg_9_ ( .D(n276), .CK(clk), .RN(n547), .Q(aluRes_q[9]) );
  DFFR_X1 aluRes_q_reg_8_ ( .D(n275), .CK(clk), .RN(n559), .Q(aluRes_q[8]) );
  DFFR_X1 aluRes_q_reg_7_ ( .D(n274), .CK(clk), .RN(n547), .Q(aluRes_q[7]) );
  DFFR_X1 aluRes_q_reg_6_ ( .D(n273), .CK(clk), .RN(n559), .Q(aluRes_q[6]) );
  DFFR_X1 aluRes_q_reg_5_ ( .D(n272), .CK(clk), .RN(n547), .Q(aluRes_q[5]) );
  DFFR_X1 aluRes_q_reg_4_ ( .D(n271), .CK(clk), .RN(n559), .Q(aluRes_q[4]) );
  DFFR_X1 aluRes_q_reg_3_ ( .D(n270), .CK(clk), .RN(n547), .Q(aluRes_q[3]) );
  DFFR_X1 aluRes_q_reg_2_ ( .D(n269), .CK(clk), .RN(n560), .Q(aluRes_q[2]) );
  DFFR_X1 aluRes_q_reg_1_ ( .D(n268), .CK(clk), .RN(n546), .Q(aluRes_q[1]) );
  DFFR_X1 aluRes_q_reg_0_ ( .D(n267), .CK(clk), .RN(n559), .Q(aluRes_q[0]) );
  DFFR_X1 regDst_q_reg ( .D(n266), .CK(clk), .RN(n554), .Q(regDst_q) );
  DFFR_X1 memRd_q_reg ( .D(n265), .CK(clk), .RN(n553), .Q(memRd_q) );
  DFFR_X1 memWr_q_reg ( .D(n264), .CK(clk), .RN(n548), .Q(memWr_q) );
  DFFR_X1 regWr_q_reg ( .D(n263), .CK(clk), .RN(n546), .Q(regWr_q) );
  DFFR_X1 isZero_q_reg ( .D(n262), .CK(clk), .RN(n555), .Q(isZero_q) );
  DFFR_X1 jump_q_reg ( .D(n261), .CK(clk), .RN(n557), .Q(jump_q) );
  DFFR_X1 branch_q_reg ( .D(n260), .CK(clk), .RN(n559), .Q(branch_q) );
  DFFR_X1 jr_q_reg ( .D(n259), .CK(clk), .RN(n547), .Q(jr_q) );
  DFFR_X1 link_q_reg ( .D(n258), .CK(clk), .RN(n546), .Q(link_q) );
  DFFR_X1 op0_q_reg ( .D(n257), .CK(clk), .RN(n557), .Q(op0_q) );
  DFFR_X1 fp_q_reg ( .D(n256), .CK(clk), .RN(n551), .Q(fp_q) );
  DFFR_X1 memWrData_sel_q_reg_1_ ( .D(n255), .CK(clk), .RN(n552), .Q(
        memWrData_sel_q[1]) );
  DFFR_X1 memWrData_sel_q_reg_0_ ( .D(n254), .CK(clk), .RN(n558), .Q(
        memWrData_sel_q[0]) );
  INV_X1 U3 ( .A(n1), .ZN(n499) );
  AOI22_X1 U4 ( .A1(valid_d), .A2(n536), .B1(valid_q), .B2(n512), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n263) );
  AOI22_X1 U6 ( .A1(regWr_d), .A2(n536), .B1(regWr_q), .B2(n512), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n266) );
  AOI22_X1 U8 ( .A1(regDst_d), .A2(n536), .B1(regDst_q), .B2(n512), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n497) );
  AOI22_X1 U10 ( .A1(rd_d[4]), .A2(n535), .B1(rd_q[4]), .B2(n511), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n496) );
  AOI22_X1 U12 ( .A1(rd_d[3]), .A2(n535), .B1(rd_q[3]), .B2(n510), .ZN(n7) );
  INV_X1 U13 ( .A(n8), .ZN(n495) );
  AOI22_X1 U14 ( .A1(rd_d[2]), .A2(n535), .B1(rd_q[2]), .B2(n509), .ZN(n8) );
  INV_X1 U15 ( .A(n9), .ZN(n494) );
  AOI22_X1 U16 ( .A1(rd_d[1]), .A2(n535), .B1(rd_q[1]), .B2(n511), .ZN(n9) );
  INV_X1 U17 ( .A(n10), .ZN(n493) );
  AOI22_X1 U18 ( .A1(rd_d[0]), .A2(n535), .B1(rd_q[0]), .B2(n510), .ZN(n10) );
  INV_X1 U19 ( .A(n11), .ZN(n257) );
  AOI22_X1 U20 ( .A1(op0_d), .A2(n535), .B1(op0_q), .B2(n509), .ZN(n11) );
  INV_X1 U21 ( .A(n12), .ZN(n498) );
  AOI221_X1 U22 ( .B1(not_trap_q), .B2(n503), .C1(not_trap_d), .C2(n526), .A(
        n13), .ZN(n12) );
  INV_X1 U23 ( .A(n14), .ZN(n264) );
  AOI22_X1 U24 ( .A1(memWr_d), .A2(n535), .B1(memWr_q), .B2(n511), .ZN(n14) );
  INV_X1 U25 ( .A(n15), .ZN(n255) );
  AOI22_X1 U26 ( .A1(memWrData_sel_d[1]), .A2(n535), .B1(memWrData_sel_q[1]), 
        .B2(n510), .ZN(n15) );
  INV_X1 U27 ( .A(n16), .ZN(n254) );
  AOI22_X1 U28 ( .A1(memWrData_sel_d[0]), .A2(n535), .B1(memWrData_sel_q[0]), 
        .B2(n509), .ZN(n16) );
  INV_X1 U29 ( .A(n17), .ZN(n265) );
  AOI22_X1 U30 ( .A1(memRd_d), .A2(n535), .B1(memRd_q), .B2(n511), .ZN(n17) );
  INV_X1 U31 ( .A(n18), .ZN(n258) );
  AOI22_X1 U32 ( .A1(link_d), .A2(n535), .B1(link_q), .B2(n510), .ZN(n18) );
  INV_X1 U33 ( .A(n19), .ZN(n261) );
  AOI22_X1 U34 ( .A1(jump_d), .A2(n535), .B1(jump_q), .B2(n509), .ZN(n19) );
  INV_X1 U35 ( .A(n20), .ZN(n259) );
  AOI22_X1 U36 ( .A1(jr_d), .A2(n534), .B1(jr_q), .B2(n511), .ZN(n20) );
  INV_X1 U37 ( .A(n21), .ZN(n262) );
  AOI22_X1 U38 ( .A1(isZero_d), .A2(n534), .B1(isZero_q), .B2(n511), .ZN(n21)
         );
  INV_X1 U39 ( .A(n22), .ZN(n468) );
  AOI22_X1 U40 ( .A1(instr_d[9]), .A2(n534), .B1(instr_q[9]), .B2(n511), .ZN(
        n22) );
  INV_X1 U41 ( .A(n23), .ZN(n467) );
  AOI22_X1 U42 ( .A1(instr_d[8]), .A2(n534), .B1(instr_q[8]), .B2(n511), .ZN(
        n23) );
  INV_X1 U43 ( .A(n24), .ZN(n466) );
  AOI22_X1 U44 ( .A1(instr_d[7]), .A2(n534), .B1(instr_q[7]), .B2(n511), .ZN(
        n24) );
  INV_X1 U45 ( .A(n25), .ZN(n465) );
  AOI22_X1 U46 ( .A1(instr_d[6]), .A2(n534), .B1(instr_q[6]), .B2(n511), .ZN(
        n25) );
  INV_X1 U47 ( .A(n26), .ZN(n464) );
  AOI22_X1 U48 ( .A1(instr_d[5]), .A2(n534), .B1(instr_q[5]), .B2(n511), .ZN(
        n26) );
  INV_X1 U49 ( .A(n27), .ZN(n463) );
  AOI221_X1 U50 ( .B1(instr_q[4]), .B2(n503), .C1(instr_d[4]), .C2(n526), .A(
        n13), .ZN(n27) );
  INV_X1 U51 ( .A(n28), .ZN(n462) );
  AOI22_X1 U52 ( .A1(instr_d[3]), .A2(n534), .B1(instr_q[3]), .B2(n511), .ZN(
        n28) );
  INV_X1 U53 ( .A(n29), .ZN(n490) );
  AOI22_X1 U54 ( .A1(instr_d[31]), .A2(n534), .B1(instr_q[31]), .B2(n511), 
        .ZN(n29) );
  INV_X1 U55 ( .A(n30), .ZN(n489) );
  AOI22_X1 U56 ( .A1(instr_d[30]), .A2(n534), .B1(instr_q[30]), .B2(n511), 
        .ZN(n30) );
  INV_X1 U57 ( .A(n31), .ZN(n461) );
  AOI221_X1 U58 ( .B1(instr_q[2]), .B2(n503), .C1(instr_d[2]), .C2(n526), .A(
        n13), .ZN(n31) );
  INV_X1 U59 ( .A(n32), .ZN(n488) );
  AOI22_X1 U60 ( .A1(instr_d[29]), .A2(n534), .B1(instr_q[29]), .B2(n511), 
        .ZN(n32) );
  INV_X1 U61 ( .A(n33), .ZN(n487) );
  AOI22_X1 U62 ( .A1(instr_d[28]), .A2(n534), .B1(instr_q[28]), .B2(n511), 
        .ZN(n33) );
  INV_X1 U63 ( .A(n34), .ZN(n486) );
  AOI22_X1 U64 ( .A1(instr_d[27]), .A2(n533), .B1(instr_q[27]), .B2(n510), 
        .ZN(n34) );
  INV_X1 U65 ( .A(n35), .ZN(n485) );
  AOI22_X1 U66 ( .A1(instr_d[26]), .A2(n533), .B1(instr_q[26]), .B2(n510), 
        .ZN(n35) );
  INV_X1 U67 ( .A(n36), .ZN(n484) );
  AOI22_X1 U68 ( .A1(instr_d[25]), .A2(n533), .B1(instr_q[25]), .B2(n510), 
        .ZN(n36) );
  INV_X1 U69 ( .A(n37), .ZN(n483) );
  AOI22_X1 U70 ( .A1(instr_d[24]), .A2(n533), .B1(instr_q[24]), .B2(n510), 
        .ZN(n37) );
  INV_X1 U71 ( .A(n38), .ZN(n482) );
  AOI22_X1 U72 ( .A1(instr_d[23]), .A2(n533), .B1(instr_q[23]), .B2(n510), 
        .ZN(n38) );
  INV_X1 U73 ( .A(n39), .ZN(n481) );
  AOI22_X1 U74 ( .A1(instr_d[22]), .A2(n533), .B1(instr_q[22]), .B2(n510), 
        .ZN(n39) );
  INV_X1 U75 ( .A(n40), .ZN(n480) );
  AOI22_X1 U76 ( .A1(instr_d[21]), .A2(n533), .B1(instr_q[21]), .B2(n510), 
        .ZN(n40) );
  INV_X1 U77 ( .A(n41), .ZN(n479) );
  AOI22_X1 U78 ( .A1(instr_d[20]), .A2(n533), .B1(instr_q[20]), .B2(n510), 
        .ZN(n41) );
  INV_X1 U79 ( .A(n42), .ZN(n460) );
  AOI22_X1 U80 ( .A1(instr_d[1]), .A2(n533), .B1(instr_q[1]), .B2(n510), .ZN(
        n42) );
  INV_X1 U81 ( .A(n43), .ZN(n478) );
  AOI22_X1 U82 ( .A1(instr_d[19]), .A2(n533), .B1(instr_q[19]), .B2(n510), 
        .ZN(n43) );
  INV_X1 U83 ( .A(n44), .ZN(n477) );
  AOI22_X1 U84 ( .A1(instr_d[18]), .A2(n533), .B1(instr_q[18]), .B2(n510), 
        .ZN(n44) );
  INV_X1 U85 ( .A(n45), .ZN(n476) );
  AOI22_X1 U86 ( .A1(instr_d[17]), .A2(n533), .B1(instr_q[17]), .B2(n510), 
        .ZN(n45) );
  INV_X1 U87 ( .A(n46), .ZN(n475) );
  AOI22_X1 U88 ( .A1(instr_d[16]), .A2(n532), .B1(instr_q[16]), .B2(n509), 
        .ZN(n46) );
  INV_X1 U89 ( .A(n47), .ZN(n474) );
  AOI22_X1 U90 ( .A1(instr_d[15]), .A2(n532), .B1(instr_q[15]), .B2(n509), 
        .ZN(n47) );
  INV_X1 U91 ( .A(n48), .ZN(n473) );
  AOI22_X1 U92 ( .A1(instr_d[14]), .A2(n532), .B1(instr_q[14]), .B2(n509), 
        .ZN(n48) );
  INV_X1 U93 ( .A(n49), .ZN(n472) );
  AOI22_X1 U94 ( .A1(instr_d[13]), .A2(n532), .B1(instr_q[13]), .B2(n509), 
        .ZN(n49) );
  INV_X1 U95 ( .A(n50), .ZN(n471) );
  AOI22_X1 U96 ( .A1(instr_d[12]), .A2(n532), .B1(instr_q[12]), .B2(n509), 
        .ZN(n50) );
  INV_X1 U97 ( .A(n51), .ZN(n470) );
  AOI22_X1 U98 ( .A1(instr_d[11]), .A2(n532), .B1(instr_q[11]), .B2(n509), 
        .ZN(n51) );
  INV_X1 U99 ( .A(n52), .ZN(n469) );
  AOI22_X1 U100 ( .A1(instr_d[10]), .A2(n532), .B1(instr_q[10]), .B2(n509), 
        .ZN(n52) );
  INV_X1 U101 ( .A(n53), .ZN(n459) );
  AOI221_X1 U102 ( .B1(instr_q[0]), .B2(n503), .C1(instr_d[0]), .C2(n526), .A(
        n13), .ZN(n53) );
  NOR2_X1 U103 ( .A1(n522), .A2(ctrl[0]), .ZN(n13) );
  INV_X1 U104 ( .A(n54), .ZN(n436) );
  AOI22_X1 U105 ( .A1(incPC_d[9]), .A2(n532), .B1(incPC_q[9]), .B2(n509), .ZN(
        n54) );
  INV_X1 U106 ( .A(n55), .ZN(n435) );
  AOI22_X1 U107 ( .A1(incPC_d[8]), .A2(n532), .B1(incPC_q[8]), .B2(n509), .ZN(
        n55) );
  INV_X1 U108 ( .A(n56), .ZN(n434) );
  AOI22_X1 U109 ( .A1(incPC_d[7]), .A2(n532), .B1(incPC_q[7]), .B2(n509), .ZN(
        n56) );
  INV_X1 U110 ( .A(n57), .ZN(n433) );
  AOI22_X1 U111 ( .A1(incPC_d[6]), .A2(n532), .B1(incPC_q[6]), .B2(n509), .ZN(
        n57) );
  INV_X1 U112 ( .A(n58), .ZN(n432) );
  AOI22_X1 U113 ( .A1(incPC_d[5]), .A2(n532), .B1(incPC_q[5]), .B2(n509), .ZN(
        n58) );
  INV_X1 U114 ( .A(n59), .ZN(n431) );
  AOI22_X1 U115 ( .A1(incPC_d[4]), .A2(n531), .B1(incPC_q[4]), .B2(n508), .ZN(
        n59) );
  INV_X1 U116 ( .A(n60), .ZN(n430) );
  AOI22_X1 U117 ( .A1(incPC_d[3]), .A2(n531), .B1(incPC_q[3]), .B2(n508), .ZN(
        n60) );
  INV_X1 U118 ( .A(n61), .ZN(n458) );
  AOI22_X1 U119 ( .A1(incPC_d[31]), .A2(n531), .B1(incPC_q[31]), .B2(n508), 
        .ZN(n61) );
  INV_X1 U120 ( .A(n62), .ZN(n457) );
  AOI22_X1 U121 ( .A1(incPC_d[30]), .A2(n531), .B1(incPC_q[30]), .B2(n508), 
        .ZN(n62) );
  INV_X1 U122 ( .A(n63), .ZN(n429) );
  AOI22_X1 U123 ( .A1(incPC_d[2]), .A2(n531), .B1(incPC_q[2]), .B2(n508), .ZN(
        n63) );
  INV_X1 U124 ( .A(n64), .ZN(n456) );
  AOI22_X1 U125 ( .A1(incPC_d[29]), .A2(n531), .B1(incPC_q[29]), .B2(n508), 
        .ZN(n64) );
  INV_X1 U126 ( .A(n65), .ZN(n455) );
  AOI22_X1 U127 ( .A1(incPC_d[28]), .A2(n531), .B1(incPC_q[28]), .B2(n508), 
        .ZN(n65) );
  INV_X1 U128 ( .A(n66), .ZN(n454) );
  AOI22_X1 U129 ( .A1(incPC_d[27]), .A2(n531), .B1(incPC_q[27]), .B2(n508), 
        .ZN(n66) );
  INV_X1 U130 ( .A(n67), .ZN(n453) );
  AOI22_X1 U131 ( .A1(incPC_d[26]), .A2(n531), .B1(incPC_q[26]), .B2(n508), 
        .ZN(n67) );
  INV_X1 U132 ( .A(n68), .ZN(n452) );
  AOI22_X1 U133 ( .A1(incPC_d[25]), .A2(n531), .B1(incPC_q[25]), .B2(n508), 
        .ZN(n68) );
  INV_X1 U134 ( .A(n69), .ZN(n451) );
  AOI22_X1 U135 ( .A1(incPC_d[24]), .A2(n531), .B1(incPC_q[24]), .B2(n508), 
        .ZN(n69) );
  INV_X1 U136 ( .A(n70), .ZN(n450) );
  AOI22_X1 U137 ( .A1(incPC_d[23]), .A2(n530), .B1(incPC_q[23]), .B2(n507), 
        .ZN(n70) );
  INV_X1 U138 ( .A(n71), .ZN(n449) );
  AOI22_X1 U139 ( .A1(incPC_d[22]), .A2(n530), .B1(incPC_q[22]), .B2(n507), 
        .ZN(n71) );
  INV_X1 U140 ( .A(n72), .ZN(n448) );
  AOI22_X1 U141 ( .A1(incPC_d[21]), .A2(n530), .B1(incPC_q[21]), .B2(n507), 
        .ZN(n72) );
  INV_X1 U142 ( .A(n73), .ZN(n447) );
  AOI22_X1 U143 ( .A1(incPC_d[20]), .A2(n530), .B1(incPC_q[20]), .B2(n507), 
        .ZN(n73) );
  INV_X1 U144 ( .A(n74), .ZN(n428) );
  AOI22_X1 U145 ( .A1(incPC_d[1]), .A2(n530), .B1(incPC_q[1]), .B2(n507), .ZN(
        n74) );
  INV_X1 U146 ( .A(n75), .ZN(n446) );
  AOI22_X1 U147 ( .A1(incPC_d[19]), .A2(n530), .B1(incPC_q[19]), .B2(n507), 
        .ZN(n75) );
  INV_X1 U148 ( .A(n76), .ZN(n445) );
  AOI22_X1 U149 ( .A1(incPC_d[18]), .A2(n530), .B1(incPC_q[18]), .B2(n507), 
        .ZN(n76) );
  INV_X1 U150 ( .A(n77), .ZN(n444) );
  AOI22_X1 U151 ( .A1(incPC_d[17]), .A2(n530), .B1(incPC_q[17]), .B2(n507), 
        .ZN(n77) );
  INV_X1 U152 ( .A(n78), .ZN(n443) );
  AOI22_X1 U153 ( .A1(incPC_d[16]), .A2(n530), .B1(incPC_q[16]), .B2(n507), 
        .ZN(n78) );
  INV_X1 U154 ( .A(n79), .ZN(n442) );
  AOI22_X1 U155 ( .A1(incPC_d[15]), .A2(n530), .B1(incPC_q[15]), .B2(n507), 
        .ZN(n79) );
  INV_X1 U156 ( .A(n80), .ZN(n441) );
  AOI22_X1 U157 ( .A1(incPC_d[14]), .A2(n530), .B1(incPC_q[14]), .B2(n507), 
        .ZN(n80) );
  INV_X1 U158 ( .A(n81), .ZN(n440) );
  AOI22_X1 U159 ( .A1(incPC_d[13]), .A2(n530), .B1(incPC_q[13]), .B2(n507), 
        .ZN(n81) );
  INV_X1 U160 ( .A(n82), .ZN(n439) );
  AOI22_X1 U161 ( .A1(incPC_d[12]), .A2(n529), .B1(incPC_q[12]), .B2(n506), 
        .ZN(n82) );
  INV_X1 U162 ( .A(n83), .ZN(n438) );
  AOI22_X1 U163 ( .A1(incPC_d[11]), .A2(n529), .B1(incPC_q[11]), .B2(n506), 
        .ZN(n83) );
  INV_X1 U164 ( .A(n84), .ZN(n437) );
  AOI22_X1 U165 ( .A1(incPC_d[10]), .A2(n529), .B1(incPC_q[10]), .B2(n506), 
        .ZN(n84) );
  INV_X1 U166 ( .A(n85), .ZN(n427) );
  AOI22_X1 U167 ( .A1(incPC_d[0]), .A2(n529), .B1(incPC_q[0]), .B2(n506), .ZN(
        n85) );
  INV_X1 U168 ( .A(n86), .ZN(n340) );
  AOI22_X1 U169 ( .A1(imm32_d[9]), .A2(n529), .B1(imm32_q[9]), .B2(n506), .ZN(
        n86) );
  INV_X1 U170 ( .A(n87), .ZN(n339) );
  AOI22_X1 U171 ( .A1(imm32_d[8]), .A2(n529), .B1(imm32_q[8]), .B2(n506), .ZN(
        n87) );
  INV_X1 U172 ( .A(n88), .ZN(n338) );
  AOI22_X1 U173 ( .A1(imm32_d[7]), .A2(n529), .B1(imm32_q[7]), .B2(n506), .ZN(
        n88) );
  INV_X1 U174 ( .A(n89), .ZN(n337) );
  AOI22_X1 U175 ( .A1(imm32_d[6]), .A2(n529), .B1(imm32_q[6]), .B2(n506), .ZN(
        n89) );
  INV_X1 U176 ( .A(n90), .ZN(n336) );
  AOI22_X1 U177 ( .A1(imm32_d[5]), .A2(n529), .B1(imm32_q[5]), .B2(n506), .ZN(
        n90) );
  INV_X1 U178 ( .A(n91), .ZN(n335) );
  AOI22_X1 U179 ( .A1(imm32_d[4]), .A2(n529), .B1(imm32_q[4]), .B2(n506), .ZN(
        n91) );
  INV_X1 U180 ( .A(n92), .ZN(n334) );
  AOI22_X1 U181 ( .A1(imm32_d[3]), .A2(n529), .B1(imm32_q[3]), .B2(n506), .ZN(
        n92) );
  INV_X1 U182 ( .A(n93), .ZN(n362) );
  AOI22_X1 U183 ( .A1(imm32_d[31]), .A2(n529), .B1(imm32_q[31]), .B2(n506), 
        .ZN(n93) );
  INV_X1 U184 ( .A(n94), .ZN(n361) );
  AOI22_X1 U185 ( .A1(imm32_d[30]), .A2(n528), .B1(imm32_q[30]), .B2(n505), 
        .ZN(n94) );
  INV_X1 U186 ( .A(n95), .ZN(n333) );
  AOI22_X1 U187 ( .A1(imm32_d[2]), .A2(n528), .B1(imm32_q[2]), .B2(n505), .ZN(
        n95) );
  INV_X1 U188 ( .A(n96), .ZN(n360) );
  AOI22_X1 U189 ( .A1(imm32_d[29]), .A2(n528), .B1(imm32_q[29]), .B2(n505), 
        .ZN(n96) );
  INV_X1 U190 ( .A(n97), .ZN(n359) );
  AOI22_X1 U191 ( .A1(imm32_d[28]), .A2(n528), .B1(imm32_q[28]), .B2(n505), 
        .ZN(n97) );
  INV_X1 U192 ( .A(n98), .ZN(n358) );
  AOI22_X1 U193 ( .A1(imm32_d[27]), .A2(n528), .B1(imm32_q[27]), .B2(n505), 
        .ZN(n98) );
  INV_X1 U194 ( .A(n99), .ZN(n357) );
  AOI22_X1 U195 ( .A1(imm32_d[26]), .A2(n528), .B1(imm32_q[26]), .B2(n505), 
        .ZN(n99) );
  INV_X1 U196 ( .A(n100), .ZN(n356) );
  AOI22_X1 U197 ( .A1(imm32_d[25]), .A2(n528), .B1(imm32_q[25]), .B2(n505), 
        .ZN(n100) );
  INV_X1 U198 ( .A(n101), .ZN(n355) );
  AOI22_X1 U199 ( .A1(imm32_d[24]), .A2(n528), .B1(imm32_q[24]), .B2(n505), 
        .ZN(n101) );
  INV_X1 U200 ( .A(n102), .ZN(n354) );
  AOI22_X1 U201 ( .A1(imm32_d[23]), .A2(n528), .B1(imm32_q[23]), .B2(n505), 
        .ZN(n102) );
  INV_X1 U202 ( .A(n103), .ZN(n353) );
  AOI22_X1 U203 ( .A1(imm32_d[22]), .A2(n528), .B1(imm32_q[22]), .B2(n505), 
        .ZN(n103) );
  INV_X1 U204 ( .A(n104), .ZN(n352) );
  AOI22_X1 U205 ( .A1(imm32_d[21]), .A2(n528), .B1(imm32_q[21]), .B2(n505), 
        .ZN(n104) );
  INV_X1 U206 ( .A(n105), .ZN(n351) );
  AOI22_X1 U207 ( .A1(imm32_d[20]), .A2(n527), .B1(imm32_q[20]), .B2(n504), 
        .ZN(n105) );
  INV_X1 U208 ( .A(n106), .ZN(n332) );
  AOI22_X1 U209 ( .A1(imm32_d[1]), .A2(n527), .B1(imm32_q[1]), .B2(n504), .ZN(
        n106) );
  INV_X1 U210 ( .A(n107), .ZN(n350) );
  AOI22_X1 U211 ( .A1(imm32_d[19]), .A2(n527), .B1(imm32_q[19]), .B2(n504), 
        .ZN(n107) );
  INV_X1 U212 ( .A(n108), .ZN(n349) );
  AOI22_X1 U213 ( .A1(imm32_d[18]), .A2(n527), .B1(imm32_q[18]), .B2(n504), 
        .ZN(n108) );
  INV_X1 U214 ( .A(n109), .ZN(n348) );
  AOI22_X1 U215 ( .A1(imm32_d[17]), .A2(n528), .B1(imm32_q[17]), .B2(n505), 
        .ZN(n109) );
  INV_X1 U216 ( .A(n110), .ZN(n347) );
  AOI22_X1 U217 ( .A1(imm32_d[16]), .A2(n527), .B1(imm32_q[16]), .B2(n504), 
        .ZN(n110) );
  INV_X1 U218 ( .A(n111), .ZN(n346) );
  AOI22_X1 U219 ( .A1(imm32_d[15]), .A2(n527), .B1(imm32_q[15]), .B2(n504), 
        .ZN(n111) );
  INV_X1 U220 ( .A(n112), .ZN(n345) );
  AOI22_X1 U221 ( .A1(imm32_d[14]), .A2(n527), .B1(imm32_q[14]), .B2(n504), 
        .ZN(n112) );
  INV_X1 U222 ( .A(n113), .ZN(n344) );
  AOI22_X1 U223 ( .A1(imm32_d[13]), .A2(n527), .B1(imm32_q[13]), .B2(n504), 
        .ZN(n113) );
  INV_X1 U224 ( .A(n114), .ZN(n343) );
  AOI22_X1 U225 ( .A1(imm32_d[12]), .A2(n527), .B1(imm32_q[12]), .B2(n504), 
        .ZN(n114) );
  INV_X1 U226 ( .A(n115), .ZN(n342) );
  AOI22_X1 U227 ( .A1(imm32_d[11]), .A2(n527), .B1(imm32_q[11]), .B2(n504), 
        .ZN(n115) );
  INV_X1 U228 ( .A(n116), .ZN(n341) );
  AOI22_X1 U229 ( .A1(imm32_d[10]), .A2(n527), .B1(imm32_q[10]), .B2(n504), 
        .ZN(n116) );
  INV_X1 U230 ( .A(n117), .ZN(n331) );
  AOI22_X1 U231 ( .A1(imm32_d[0]), .A2(n526), .B1(imm32_q[0]), .B2(n503), .ZN(
        n117) );
  INV_X1 U232 ( .A(n118), .ZN(n256) );
  AOI22_X1 U233 ( .A1(fp_d), .A2(n527), .B1(fp_q), .B2(n504), .ZN(n118) );
  INV_X1 U234 ( .A(n119), .ZN(n492) );
  AOI22_X1 U235 ( .A1(dSize_d[1]), .A2(n120), .B1(dSize_q[1]), .B2(n121), .ZN(
        n119) );
  INV_X1 U236 ( .A(n122), .ZN(n491) );
  AOI22_X1 U237 ( .A1(dSize_d[0]), .A2(n120), .B1(dSize_q[0]), .B2(n121), .ZN(
        n122) );
  INV_X1 U238 ( .A(n121), .ZN(n120) );
  NAND2_X1 U239 ( .A1(n561), .A2(n524), .ZN(n121) );
  INV_X1 U240 ( .A(n123), .ZN(n308) );
  AOI22_X1 U241 ( .A1(busFP_d[9]), .A2(n526), .B1(busFP_q[9]), .B2(n503), .ZN(
        n123) );
  INV_X1 U242 ( .A(n124), .ZN(n307) );
  AOI22_X1 U243 ( .A1(busFP_d[8]), .A2(n526), .B1(busFP_q[8]), .B2(n503), .ZN(
        n124) );
  INV_X1 U244 ( .A(n125), .ZN(n306) );
  AOI22_X1 U245 ( .A1(busFP_d[7]), .A2(n526), .B1(busFP_q[7]), .B2(n503), .ZN(
        n125) );
  INV_X1 U246 ( .A(n126), .ZN(n305) );
  AOI22_X1 U247 ( .A1(busFP_d[6]), .A2(n526), .B1(busFP_q[6]), .B2(n503), .ZN(
        n126) );
  INV_X1 U248 ( .A(n127), .ZN(n304) );
  AOI22_X1 U249 ( .A1(busFP_d[5]), .A2(n526), .B1(busFP_q[5]), .B2(n503), .ZN(
        n127) );
  INV_X1 U250 ( .A(n128), .ZN(n303) );
  AOI22_X1 U251 ( .A1(busFP_d[4]), .A2(n526), .B1(busFP_q[4]), .B2(n503), .ZN(
        n128) );
  INV_X1 U252 ( .A(n129), .ZN(n302) );
  AOI22_X1 U253 ( .A1(busFP_d[3]), .A2(n531), .B1(busFP_q[3]), .B2(n508), .ZN(
        n129) );
  INV_X1 U254 ( .A(n130), .ZN(n330) );
  AOI22_X1 U255 ( .A1(busFP_d[31]), .A2(n544), .B1(busFP_q[31]), .B2(n521), 
        .ZN(n130) );
  INV_X1 U256 ( .A(n131), .ZN(n329) );
  AOI22_X1 U257 ( .A1(busFP_d[30]), .A2(n535), .B1(busFP_q[30]), .B2(n522), 
        .ZN(n131) );
  INV_X1 U258 ( .A(n132), .ZN(n301) );
  AOI22_X1 U259 ( .A1(busFP_d[2]), .A2(n533), .B1(busFP_q[2]), .B2(n522), .ZN(
        n132) );
  INV_X1 U260 ( .A(n133), .ZN(n328) );
  AOI22_X1 U261 ( .A1(busFP_d[29]), .A2(n534), .B1(busFP_q[29]), .B2(n522), 
        .ZN(n133) );
  INV_X1 U262 ( .A(n134), .ZN(n327) );
  AOI22_X1 U263 ( .A1(busFP_d[28]), .A2(n545), .B1(busFP_q[28]), .B2(n522), 
        .ZN(n134) );
  INV_X1 U264 ( .A(n135), .ZN(n326) );
  AOI22_X1 U265 ( .A1(busFP_d[27]), .A2(n545), .B1(busFP_q[27]), .B2(n521), 
        .ZN(n135) );
  INV_X1 U266 ( .A(n136), .ZN(n325) );
  AOI22_X1 U267 ( .A1(busFP_d[26]), .A2(n545), .B1(busFP_q[26]), .B2(n521), 
        .ZN(n136) );
  INV_X1 U268 ( .A(n137), .ZN(n324) );
  AOI22_X1 U269 ( .A1(busFP_d[25]), .A2(n545), .B1(busFP_q[25]), .B2(n521), 
        .ZN(n137) );
  INV_X1 U270 ( .A(n138), .ZN(n323) );
  AOI22_X1 U271 ( .A1(busFP_d[24]), .A2(n545), .B1(busFP_q[24]), .B2(n521), 
        .ZN(n138) );
  INV_X1 U272 ( .A(n139), .ZN(n322) );
  AOI22_X1 U273 ( .A1(busFP_d[23]), .A2(n545), .B1(busFP_q[23]), .B2(n521), 
        .ZN(n139) );
  INV_X1 U274 ( .A(n140), .ZN(n321) );
  AOI22_X1 U275 ( .A1(busFP_d[22]), .A2(n545), .B1(busFP_q[22]), .B2(n521), 
        .ZN(n140) );
  INV_X1 U276 ( .A(n141), .ZN(n320) );
  AOI22_X1 U277 ( .A1(busFP_d[21]), .A2(n545), .B1(busFP_q[21]), .B2(n521), 
        .ZN(n141) );
  INV_X1 U278 ( .A(n142), .ZN(n319) );
  AOI22_X1 U279 ( .A1(busFP_d[20]), .A2(n545), .B1(busFP_q[20]), .B2(n521), 
        .ZN(n142) );
  INV_X1 U280 ( .A(n143), .ZN(n300) );
  AOI22_X1 U281 ( .A1(busFP_d[1]), .A2(n545), .B1(busFP_q[1]), .B2(n521), .ZN(
        n143) );
  INV_X1 U282 ( .A(n144), .ZN(n318) );
  AOI22_X1 U283 ( .A1(busFP_d[19]), .A2(n545), .B1(busFP_q[19]), .B2(n521), 
        .ZN(n144) );
  INV_X1 U284 ( .A(n145), .ZN(n317) );
  AOI22_X1 U285 ( .A1(busFP_d[18]), .A2(n545), .B1(busFP_q[18]), .B2(n520), 
        .ZN(n145) );
  INV_X1 U286 ( .A(n146), .ZN(n316) );
  AOI22_X1 U287 ( .A1(busFP_d[17]), .A2(n544), .B1(busFP_q[17]), .B2(n521), 
        .ZN(n146) );
  INV_X1 U288 ( .A(n147), .ZN(n315) );
  AOI22_X1 U289 ( .A1(busFP_d[16]), .A2(n544), .B1(busFP_q[16]), .B2(n520), 
        .ZN(n147) );
  INV_X1 U290 ( .A(n148), .ZN(n314) );
  AOI22_X1 U291 ( .A1(busFP_d[15]), .A2(n544), .B1(busFP_q[15]), .B2(n520), 
        .ZN(n148) );
  INV_X1 U292 ( .A(n149), .ZN(n313) );
  AOI22_X1 U293 ( .A1(busFP_d[14]), .A2(n544), .B1(busFP_q[14]), .B2(n520), 
        .ZN(n149) );
  INV_X1 U294 ( .A(n150), .ZN(n312) );
  AOI22_X1 U295 ( .A1(busFP_d[13]), .A2(n544), .B1(busFP_q[13]), .B2(n520), 
        .ZN(n150) );
  INV_X1 U296 ( .A(n151), .ZN(n311) );
  AOI22_X1 U297 ( .A1(busFP_d[12]), .A2(n544), .B1(busFP_q[12]), .B2(n520), 
        .ZN(n151) );
  INV_X1 U298 ( .A(n152), .ZN(n310) );
  AOI22_X1 U299 ( .A1(busFP_d[11]), .A2(n544), .B1(busFP_q[11]), .B2(n520), 
        .ZN(n152) );
  INV_X1 U300 ( .A(n153), .ZN(n309) );
  AOI22_X1 U301 ( .A1(busFP_d[10]), .A2(n544), .B1(busFP_q[10]), .B2(n520), 
        .ZN(n153) );
  INV_X1 U302 ( .A(n154), .ZN(n299) );
  AOI22_X1 U303 ( .A1(busFP_d[0]), .A2(n544), .B1(busFP_q[0]), .B2(n520), .ZN(
        n154) );
  INV_X1 U304 ( .A(n155), .ZN(n372) );
  AOI22_X1 U305 ( .A1(busB_d[9]), .A2(n544), .B1(busB_q[9]), .B2(n519), .ZN(
        n155) );
  INV_X1 U306 ( .A(n156), .ZN(n371) );
  AOI22_X1 U307 ( .A1(busB_d[8]), .A2(n544), .B1(busB_q[8]), .B2(n520), .ZN(
        n156) );
  INV_X1 U308 ( .A(n157), .ZN(n370) );
  AOI22_X1 U309 ( .A1(busB_d[7]), .A2(n544), .B1(busB_q[7]), .B2(n520), .ZN(
        n157) );
  INV_X1 U310 ( .A(n158), .ZN(n369) );
  AOI22_X1 U311 ( .A1(busB_d[6]), .A2(n543), .B1(busB_q[6]), .B2(n520), .ZN(
        n158) );
  INV_X1 U312 ( .A(n159), .ZN(n368) );
  AOI22_X1 U313 ( .A1(busB_d[5]), .A2(n543), .B1(busB_q[5]), .B2(n519), .ZN(
        n159) );
  INV_X1 U314 ( .A(n160), .ZN(n367) );
  AOI22_X1 U315 ( .A1(busB_d[4]), .A2(n543), .B1(busB_q[4]), .B2(n519), .ZN(
        n160) );
  INV_X1 U316 ( .A(n161), .ZN(n366) );
  AOI22_X1 U317 ( .A1(busB_d[3]), .A2(n543), .B1(busB_q[3]), .B2(n519), .ZN(
        n161) );
  INV_X1 U318 ( .A(n162), .ZN(n394) );
  AOI22_X1 U319 ( .A1(busB_d[31]), .A2(n543), .B1(busB_q[31]), .B2(n519), .ZN(
        n162) );
  INV_X1 U320 ( .A(n163), .ZN(n393) );
  AOI22_X1 U321 ( .A1(busB_d[30]), .A2(n543), .B1(busB_q[30]), .B2(n519), .ZN(
        n163) );
  INV_X1 U322 ( .A(n164), .ZN(n365) );
  AOI22_X1 U323 ( .A1(busB_d[2]), .A2(n543), .B1(busB_q[2]), .B2(n519), .ZN(
        n164) );
  INV_X1 U324 ( .A(n165), .ZN(n392) );
  AOI22_X1 U325 ( .A1(busB_d[29]), .A2(n543), .B1(busB_q[29]), .B2(n519), .ZN(
        n165) );
  INV_X1 U326 ( .A(n166), .ZN(n391) );
  AOI22_X1 U327 ( .A1(busB_d[28]), .A2(n543), .B1(busB_q[28]), .B2(n519), .ZN(
        n166) );
  INV_X1 U328 ( .A(n167), .ZN(n390) );
  AOI22_X1 U329 ( .A1(busB_d[27]), .A2(n543), .B1(busB_q[27]), .B2(n519), .ZN(
        n167) );
  INV_X1 U330 ( .A(n168), .ZN(n389) );
  AOI22_X1 U331 ( .A1(busB_d[26]), .A2(n543), .B1(busB_q[26]), .B2(n519), .ZN(
        n168) );
  INV_X1 U332 ( .A(n169), .ZN(n388) );
  AOI22_X1 U333 ( .A1(busB_d[25]), .A2(n543), .B1(busB_q[25]), .B2(n519), .ZN(
        n169) );
  INV_X1 U334 ( .A(n170), .ZN(n387) );
  AOI22_X1 U335 ( .A1(busB_d[24]), .A2(n542), .B1(busB_q[24]), .B2(n518), .ZN(
        n170) );
  INV_X1 U336 ( .A(n171), .ZN(n386) );
  AOI22_X1 U337 ( .A1(busB_d[23]), .A2(n542), .B1(busB_q[23]), .B2(n518), .ZN(
        n171) );
  INV_X1 U338 ( .A(n172), .ZN(n385) );
  AOI22_X1 U339 ( .A1(busB_d[22]), .A2(n542), .B1(busB_q[22]), .B2(n518), .ZN(
        n172) );
  INV_X1 U340 ( .A(n173), .ZN(n384) );
  AOI22_X1 U341 ( .A1(busB_d[21]), .A2(n542), .B1(busB_q[21]), .B2(n518), .ZN(
        n173) );
  INV_X1 U342 ( .A(n174), .ZN(n383) );
  AOI22_X1 U343 ( .A1(busB_d[20]), .A2(n542), .B1(busB_q[20]), .B2(n518), .ZN(
        n174) );
  INV_X1 U344 ( .A(n175), .ZN(n364) );
  AOI22_X1 U345 ( .A1(busB_d[1]), .A2(n542), .B1(busB_q[1]), .B2(n518), .ZN(
        n175) );
  INV_X1 U346 ( .A(n176), .ZN(n382) );
  AOI22_X1 U347 ( .A1(busB_d[19]), .A2(n542), .B1(busB_q[19]), .B2(n518), .ZN(
        n176) );
  INV_X1 U348 ( .A(n177), .ZN(n381) );
  AOI22_X1 U349 ( .A1(busB_d[18]), .A2(n542), .B1(busB_q[18]), .B2(n518), .ZN(
        n177) );
  INV_X1 U350 ( .A(n178), .ZN(n380) );
  AOI22_X1 U351 ( .A1(busB_d[17]), .A2(n542), .B1(busB_q[17]), .B2(n518), .ZN(
        n178) );
  INV_X1 U352 ( .A(n179), .ZN(n379) );
  AOI22_X1 U353 ( .A1(busB_d[16]), .A2(n542), .B1(busB_q[16]), .B2(n518), .ZN(
        n179) );
  INV_X1 U354 ( .A(n180), .ZN(n378) );
  AOI22_X1 U355 ( .A1(busB_d[15]), .A2(n542), .B1(busB_q[15]), .B2(n518), .ZN(
        n180) );
  INV_X1 U356 ( .A(n181), .ZN(n377) );
  AOI22_X1 U357 ( .A1(busB_d[14]), .A2(n542), .B1(busB_q[14]), .B2(n518), .ZN(
        n181) );
  INV_X1 U358 ( .A(n182), .ZN(n376) );
  AOI22_X1 U359 ( .A1(busB_d[13]), .A2(n541), .B1(busB_q[13]), .B2(n517), .ZN(
        n182) );
  INV_X1 U360 ( .A(n183), .ZN(n375) );
  AOI22_X1 U361 ( .A1(busB_d[12]), .A2(n541), .B1(busB_q[12]), .B2(n517), .ZN(
        n183) );
  INV_X1 U362 ( .A(n184), .ZN(n374) );
  AOI22_X1 U363 ( .A1(busB_d[11]), .A2(n541), .B1(busB_q[11]), .B2(n517), .ZN(
        n184) );
  INV_X1 U364 ( .A(n185), .ZN(n373) );
  AOI22_X1 U365 ( .A1(busB_d[10]), .A2(n541), .B1(busB_q[10]), .B2(n517), .ZN(
        n185) );
  INV_X1 U366 ( .A(n186), .ZN(n363) );
  AOI22_X1 U367 ( .A1(busB_d[0]), .A2(n541), .B1(busB_q[0]), .B2(n517), .ZN(
        n186) );
  INV_X1 U368 ( .A(n187), .ZN(n404) );
  AOI22_X1 U369 ( .A1(busA_d[9]), .A2(n541), .B1(busA_q[9]), .B2(n517), .ZN(
        n187) );
  INV_X1 U370 ( .A(n188), .ZN(n403) );
  AOI22_X1 U371 ( .A1(busA_d[8]), .A2(n541), .B1(busA_q[8]), .B2(n517), .ZN(
        n188) );
  INV_X1 U372 ( .A(n189), .ZN(n402) );
  AOI22_X1 U373 ( .A1(busA_d[7]), .A2(n541), .B1(busA_q[7]), .B2(n517), .ZN(
        n189) );
  INV_X1 U374 ( .A(n190), .ZN(n401) );
  AOI22_X1 U375 ( .A1(busA_d[6]), .A2(n541), .B1(busA_q[6]), .B2(n517), .ZN(
        n190) );
  INV_X1 U376 ( .A(n191), .ZN(n400) );
  AOI22_X1 U377 ( .A1(busA_d[5]), .A2(n541), .B1(busA_q[5]), .B2(n517), .ZN(
        n191) );
  INV_X1 U378 ( .A(n192), .ZN(n399) );
  AOI22_X1 U379 ( .A1(busA_d[4]), .A2(n541), .B1(busA_q[4]), .B2(n517), .ZN(
        n192) );
  INV_X1 U380 ( .A(n193), .ZN(n398) );
  AOI22_X1 U381 ( .A1(busA_d[3]), .A2(n540), .B1(busA_q[3]), .B2(n516), .ZN(
        n193) );
  INV_X1 U382 ( .A(n194), .ZN(n426) );
  AOI22_X1 U383 ( .A1(busA_d[31]), .A2(n540), .B1(busA_q[31]), .B2(n516), .ZN(
        n194) );
  INV_X1 U384 ( .A(n195), .ZN(n425) );
  AOI22_X1 U385 ( .A1(busA_d[30]), .A2(n540), .B1(busA_q[30]), .B2(n516), .ZN(
        n195) );
  INV_X1 U386 ( .A(n196), .ZN(n397) );
  AOI22_X1 U387 ( .A1(busA_d[2]), .A2(n540), .B1(busA_q[2]), .B2(n516), .ZN(
        n196) );
  INV_X1 U388 ( .A(n197), .ZN(n424) );
  AOI22_X1 U389 ( .A1(busA_d[29]), .A2(n540), .B1(busA_q[29]), .B2(n516), .ZN(
        n197) );
  INV_X1 U390 ( .A(n198), .ZN(n423) );
  AOI22_X1 U391 ( .A1(busA_d[28]), .A2(n540), .B1(busA_q[28]), .B2(n516), .ZN(
        n198) );
  INV_X1 U392 ( .A(n199), .ZN(n422) );
  AOI22_X1 U393 ( .A1(busA_d[27]), .A2(n540), .B1(busA_q[27]), .B2(n516), .ZN(
        n199) );
  INV_X1 U394 ( .A(n200), .ZN(n421) );
  AOI22_X1 U395 ( .A1(busA_d[26]), .A2(n540), .B1(busA_q[26]), .B2(n516), .ZN(
        n200) );
  INV_X1 U396 ( .A(n201), .ZN(n420) );
  AOI22_X1 U397 ( .A1(busA_d[25]), .A2(n540), .B1(busA_q[25]), .B2(n516), .ZN(
        n201) );
  INV_X1 U398 ( .A(n202), .ZN(n419) );
  AOI22_X1 U399 ( .A1(busA_d[24]), .A2(n540), .B1(busA_q[24]), .B2(n516), .ZN(
        n202) );
  INV_X1 U400 ( .A(n203), .ZN(n418) );
  AOI22_X1 U401 ( .A1(busA_d[23]), .A2(n540), .B1(busA_q[23]), .B2(n516), .ZN(
        n203) );
  INV_X1 U402 ( .A(n204), .ZN(n417) );
  AOI22_X1 U403 ( .A1(busA_d[22]), .A2(n540), .B1(busA_q[22]), .B2(n516), .ZN(
        n204) );
  INV_X1 U404 ( .A(n205), .ZN(n416) );
  AOI22_X1 U405 ( .A1(busA_d[21]), .A2(n539), .B1(busA_q[21]), .B2(n515), .ZN(
        n205) );
  INV_X1 U406 ( .A(n206), .ZN(n415) );
  AOI22_X1 U407 ( .A1(busA_d[20]), .A2(n539), .B1(busA_q[20]), .B2(n515), .ZN(
        n206) );
  INV_X1 U408 ( .A(n207), .ZN(n396) );
  AOI22_X1 U409 ( .A1(busA_d[1]), .A2(n539), .B1(busA_q[1]), .B2(n515), .ZN(
        n207) );
  INV_X1 U410 ( .A(n208), .ZN(n414) );
  AOI22_X1 U411 ( .A1(busA_d[19]), .A2(n539), .B1(busA_q[19]), .B2(n515), .ZN(
        n208) );
  INV_X1 U412 ( .A(n209), .ZN(n413) );
  AOI22_X1 U413 ( .A1(busA_d[18]), .A2(n539), .B1(busA_q[18]), .B2(n515), .ZN(
        n209) );
  INV_X1 U414 ( .A(n210), .ZN(n412) );
  AOI22_X1 U415 ( .A1(busA_d[17]), .A2(n539), .B1(busA_q[17]), .B2(n515), .ZN(
        n210) );
  INV_X1 U416 ( .A(n211), .ZN(n411) );
  AOI22_X1 U417 ( .A1(busA_d[16]), .A2(n539), .B1(busA_q[16]), .B2(n515), .ZN(
        n211) );
  INV_X1 U418 ( .A(n212), .ZN(n410) );
  AOI22_X1 U419 ( .A1(busA_d[15]), .A2(n539), .B1(busA_q[15]), .B2(n515), .ZN(
        n212) );
  INV_X1 U420 ( .A(n213), .ZN(n409) );
  AOI22_X1 U421 ( .A1(busA_d[14]), .A2(n539), .B1(busA_q[14]), .B2(n515), .ZN(
        n213) );
  INV_X1 U422 ( .A(n214), .ZN(n408) );
  AOI22_X1 U423 ( .A1(busA_d[13]), .A2(n539), .B1(busA_q[13]), .B2(n515), .ZN(
        n214) );
  INV_X1 U424 ( .A(n215), .ZN(n407) );
  AOI22_X1 U425 ( .A1(busA_d[12]), .A2(n539), .B1(busA_q[12]), .B2(n515), .ZN(
        n215) );
  INV_X1 U426 ( .A(n216), .ZN(n406) );
  AOI22_X1 U427 ( .A1(busA_d[11]), .A2(n539), .B1(busA_q[11]), .B2(n515), .ZN(
        n216) );
  INV_X1 U428 ( .A(n217), .ZN(n405) );
  AOI22_X1 U429 ( .A1(busA_d[10]), .A2(n538), .B1(busA_q[10]), .B2(n514), .ZN(
        n217) );
  INV_X1 U430 ( .A(n218), .ZN(n395) );
  AOI22_X1 U431 ( .A1(busA_d[0]), .A2(n538), .B1(busA_q[0]), .B2(n514), .ZN(
        n218) );
  INV_X1 U432 ( .A(n219), .ZN(n260) );
  AOI22_X1 U433 ( .A1(branch_d), .A2(n538), .B1(branch_q), .B2(n514), .ZN(n219) );
  INV_X1 U434 ( .A(n220), .ZN(n276) );
  AOI22_X1 U435 ( .A1(aluRes_d[9]), .A2(n538), .B1(aluRes_q[9]), .B2(n514), 
        .ZN(n220) );
  INV_X1 U436 ( .A(n221), .ZN(n275) );
  AOI22_X1 U437 ( .A1(aluRes_d[8]), .A2(n538), .B1(aluRes_q[8]), .B2(n514), 
        .ZN(n221) );
  INV_X1 U438 ( .A(n222), .ZN(n274) );
  AOI22_X1 U439 ( .A1(aluRes_d[7]), .A2(n538), .B1(aluRes_q[7]), .B2(n514), 
        .ZN(n222) );
  INV_X1 U440 ( .A(n223), .ZN(n273) );
  AOI22_X1 U441 ( .A1(aluRes_d[6]), .A2(n538), .B1(aluRes_q[6]), .B2(n514), 
        .ZN(n223) );
  INV_X1 U442 ( .A(n224), .ZN(n272) );
  AOI22_X1 U443 ( .A1(aluRes_d[5]), .A2(n538), .B1(aluRes_q[5]), .B2(n514), 
        .ZN(n224) );
  INV_X1 U444 ( .A(n225), .ZN(n271) );
  AOI22_X1 U445 ( .A1(aluRes_d[4]), .A2(n538), .B1(aluRes_q[4]), .B2(n514), 
        .ZN(n225) );
  INV_X1 U446 ( .A(n226), .ZN(n270) );
  AOI22_X1 U447 ( .A1(aluRes_d[3]), .A2(n538), .B1(aluRes_q[3]), .B2(n514), 
        .ZN(n226) );
  INV_X1 U448 ( .A(n227), .ZN(n298) );
  AOI22_X1 U449 ( .A1(aluRes_d[31]), .A2(n538), .B1(aluRes_q[31]), .B2(n514), 
        .ZN(n227) );
  INV_X1 U450 ( .A(n228), .ZN(n297) );
  AOI22_X1 U451 ( .A1(aluRes_d[30]), .A2(n538), .B1(aluRes_q[30]), .B2(n514), 
        .ZN(n228) );
  INV_X1 U452 ( .A(n229), .ZN(n269) );
  AOI22_X1 U453 ( .A1(aluRes_d[2]), .A2(n537), .B1(aluRes_q[2]), .B2(n513), 
        .ZN(n229) );
  INV_X1 U454 ( .A(n230), .ZN(n296) );
  AOI22_X1 U455 ( .A1(aluRes_d[29]), .A2(n537), .B1(aluRes_q[29]), .B2(n513), 
        .ZN(n230) );
  INV_X1 U456 ( .A(n231), .ZN(n295) );
  AOI22_X1 U457 ( .A1(aluRes_d[28]), .A2(n537), .B1(aluRes_q[28]), .B2(n513), 
        .ZN(n231) );
  INV_X1 U458 ( .A(n232), .ZN(n294) );
  AOI22_X1 U459 ( .A1(aluRes_d[27]), .A2(n537), .B1(aluRes_q[27]), .B2(n513), 
        .ZN(n232) );
  INV_X1 U460 ( .A(n233), .ZN(n293) );
  AOI22_X1 U461 ( .A1(aluRes_d[26]), .A2(n537), .B1(aluRes_q[26]), .B2(n513), 
        .ZN(n233) );
  INV_X1 U462 ( .A(n234), .ZN(n292) );
  AOI22_X1 U463 ( .A1(aluRes_d[25]), .A2(n537), .B1(aluRes_q[25]), .B2(n513), 
        .ZN(n234) );
  INV_X1 U464 ( .A(n235), .ZN(n291) );
  AOI22_X1 U465 ( .A1(aluRes_d[24]), .A2(n537), .B1(aluRes_q[24]), .B2(n513), 
        .ZN(n235) );
  INV_X1 U466 ( .A(n236), .ZN(n290) );
  AOI22_X1 U467 ( .A1(aluRes_d[23]), .A2(n537), .B1(aluRes_q[23]), .B2(n513), 
        .ZN(n236) );
  INV_X1 U468 ( .A(n237), .ZN(n289) );
  AOI22_X1 U469 ( .A1(aluRes_d[22]), .A2(n537), .B1(aluRes_q[22]), .B2(n513), 
        .ZN(n237) );
  INV_X1 U470 ( .A(n238), .ZN(n288) );
  AOI22_X1 U471 ( .A1(aluRes_d[21]), .A2(n537), .B1(aluRes_q[21]), .B2(n513), 
        .ZN(n238) );
  INV_X1 U472 ( .A(n239), .ZN(n287) );
  AOI22_X1 U473 ( .A1(aluRes_d[20]), .A2(n537), .B1(aluRes_q[20]), .B2(n513), 
        .ZN(n239) );
  INV_X1 U474 ( .A(n240), .ZN(n268) );
  AOI22_X1 U475 ( .A1(aluRes_d[1]), .A2(n537), .B1(aluRes_q[1]), .B2(n513), 
        .ZN(n240) );
  INV_X1 U476 ( .A(n241), .ZN(n286) );
  AOI22_X1 U477 ( .A1(aluRes_d[19]), .A2(n536), .B1(aluRes_q[19]), .B2(n512), 
        .ZN(n241) );
  INV_X1 U478 ( .A(n242), .ZN(n285) );
  AOI22_X1 U479 ( .A1(aluRes_d[18]), .A2(n536), .B1(aluRes_q[18]), .B2(n512), 
        .ZN(n242) );
  INV_X1 U480 ( .A(n243), .ZN(n284) );
  AOI22_X1 U481 ( .A1(aluRes_d[17]), .A2(n536), .B1(aluRes_q[17]), .B2(n512), 
        .ZN(n243) );
  INV_X1 U482 ( .A(n244), .ZN(n283) );
  AOI22_X1 U483 ( .A1(aluRes_d[16]), .A2(n536), .B1(aluRes_q[16]), .B2(n512), 
        .ZN(n244) );
  INV_X1 U484 ( .A(n245), .ZN(n282) );
  AOI22_X1 U485 ( .A1(aluRes_d[15]), .A2(n536), .B1(aluRes_q[15]), .B2(n512), 
        .ZN(n245) );
  INV_X1 U486 ( .A(n246), .ZN(n281) );
  AOI22_X1 U487 ( .A1(aluRes_d[14]), .A2(n536), .B1(aluRes_q[14]), .B2(n512), 
        .ZN(n246) );
  INV_X1 U488 ( .A(n247), .ZN(n280) );
  AOI22_X1 U489 ( .A1(aluRes_d[13]), .A2(n536), .B1(aluRes_q[13]), .B2(n512), 
        .ZN(n247) );
  INV_X1 U490 ( .A(n248), .ZN(n279) );
  AOI22_X1 U491 ( .A1(aluRes_d[12]), .A2(n536), .B1(aluRes_q[12]), .B2(n512), 
        .ZN(n248) );
  INV_X1 U492 ( .A(n249), .ZN(n278) );
  AOI22_X1 U493 ( .A1(aluRes_d[11]), .A2(n536), .B1(aluRes_q[11]), .B2(n512), 
        .ZN(n249) );
  INV_X1 U494 ( .A(n250), .ZN(n277) );
  AOI22_X1 U495 ( .A1(aluRes_d[10]), .A2(n541), .B1(aluRes_q[10]), .B2(n517), 
        .ZN(n250) );
  INV_X1 U496 ( .A(n251), .ZN(n267) );
  AOI22_X1 U497 ( .A1(aluRes_d[0]), .A2(n526), .B1(aluRes_q[0]), .B2(n503), 
        .ZN(n251) );
  INV_X1 U498 ( .A(n252), .ZN(n3) );
  OAI21_X1 U499 ( .B1(ctrl[1]), .B2(ctrl[0]), .A(n253), .ZN(n252) );
  INV_X1 U500 ( .A(n253), .ZN(n2) );
  NAND2_X1 U501 ( .A1(ctrl[1]), .A2(ctrl[0]), .ZN(n253) );
  BUF_X4 U502 ( .A(n502), .Z(n513) );
  BUF_X4 U503 ( .A(n525), .Z(n537) );
  BUF_X4 U504 ( .A(n525), .Z(n545) );
  BUF_X4 U505 ( .A(n500), .Z(n522) );
  BUF_X4 U506 ( .A(n501), .Z(n521) );
  BUF_X4 U507 ( .A(n502), .Z(n504) );
  BUF_X4 U508 ( .A(n525), .Z(n527) );
  BUF_X4 U509 ( .A(n501), .Z(n505) );
  BUF_X4 U510 ( .A(n524), .Z(n528) );
  BUF_X4 U511 ( .A(n502), .Z(n520) );
  BUF_X4 U512 ( .A(n502), .Z(n518) );
  BUF_X4 U513 ( .A(n525), .Z(n542) );
  BUF_X4 U514 ( .A(n502), .Z(n519) );
  BUF_X4 U515 ( .A(n525), .Z(n543) );
  BUF_X4 U516 ( .A(n502), .Z(n517) );
  BUF_X4 U517 ( .A(n525), .Z(n541) );
  BUF_X4 U518 ( .A(n501), .Z(n514) );
  BUF_X4 U519 ( .A(n524), .Z(n538) );
  BUF_X4 U520 ( .A(n501), .Z(n515) );
  BUF_X4 U521 ( .A(n524), .Z(n539) );
  BUF_X4 U522 ( .A(n501), .Z(n516) );
  BUF_X4 U523 ( .A(n524), .Z(n540) );
  BUF_X4 U524 ( .A(n501), .Z(n506) );
  BUF_X4 U525 ( .A(n524), .Z(n529) );
  BUF_X4 U526 ( .A(n502), .Z(n507) );
  BUF_X4 U527 ( .A(n525), .Z(n530) );
  BUF_X4 U528 ( .A(n501), .Z(n508) );
  BUF_X4 U529 ( .A(n524), .Z(n531) );
  BUF_X4 U530 ( .A(n523), .Z(n532) );
  BUF_X4 U531 ( .A(n523), .Z(n533) );
  BUF_X4 U532 ( .A(n523), .Z(n534) );
  BUF_X4 U533 ( .A(n500), .Z(n503) );
  BUF_X4 U534 ( .A(n523), .Z(n526) );
  BUF_X4 U535 ( .A(n501), .Z(n512) );
  BUF_X4 U536 ( .A(n524), .Z(n536) );
  BUF_X4 U537 ( .A(rst), .Z(n546) );
  BUF_X4 U538 ( .A(rst), .Z(n547) );
  BUF_X4 U539 ( .A(rst), .Z(n548) );
  BUF_X4 U540 ( .A(rst), .Z(n549) );
  BUF_X4 U541 ( .A(rst), .Z(n550) );
  BUF_X4 U542 ( .A(rst), .Z(n551) );
  BUF_X4 U543 ( .A(rst), .Z(n552) );
  BUF_X4 U544 ( .A(rst), .Z(n556) );
  BUF_X4 U545 ( .A(rst), .Z(n553) );
  BUF_X4 U546 ( .A(rst), .Z(n561) );
  BUF_X4 U547 ( .A(n500), .Z(n511) );
  BUF_X4 U548 ( .A(n500), .Z(n510) );
  BUF_X4 U549 ( .A(n500), .Z(n509) );
  BUF_X4 U550 ( .A(n523), .Z(n544) );
  BUF_X4 U551 ( .A(n523), .Z(n535) );
  BUF_X4 U552 ( .A(rst), .Z(n555) );
  BUF_X4 U553 ( .A(rst), .Z(n554) );
  BUF_X4 U554 ( .A(n3), .Z(n502) );
  BUF_X4 U555 ( .A(n3), .Z(n501) );
  BUF_X4 U556 ( .A(n3), .Z(n500) );
  BUF_X4 U557 ( .A(n2), .Z(n525) );
  BUF_X4 U558 ( .A(n2), .Z(n524) );
  BUF_X4 U559 ( .A(n2), .Z(n523) );
  BUF_X4 U560 ( .A(rst), .Z(n560) );
  BUF_X4 U561 ( .A(rst), .Z(n559) );
  BUF_X4 U562 ( .A(rst), .Z(n558) );
  BUF_X4 U563 ( .A(rst), .Z(n557) );
endmodule

