`ifndef _constants_vh_
`define _constants_vh_

// Register 0 index
`define R0      5'b0

// Pipeline register controls
`define SQUASH  2'b00
`define GO      2'b11
`define STALL   2'b01

// Instructions
`define NOP     32'h15

`endif //_constants_vh_