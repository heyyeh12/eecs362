module if_id(clk, rst, incPC_d, instr_d, incPC_q, instr_q);

input clk, rst;
input [31:0] incPC_d, instr_d;
output [31:0] incPC_q, instr_q;


endmodule