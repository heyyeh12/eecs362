
module multiplier ( a, b, control, product_in, product_out );
  input [31:0] a;
  input [31:0] b;
  input [1:0] control;
  input [31:0] product_in;
  output [31:0] product_out;
  wire   net253043, net253044, net253049, net253050, net253056, net253057,
         net253059, net253064, net253067, net253103, net253109, net253111,
         net253156, net253163, net253173, net253176, net253177, net253179,
         net253182, net253183, net253185, net253187, net253188, net253191,
         net253192, net253193, net253194, net253198, net253204, net253205,
         net253208, net253209, net253220, net253231, net253237, net253246,
         net253270, net253271, net253272, net253273, net253274, net253278,
         net253279, net253280, net253286, net253287, net253289, net253294,
         net253295, net253296, net253301, net253304, net253308, net253322,
         net253323, net253327, net253380, net253385, net253386, net253388,
         net253390, net253391, net253392, net253393, net253396, net253398,
         net253401, net253402, net253406, net253407, net253411, net253415,
         net253419, net253421, net253425, net253431, net253442, net253443,
         net253444, net253445, net253446, net253447, net253448, net253449,
         net253450, net253451, net253452, net253453, net253457, net253458,
         net253460, net253462, net253463, net253519, net253522, net253525,
         net253533, net253535, net253547, net253553, net253557, net253564,
         net253569, net253570, net253571, net253572, net253579, net253584,
         net253586, net253588, net253591, net253592, net253643, net253646,
         net253647, net253656, net253657, net253659, net253660, net253693,
         net253694, net253697, net253701, net253762, net253763, net253764,
         net253765, net253770, net253772, net253776, net253780, net253797,
         net253808, net253810, net253815, net253816, net253819, net253820,
         net253823, net253824, net253913, net253936, net253986, net253987,
         net254001, net254004, net254051, net254052, net254054, net254057,
         net254058, net254059, net254082, net254083, net254084, net254085,
         net254086, net254094, net254179, net254184, net254188, net254189,
         net254191, net254192, net254234, net254235, net254242, net254255,
         net254283, net254285, net254290, net254291, net254293, net254296,
         net254298, net254302, net254306, net254363, net254364, net254366,
         net254390, net254411, net254414, net254415, net254459, net254464,
         net254465, net254467, net254468, net254470, net254562, net254566,
         net254567, net254575, net254576, net254577, net254628, net254631,
         net254633, net254634, net254635, net254656, net254666, net254669,
         net254670, net254671, net254675, net254681, net254682, net254683,
         net254684, net254687, net254688, net254689, net254693, net254696,
         net254756, net254760, net254761, net254766, net254767, net254770,
         net254807, net254856, net254857, net254858, net254861, net254862,
         net254864, net254869, net254871, net254872, net254873, net254932,
         net254939, net254940, net254948, net254949, net254952, net254992,
         net255040, net255044, net255045, net255046, net255047, net255089,
         net255090, net255091, net255092, net255096, net255097, net255098,
         net255101, net255102, net255104, net255105, net255106, net255164,
         net255165, net255166, net255167, net255179, net255217, net255218,
         net255223, net255225, net255226, net255229, net255231, net255232,
         net255244, net255247, net255284, net255318, net255319, net255322,
         net255324, net255328, net255341, net255374, net255375, net255376,
         net255378, net255379, net255380, net255383, net255409, net255413,
         net255425, net255426, net255428, net255429, net255430, net255433,
         net255434, net255437, net255438, net255445, net255453, net255454,
         net255456, net255457, net255458, net255459, net255484, net255489,
         net255490, net255498, net255504, net255505, net255506, net255507,
         net255533, net255537, net255538, net255540, net255542, net255543,
         net255581, net255582, net255587, net255591, net255593, net255594,
         net255605, net255606, net255611, net255616, net255624, net255626,
         net255627, net255629, net255699, net255702, net255703, net255705,
         net255708, net255714, net255718, net255720, net255721, net255724,
         net255725, net255726, net255727, net255770, net255773, net255775,
         net255776, net255777, net255779, net255785, net255790, net255855,
         net255856, net255872, net255874, net255878, net255910, net255915,
         net255916, net255929, net255936, net256018, net256032, net256033,
         net256050, net256077, net256089, net256087, net256099, net256097,
         net256095, net256111, net256105, net256119, net256117, net256127,
         net256125, net256139, net256137, net256135, net256145, net256143,
         net256141, net256153, net256151, net256147, net256159, net256157,
         net256167, net256165, net256175, net256173, net256184, net256183,
         net256290, net256303, net256306, net256305, net256334, net256362,
         net256371, net256375, net256376, net256388, net256402, net256420,
         net256527, net256541, net256556, net256555, net256583, net256582,
         net256742, net256741, net256796, net256795, net256823, net256839,
         net256843, net256860, net256874, net256907, net256909, net256927,
         net256966, net256982, net257023, net257044, net257052, net257069,
         net257068, net257109, net257127, net257159, net257171, net257211,
         net257239, net257240, net257266, net257283, net257296, net257295,
         net257343, net257401, net257407, net257456, net257481, net257485,
         net257484, net257560, net257565, net257564, net257586, net257590,
         net257589, net257630, net257650, net257661, net257672, net257678,
         net257702, net257721, net257720, net257752, net257779, net257778,
         net257828, net257838, net257864, net257880, net257953, net257979,
         net258044, net258069, net256296, net255436, net255435, net256115,
         net254140, net254050, net257522, net255583, net255443, net255442,
         net255441, net255221, net255220, net255219, net256958, net253394,
         net253320, net258007, net257031, net253689, net257435, net256800,
         net253429, net253427, net253424, net253414, net253405, net253315,
         net253206, net257772, net255875, net255870, net255617, net254711,
         net254709, net254695, net256680, net256678, net254461, net254673,
         net254570, net254463, net254462, net253804, net257392, net256627,
         net256584, net254947, net256879, net254708, net254367, net255706,
         net255427, net256060, net256059, net256058, net256054, net256748,
         net256747, net256746, net255592, net255590, net255589, net255588,
         net255585, net255584, net255548, net255547, net255546, net255440,
         net255439, net257153, net253395, net253324, net253316, net253306,
         net253305, net253169, net253775, net253653, net255100, net255099,
         net254942, net254868, net253291, net253180, net253178, net253164,
         net257363, net256990, net255320, net257693, net255619, net255618,
         net255431, net257796, net257442, net253651, net253641, net253640,
         net253583, net253582, net253580, net253441, net253423, net253422,
         net257439, net253988, net253985, net253984, net253983, net253802,
         net253801, net253806, net253805, net253800, net253761, net253758,
         net253756, net253688, net253652, net253650, net257677, net257469,
         net256045, net256044, net256042, net256041, net256040, net256039,
         net255868, net257918, net254941, net254935, net254934, net254933,
         net254867, net254755, net254238, net254233, net256421, net256069,
         net256055, net255964, net255877, net257981, net257980, net253691,
         net253690, net253687, net253685, net253662, net253433, net257254,
         net256947, net254361, net254297, net254289, net254284, net254239,
         net254237, net254232, net254231, net254147, net254145, net254143,
         net254142, net253190, net253189, net253162, net253161, net253160,
         net253058, net253039, net253038, net255329, net255327, net255325,
         net255107, net257782, net256062, net256061, net256870, net255545,
         net255503, net255502, net255501, net255500, net255499, net255335,
         net255333, net255332, net255331, net255967, net255966, net255914,
         net256103, net256101, net253302, net253166, net253165, net253053,
         net257585, net257482, net256401, net255871, net255867, net255854,
         net255853, net255852, net255796, net255795, net255622, net255613,
         net255488, net255407, net256063, net257064, net256953, net254870,
         net254865, net254863, net254753, net254752, net254751, net254690,
         net254680, net254574, net254573, net254572, net256179, net254183,
         net254182, net254181, net254180, net254150, net254149, net257703,
         net256974, net256700, net254748, net254747, net254746, net254744,
         net254743, net254571, net254460, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115;

  NAND2_X1 U1133 ( .A1(n3789), .A2(net257211), .ZN(n3769) );
  NOR2_X1 U1134 ( .A1(net257672), .A2(n3770), .ZN(n3771) );
  INV_X4 U1135 ( .A(net253445), .ZN(net257828) );
  AOI21_X4 U1136 ( .B1(net254054), .B2(n3413), .A(n3630), .ZN(n3466) );
  INV_X4 U1137 ( .A(net254180), .ZN(n1104) );
  INV_X4 U1138 ( .A(net254180), .ZN(net254150) );
  NOR2_X1 U1139 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  INV_X4 U1140 ( .A(n2833), .ZN(n2760) );
  NAND2_X4 U1141 ( .A1(n1393), .A2(n1394), .ZN(n1396) );
  INV_X2 U1142 ( .A(n1860), .ZN(n1861) );
  INV_X2 U1143 ( .A(n3690), .ZN(n1334) );
  INV_X2 U1144 ( .A(n1667), .ZN(n1105) );
  INV_X4 U1146 ( .A(n1106), .ZN(n1107) );
  NAND2_X1 U1147 ( .A1(net254462), .A2(net254463), .ZN(n1259) );
  CLKBUF_X1 U1148 ( .A(net254464), .Z(n1374) );
  OAI221_X1 U1149 ( .B1(net253308), .B2(n3918), .C1(n3917), .C2(net256184), 
        .A(n3916), .ZN(net253304) );
  NOR2_X1 U1150 ( .A1(n1723), .A2(net253304), .ZN(net253306) );
  INV_X1 U1151 ( .A(n2180), .ZN(n2181) );
  INV_X2 U1152 ( .A(net254182), .ZN(n1254) );
  NAND2_X4 U1153 ( .A1(net253763), .A2(net253762), .ZN(n1108) );
  NAND2_X2 U1154 ( .A1(net253763), .A2(net253762), .ZN(net253447) );
  NAND2_X4 U1155 ( .A1(n3161), .A2(n1776), .ZN(n3079) );
  NAND2_X2 U1156 ( .A1(n1580), .A2(n3265), .ZN(n1582) );
  INV_X8 U1157 ( .A(net257980), .ZN(net257981) );
  INV_X8 U1158 ( .A(net254001), .ZN(net254289) );
  OAI21_X2 U1159 ( .B1(net254293), .B2(n3248), .A(n3324), .ZN(n1109) );
  NAND2_X2 U1160 ( .A1(net254239), .A2(n1488), .ZN(n1632) );
  INV_X4 U1162 ( .A(n1386), .ZN(n1110) );
  INV_X8 U1163 ( .A(net255375), .ZN(n1386) );
  NAND2_X2 U1164 ( .A1(net255229), .A2(net255331), .ZN(net255375) );
  NAND2_X1 U1166 ( .A1(n3337), .A2(n1933), .ZN(n2003) );
  NAND2_X2 U1167 ( .A1(n1582), .A2(n1581), .ZN(n1956) );
  NAND2_X4 U1168 ( .A1(n2785), .A2(n2784), .ZN(n1111) );
  BUF_X16 U1169 ( .A(n4004), .Z(n1112) );
  INV_X4 U1170 ( .A(net253458), .ZN(net253453) );
  OAI211_X2 U1171 ( .C1(n3531), .C2(n1892), .A(n1436), .B(n3529), .ZN(n1113)
         );
  NAND2_X2 U1173 ( .A1(n3604), .A2(n3550), .ZN(n3383) );
  INV_X1 U1174 ( .A(n3938), .ZN(n1114) );
  INV_X2 U1175 ( .A(n1114), .ZN(n1115) );
  OAI21_X4 U1176 ( .B1(n3288), .B2(n1910), .A(n1777), .ZN(n1931) );
  NAND2_X2 U1177 ( .A1(n3942), .A2(n3897), .ZN(n3846) );
  INV_X4 U1178 ( .A(net254237), .ZN(n1488) );
  INV_X4 U1179 ( .A(net255091), .ZN(net255319) );
  XNOR2_X1 U1181 ( .A(n3970), .B(n4010), .ZN(n1116) );
  NOR2_X2 U1182 ( .A1(net257980), .A2(net253662), .ZN(net253691) );
  XNOR2_X2 U1183 ( .A(n2526), .B(n2683), .ZN(n1117) );
  NAND2_X2 U1184 ( .A1(n1486), .A2(n1487), .ZN(net256796) );
  NAND2_X2 U1185 ( .A1(n1484), .A2(n1485), .ZN(n1487) );
  NAND2_X4 U1186 ( .A1(net255100), .A2(net255099), .ZN(n1118) );
  NAND2_X4 U1187 ( .A1(net255100), .A2(net255099), .ZN(n1119) );
  INV_X2 U1188 ( .A(n1697), .ZN(n1248) );
  INV_X4 U1190 ( .A(n1558), .ZN(n1559) );
  NAND3_X2 U1191 ( .A1(n3390), .A2(n3389), .A3(net257407), .ZN(n1120) );
  INV_X4 U1192 ( .A(n3034), .ZN(n2960) );
  INV_X4 U1193 ( .A(net254680), .ZN(net254870) );
  INV_X4 U1194 ( .A(n2760), .ZN(n1121) );
  INV_X2 U1195 ( .A(n2568), .ZN(n1813) );
  NAND2_X2 U1196 ( .A1(n1931), .A2(n3412), .ZN(n1122) );
  NOR2_X4 U1197 ( .A1(n3522), .A2(n3521), .ZN(n3526) );
  INV_X4 U1198 ( .A(n1947), .ZN(n1948) );
  INV_X2 U1199 ( .A(n3500), .ZN(n3102) );
  NAND2_X4 U1200 ( .A1(net253156), .A2(n3993), .ZN(n3851) );
  INV_X2 U1202 ( .A(n3475), .ZN(n1190) );
  NAND2_X4 U1203 ( .A1(net253640), .A2(net253641), .ZN(net257442) );
  NAND2_X1 U1204 ( .A1(net253640), .A2(net253641), .ZN(net257153) );
  OAI21_X4 U1205 ( .B1(net254575), .B2(net254576), .A(net257864), .ZN(n1123)
         );
  NOR3_X2 U1207 ( .A1(net253057), .A2(n1993), .A3(n3988), .ZN(n3989) );
  INV_X4 U1208 ( .A(n1881), .ZN(n1400) );
  NAND2_X2 U1209 ( .A1(net253431), .A2(n1290), .ZN(n1558) );
  NAND2_X4 U1210 ( .A1(n3624), .A2(n3623), .ZN(n1125) );
  NAND2_X2 U1211 ( .A1(n3594), .A2(n3597), .ZN(n1338) );
  BUF_X32 U1212 ( .A(net253564), .Z(net256966) );
  INV_X4 U1213 ( .A(net254284), .ZN(n1286) );
  NAND2_X2 U1215 ( .A1(n2215), .A2(n2278), .ZN(n1520) );
  OAI21_X4 U1216 ( .B1(n2947), .B2(n2946), .A(n1261), .ZN(n2747) );
  AOI21_X2 U1217 ( .B1(n2661), .B2(n1273), .A(n2660), .ZN(n2666) );
  INV_X4 U1218 ( .A(n2485), .ZN(n1126) );
  XNOR2_X2 U1219 ( .A(n1906), .B(n2858), .ZN(product_out[16]) );
  INV_X16 U1220 ( .A(n1268), .ZN(n1906) );
  INV_X4 U1221 ( .A(n2933), .ZN(n2934) );
  NAND2_X4 U1222 ( .A1(n1816), .A2(n3092), .ZN(n2933) );
  XNOR2_X1 U1223 ( .A(n1128), .B(n1127), .ZN(product_out[22]) );
  INV_X4 U1224 ( .A(n1784), .ZN(n1127) );
  INV_X4 U1226 ( .A(n1169), .ZN(n3690) );
  NOR2_X4 U1228 ( .A1(n2664), .A2(n2663), .ZN(n2544) );
  INV_X8 U1229 ( .A(n2733), .ZN(n2658) );
  INV_X4 U1230 ( .A(n3108), .ZN(n2989) );
  INV_X4 U1231 ( .A(n3496), .ZN(n3100) );
  INV_X4 U1232 ( .A(n1176), .ZN(n3095) );
  OAI21_X2 U1233 ( .B1(n3005), .B2(n1445), .A(n1176), .ZN(n3090) );
  NAND2_X1 U1234 ( .A1(n1922), .A2(n3982), .ZN(n3985) );
  XNOR2_X2 U1235 ( .A(n2847), .B(n1269), .ZN(n1129) );
  INV_X4 U1236 ( .A(n1129), .ZN(n4067) );
  CLKBUF_X3 U1237 ( .A(n3091), .Z(n1816) );
  INV_X4 U1238 ( .A(n3495), .ZN(n3101) );
  INV_X2 U1239 ( .A(n3338), .ZN(n1130) );
  NAND4_X4 U1240 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n3004)
         );
  AOI21_X2 U1242 ( .B1(n2998), .B2(n1169), .A(n2996), .ZN(n3000) );
  NAND2_X4 U1243 ( .A1(n2991), .A2(n2992), .ZN(n3002) );
  OAI211_X2 U1245 ( .C1(n3338), .C2(n1758), .A(n2003), .B(n1440), .ZN(n3339)
         );
  NAND2_X4 U1246 ( .A1(n1130), .A2(n1439), .ZN(n3104) );
  NAND2_X2 U1247 ( .A1(n3856), .A2(n1992), .ZN(n3473) );
  INV_X8 U1248 ( .A(net254949), .ZN(net255226) );
  XNOR2_X2 U1249 ( .A(n2845), .B(n1504), .ZN(n1131) );
  CLKBUF_X3 U1250 ( .A(n1958), .Z(n1972) );
  NOR2_X4 U1252 ( .A1(n1497), .A2(n3160), .ZN(n1132) );
  BUF_X4 U1253 ( .A(n3285), .Z(n1497) );
  NAND2_X4 U1254 ( .A1(n1560), .A2(n1561), .ZN(n1563) );
  INV_X4 U1255 ( .A(n3470), .ZN(n3467) );
  INV_X2 U1256 ( .A(n4102), .ZN(n1133) );
  INV_X4 U1258 ( .A(net253547), .ZN(n1568) );
  NAND2_X2 U1259 ( .A1(n1252), .A2(n1253), .ZN(n2631) );
  NAND2_X4 U1260 ( .A1(n2365), .A2(n1990), .ZN(n2335) );
  INV_X4 U1261 ( .A(net254861), .ZN(n1383) );
  NAND2_X2 U1262 ( .A1(net256953), .A2(net254673), .ZN(net254861) );
  NAND2_X4 U1263 ( .A1(n3161), .A2(n1776), .ZN(n1134) );
  XOR2_X2 U1264 ( .A(n1415), .B(n3998), .Z(n1135) );
  INV_X2 U1265 ( .A(n2584), .ZN(n1347) );
  AND2_X2 U1266 ( .A1(net256402), .A2(net255854), .ZN(n1136) );
  INV_X8 U1267 ( .A(n2447), .ZN(n2514) );
  NAND2_X2 U1268 ( .A1(a[10]), .A2(net256388), .ZN(n2447) );
  NAND2_X1 U1269 ( .A1(net256388), .A2(a[6]), .ZN(n1137) );
  INV_X8 U1270 ( .A(net256145), .ZN(net256143) );
  INV_X4 U1271 ( .A(net253246), .ZN(net256145) );
  OAI21_X4 U1272 ( .B1(n2065), .B2(n2026), .A(n2025), .ZN(n1954) );
  OR2_X2 U1273 ( .A1(n3431), .A2(n3427), .ZN(n1138) );
  NAND2_X4 U1274 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  INV_X8 U1275 ( .A(net257693), .ZN(n1258) );
  INV_X8 U1276 ( .A(n3563), .ZN(n3634) );
  INV_X2 U1277 ( .A(net255503), .ZN(net255502) );
  NAND2_X2 U1278 ( .A1(net256296), .A2(n1649), .ZN(net255503) );
  INV_X8 U1279 ( .A(n2155), .ZN(n1998) );
  INV_X8 U1280 ( .A(n2787), .ZN(n1241) );
  INV_X8 U1281 ( .A(n3597), .ZN(n1337) );
  INV_X8 U1282 ( .A(n3031), .ZN(n1479) );
  NOR2_X4 U1283 ( .A1(net254570), .A2(net254571), .ZN(net254671) );
  INV_X8 U1284 ( .A(net256582), .ZN(net256555) );
  INV_X4 U1285 ( .A(n2270), .ZN(n1804) );
  INV_X8 U1286 ( .A(n2361), .ZN(n2363) );
  INV_X8 U1287 ( .A(n2404), .ZN(n2358) );
  INV_X8 U1288 ( .A(n1705), .ZN(n1508) );
  INV_X8 U1289 ( .A(n1492), .ZN(n1707) );
  OAI21_X4 U1290 ( .B1(net254939), .B2(net254689), .A(n2811), .ZN(n1800) );
  INV_X4 U1291 ( .A(n2880), .ZN(n1303) );
  NAND2_X4 U1292 ( .A1(n1757), .A2(n2712), .ZN(n1247) );
  INV_X8 U1293 ( .A(n1679), .ZN(net257980) );
  NAND2_X4 U1294 ( .A1(n2989), .A2(n2990), .ZN(n3110) );
  INV_X4 U1295 ( .A(n3163), .ZN(n1468) );
  NAND2_X4 U1296 ( .A1(net253415), .A2(n1712), .ZN(net253422) );
  INV_X8 U1297 ( .A(n3283), .ZN(n3288) );
  INV_X8 U1298 ( .A(n3342), .ZN(n1436) );
  NAND2_X4 U1299 ( .A1(n3346), .A2(n1769), .ZN(n3534) );
  NAND2_X4 U1300 ( .A1(n3012), .A2(n3015), .ZN(n1269) );
  AOI22_X4 U1301 ( .A1(n2647), .A2(n2642), .B1(n2647), .B2(net256095), .ZN(
        n2643) );
  XOR2_X2 U1302 ( .A(n2936), .B(n3020), .Z(n1139) );
  OAI211_X2 U1303 ( .C1(n1189), .C2(net256184), .A(n4070), .B(n4069), .ZN(
        net253049) );
  NOR2_X4 U1304 ( .A1(n3494), .A2(n3781), .ZN(n1143) );
  AND2_X2 U1305 ( .A1(n1643), .A2(net253571), .ZN(n1140) );
  INV_X4 U1306 ( .A(n3497), .ZN(n3498) );
  XNOR2_X2 U1307 ( .A(n2521), .B(n1142), .ZN(n1798) );
  INV_X32 U1308 ( .A(n1794), .ZN(n1142) );
  INV_X8 U1309 ( .A(n3384), .ZN(n1540) );
  INV_X2 U1310 ( .A(n2626), .ZN(n1144) );
  NAND2_X2 U1311 ( .A1(n2391), .A2(net255498), .ZN(n1147) );
  NAND2_X4 U1312 ( .A1(n1145), .A2(n1146), .ZN(n1148) );
  NAND2_X4 U1313 ( .A1(n1147), .A2(n1148), .ZN(n2393) );
  INV_X4 U1314 ( .A(n2391), .ZN(n1145) );
  INV_X4 U1315 ( .A(net255498), .ZN(n1146) );
  NAND2_X2 U1316 ( .A1(n2721), .A2(n2720), .ZN(n1151) );
  NAND2_X4 U1317 ( .A1(n1149), .A2(n1150), .ZN(n1152) );
  NAND2_X4 U1318 ( .A1(n1151), .A2(n1152), .ZN(n2722) );
  INV_X4 U1319 ( .A(n2721), .ZN(n1149) );
  INV_X4 U1320 ( .A(n2720), .ZN(n1150) );
  NAND2_X4 U1321 ( .A1(n2392), .A2(n2393), .ZN(n2534) );
  INV_X8 U1322 ( .A(n2722), .ZN(n3007) );
  NAND2_X4 U1323 ( .A1(n1595), .A2(n1596), .ZN(n1597) );
  OAI21_X4 U1324 ( .B1(n2569), .B2(n2568), .A(n1435), .ZN(n1153) );
  NAND2_X2 U1325 ( .A1(n2403), .A2(n2404), .ZN(n1155) );
  NAND2_X4 U1326 ( .A1(n1154), .A2(n2358), .ZN(n1156) );
  NAND2_X2 U1327 ( .A1(n1155), .A2(n1156), .ZN(n2346) );
  INV_X2 U1328 ( .A(n2403), .ZN(n1154) );
  NAND2_X2 U1329 ( .A1(n2103), .A2(n2001), .ZN(n1159) );
  NAND2_X4 U1330 ( .A1(n1157), .A2(n1158), .ZN(n1160) );
  NAND2_X4 U1331 ( .A1(n1159), .A2(n1160), .ZN(n2000) );
  INV_X4 U1332 ( .A(n2103), .ZN(n1157) );
  INV_X4 U1333 ( .A(n2001), .ZN(n1158) );
  INV_X8 U1334 ( .A(n2567), .ZN(n2568) );
  NAND2_X1 U1335 ( .A1(n1390), .A2(net256165), .ZN(n2403) );
  INV_X2 U1336 ( .A(n1942), .ZN(n3190) );
  NAND2_X4 U1337 ( .A1(n1559), .A2(net253443), .ZN(n1350) );
  INV_X1 U1338 ( .A(n1991), .ZN(n1996) );
  NAND2_X4 U1339 ( .A1(n2807), .A2(n2866), .ZN(n1570) );
  INV_X4 U1340 ( .A(n2161), .ZN(n2162) );
  INV_X8 U1341 ( .A(n3385), .ZN(n3386) );
  NAND2_X4 U1342 ( .A1(n3706), .A2(net253411), .ZN(n3707) );
  INV_X8 U1343 ( .A(n2002), .ZN(n1851) );
  OAI211_X4 U1344 ( .C1(n2655), .C2(n1535), .A(n2652), .B(n2653), .ZN(n2733)
         );
  INV_X1 U1345 ( .A(net254004), .ZN(net257295) );
  INV_X4 U1346 ( .A(n1935), .ZN(n3471) );
  NAND3_X2 U1347 ( .A1(n1462), .A2(n3252), .A3(net257068), .ZN(n3389) );
  NAND3_X2 U1348 ( .A1(n3412), .A2(n1931), .A3(net257069), .ZN(n3390) );
  NOR2_X2 U1349 ( .A1(n2993), .A2(n1169), .ZN(n2994) );
  NAND2_X4 U1350 ( .A1(n3184), .A2(n3185), .ZN(n3287) );
  INV_X8 U1351 ( .A(n3334), .ZN(n1501) );
  OAI21_X2 U1352 ( .B1(n1722), .B2(net253278), .A(n1725), .ZN(n1161) );
  INV_X4 U1353 ( .A(n1746), .ZN(n1745) );
  XNOR2_X2 U1354 ( .A(n2845), .B(n1504), .ZN(n1162) );
  NAND2_X1 U1355 ( .A1(n3257), .A2(n3274), .ZN(n1165) );
  NAND2_X4 U1356 ( .A1(n1163), .A2(n1164), .ZN(n1166) );
  NAND2_X2 U1357 ( .A1(n1166), .A2(n1165), .ZN(n3258) );
  INV_X4 U1358 ( .A(n3257), .ZN(n1163) );
  INV_X8 U1360 ( .A(n3567), .ZN(n3650) );
  INV_X4 U1362 ( .A(n3621), .ZN(n1394) );
  INV_X4 U1363 ( .A(net253761), .ZN(net253652) );
  NAND2_X4 U1364 ( .A1(net253697), .A2(n1605), .ZN(n1167) );
  NAND2_X4 U1365 ( .A1(n3598), .A2(n1604), .ZN(n1605) );
  OAI22_X1 U1366 ( .A1(n2351), .A2(n3512), .B1(n4108), .B2(net256184), .ZN(
        n2929) );
  NOR2_X4 U1367 ( .A1(n3552), .A2(n3347), .ZN(n3326) );
  BUF_X4 U1368 ( .A(net253646), .Z(net258007) );
  OAI21_X4 U1369 ( .B1(n3288), .B2(n1910), .A(n3286), .ZN(n1168) );
  NAND2_X2 U1370 ( .A1(n1851), .A2(n3110), .ZN(n1169) );
  NAND2_X2 U1371 ( .A1(n1851), .A2(n3110), .ZN(n2997) );
  INV_X8 U1372 ( .A(n3587), .ZN(n3639) );
  INV_X8 U1373 ( .A(n4000), .ZN(n4002) );
  NAND2_X2 U1374 ( .A1(n3611), .A2(n3612), .ZN(n1172) );
  NAND2_X2 U1375 ( .A1(n1170), .A2(n1171), .ZN(n1173) );
  NAND2_X2 U1376 ( .A1(n1172), .A2(n1173), .ZN(net253808) );
  INV_X4 U1377 ( .A(n3611), .ZN(n1170) );
  INV_X4 U1378 ( .A(n3612), .ZN(n1171) );
  INV_X4 U1379 ( .A(n1980), .ZN(n1981) );
  NAND2_X4 U1380 ( .A1(n3004), .A2(n1418), .ZN(n1176) );
  NAND2_X2 U1381 ( .A1(n1174), .A2(n1175), .ZN(n1177) );
  NAND2_X2 U1382 ( .A1(n1176), .A2(n1177), .ZN(n1941) );
  INV_X4 U1383 ( .A(n1418), .ZN(n1175) );
  NAND2_X2 U1384 ( .A1(n1941), .A2(n1176), .ZN(n3495) );
  NAND2_X4 U1385 ( .A1(n3476), .A2(n4107), .ZN(n3257) );
  INV_X4 U1387 ( .A(net253273), .ZN(net256839) );
  NAND2_X2 U1388 ( .A1(n3379), .A2(n1179), .ZN(n1180) );
  NAND2_X2 U1389 ( .A1(n1178), .A2(n1765), .ZN(n1181) );
  NAND2_X2 U1390 ( .A1(n1180), .A2(n1181), .ZN(n1809) );
  INV_X1 U1391 ( .A(n3379), .ZN(n1178) );
  INV_X4 U1392 ( .A(n1765), .ZN(n1179) );
  XNOR2_X2 U1393 ( .A(n3431), .B(n3314), .ZN(n1182) );
  NAND2_X4 U1394 ( .A1(n3312), .A2(n3313), .ZN(n3314) );
  NAND2_X2 U1396 ( .A1(net255626), .A2(n1258), .ZN(net255591) );
  INV_X4 U1397 ( .A(n1882), .ZN(n1329) );
  INV_X8 U1398 ( .A(n2502), .ZN(n1873) );
  NAND2_X4 U1399 ( .A1(n2841), .A2(n1773), .ZN(n2941) );
  INV_X1 U1400 ( .A(n3494), .ZN(n1183) );
  NAND2_X1 U1401 ( .A1(n2840), .A2(net254856), .ZN(n1186) );
  NAND2_X4 U1402 ( .A1(n1184), .A2(n1185), .ZN(n1187) );
  NAND2_X2 U1403 ( .A1(n1186), .A2(n1187), .ZN(n2842) );
  INV_X4 U1404 ( .A(n2840), .ZN(n1184) );
  XNOR2_X2 U1406 ( .A(n1137), .B(n2436), .ZN(n1822) );
  NAND2_X4 U1407 ( .A1(n2868), .A2(n2869), .ZN(n1455) );
  INV_X4 U1408 ( .A(net253586), .ZN(n1675) );
  NAND2_X2 U1409 ( .A1(n3458), .A2(n3459), .ZN(n3549) );
  INV_X8 U1410 ( .A(n2443), .ZN(n2586) );
  INV_X2 U1411 ( .A(net257439), .ZN(net253984) );
  NAND2_X4 U1412 ( .A1(n3319), .A2(n3320), .ZN(n1544) );
  XNOR2_X2 U1413 ( .A(n2274), .B(n2263), .ZN(n1188) );
  NAND2_X2 U1414 ( .A1(n2062), .A2(n2063), .ZN(n2064) );
  NAND2_X4 U1415 ( .A1(n3665), .A2(n3718), .ZN(n3719) );
  INV_X2 U1416 ( .A(n3675), .ZN(n3673) );
  NAND3_X2 U1417 ( .A1(n2580), .A2(n2676), .A3(n2579), .ZN(n2581) );
  BUF_X8 U1418 ( .A(net254291), .Z(net257254) );
  INV_X2 U1419 ( .A(n2895), .ZN(n1814) );
  INV_X2 U1420 ( .A(n2830), .ZN(n2758) );
  XNOR2_X2 U1421 ( .A(n3396), .B(n1190), .ZN(n1189) );
  NAND2_X4 U1423 ( .A1(net254084), .A2(net254052), .ZN(net254051) );
  INV_X2 U1424 ( .A(n2385), .ZN(n1346) );
  INV_X1 U1425 ( .A(n2699), .ZN(n2454) );
  NAND2_X2 U1426 ( .A1(n3466), .A2(n1212), .ZN(n1193) );
  NAND2_X4 U1427 ( .A1(n1191), .A2(n1192), .ZN(n1194) );
  NAND2_X4 U1428 ( .A1(n1193), .A2(n1194), .ZN(n3470) );
  INV_X4 U1429 ( .A(n3466), .ZN(n1191) );
  INV_X4 U1430 ( .A(n1212), .ZN(n1192) );
  AND2_X2 U1431 ( .A1(net253647), .A2(net253646), .ZN(n1212) );
  INV_X1 U1432 ( .A(net255107), .ZN(net255102) );
  OAI21_X2 U1433 ( .B1(n1804), .B2(n2218), .A(n2315), .ZN(n2279) );
  NAND3_X2 U1434 ( .A1(n1113), .A2(n3540), .A3(n3541), .ZN(n1195) );
  NAND2_X2 U1435 ( .A1(n2514), .A2(n2513), .ZN(n1197) );
  NAND2_X4 U1436 ( .A1(n2447), .A2(n1196), .ZN(n1198) );
  NAND2_X4 U1437 ( .A1(n1197), .A2(n1198), .ZN(n2594) );
  INV_X8 U1438 ( .A(n2513), .ZN(n1196) );
  NAND2_X1 U1439 ( .A1(n3981), .A2(n3980), .ZN(n1200) );
  NAND2_X4 U1440 ( .A1(n1135), .A2(n1199), .ZN(n1201) );
  NAND2_X4 U1441 ( .A1(n1200), .A2(n1201), .ZN(net253057) );
  INV_X4 U1442 ( .A(n3980), .ZN(n1199) );
  INV_X4 U1443 ( .A(net253057), .ZN(net253209) );
  NAND2_X1 U1444 ( .A1(net254687), .A2(net254688), .ZN(n2958) );
  INV_X16 U1445 ( .A(control[0]), .ZN(net257677) );
  INV_X16 U1446 ( .A(control[0]), .ZN(n1357) );
  INV_X16 U1447 ( .A(control[0]), .ZN(n1358) );
  INV_X16 U1448 ( .A(control[0]), .ZN(n1221) );
  INV_X16 U1449 ( .A(control[0]), .ZN(n1222) );
  INV_X8 U1450 ( .A(n2323), .ZN(n2205) );
  INV_X32 U1451 ( .A(control[1]), .ZN(net257720) );
  NAND2_X2 U1452 ( .A1(net254180), .A2(net254181), .ZN(net254057) );
  INV_X8 U1453 ( .A(net253270), .ZN(net253388) );
  CLKBUF_X2 U1454 ( .A(n3141), .Z(n1202) );
  NAND2_X4 U1455 ( .A1(n3545), .A2(n3551), .ZN(n3452) );
  OAI21_X4 U1456 ( .B1(n3445), .B2(n3446), .A(n3448), .ZN(n3545) );
  INV_X4 U1457 ( .A(n2842), .ZN(n2843) );
  INV_X4 U1458 ( .A(n3849), .ZN(n3863) );
  AOI21_X2 U1459 ( .B1(n2670), .B2(n4110), .A(n1260), .ZN(n2672) );
  INV_X8 U1460 ( .A(n2669), .ZN(n2947) );
  NAND2_X4 U1461 ( .A1(n1203), .A2(n1204), .ZN(n1205) );
  NAND2_X4 U1462 ( .A1(n1205), .A2(n2028), .ZN(n2093) );
  INV_X4 U1463 ( .A(n2030), .ZN(n1203) );
  INV_X4 U1464 ( .A(n2029), .ZN(n1204) );
  NAND2_X4 U1465 ( .A1(a[2]), .A2(net257678), .ZN(n2030) );
  INV_X4 U1466 ( .A(n2093), .ZN(n2098) );
  CLKBUF_X3 U1467 ( .A(n3198), .Z(n1206) );
  INV_X4 U1468 ( .A(n1733), .ZN(net256958) );
  INV_X4 U1469 ( .A(net255226), .ZN(net256860) );
  NOR2_X2 U1470 ( .A1(net255592), .A2(net255438), .ZN(net255588) );
  NAND2_X4 U1471 ( .A1(b[16]), .A2(control[0]), .ZN(n1207) );
  INV_X4 U1472 ( .A(n2954), .ZN(n1584) );
  NAND2_X4 U1473 ( .A1(n1798), .A2(n2522), .ZN(n2525) );
  INV_X8 U1474 ( .A(n1939), .ZN(n1513) );
  NAND2_X2 U1475 ( .A1(n4012), .A2(n4011), .ZN(n3969) );
  NAND3_X4 U1476 ( .A1(n3976), .A2(n1917), .A3(n3974), .ZN(n4000) );
  INV_X8 U1477 ( .A(n3973), .ZN(n3974) );
  NOR2_X4 U1478 ( .A1(n3858), .A2(n3857), .ZN(n1262) );
  OAI21_X4 U1479 ( .B1(net257239), .B2(net254306), .A(n1668), .ZN(net254297)
         );
  NOR2_X4 U1480 ( .A1(n3690), .A2(net256095), .ZN(n2991) );
  INV_X8 U1481 ( .A(n1855), .ZN(n2790) );
  INV_X4 U1482 ( .A(n1748), .ZN(n1747) );
  NAND2_X1 U1483 ( .A1(n3991), .A2(n1973), .ZN(n1210) );
  NAND2_X4 U1484 ( .A1(n1208), .A2(n1209), .ZN(n1211) );
  NAND2_X2 U1485 ( .A1(n1210), .A2(n1211), .ZN(product_out[30]) );
  INV_X4 U1486 ( .A(n3991), .ZN(n1208) );
  INV_X4 U1487 ( .A(n1973), .ZN(n1209) );
  NAND2_X2 U1488 ( .A1(n1587), .A2(n1241), .ZN(n1243) );
  NAND2_X1 U1489 ( .A1(n2135), .A2(n2134), .ZN(n2138) );
  INV_X2 U1491 ( .A(n2109), .ZN(n1551) );
  NAND2_X4 U1492 ( .A1(n2151), .A2(n2187), .ZN(n2226) );
  INV_X2 U1493 ( .A(n2082), .ZN(n1572) );
  NAND2_X4 U1494 ( .A1(n2266), .A2(n2265), .ZN(n2267) );
  NAND2_X4 U1495 ( .A1(n2191), .A2(n2190), .ZN(n2140) );
  NAND3_X1 U1496 ( .A1(net257044), .A2(net253058), .A3(net253059), .ZN(
        net253056) );
  NAND3_X1 U1497 ( .A1(net253058), .A2(net253208), .A3(net253059), .ZN(
        net257661) );
  NAND2_X1 U1498 ( .A1(n3860), .A2(net253173), .ZN(n1215) );
  NAND2_X2 U1499 ( .A1(n1213), .A2(n1214), .ZN(n1216) );
  NAND2_X2 U1500 ( .A1(n1215), .A2(n1216), .ZN(n3927) );
  INV_X2 U1501 ( .A(n3860), .ZN(n1213) );
  INV_X1 U1502 ( .A(net253173), .ZN(n1214) );
  NAND2_X4 U1503 ( .A1(product_in[28]), .A2(net256095), .ZN(net253173) );
  NAND2_X1 U1504 ( .A1(n2230), .A2(n2268), .ZN(n2165) );
  AOI21_X2 U1505 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3946) );
  NAND2_X2 U1506 ( .A1(n3940), .A2(n1833), .ZN(n3943) );
  NAND2_X4 U1507 ( .A1(n1136), .A2(net255856), .ZN(net255852) );
  INV_X16 U1508 ( .A(net256401), .ZN(net256402) );
  INV_X1 U1509 ( .A(net255868), .ZN(net255854) );
  INV_X32 U1510 ( .A(control[1]), .ZN(net256077) );
  NAND2_X2 U1511 ( .A1(n1248), .A2(net255040), .ZN(n1219) );
  NAND2_X4 U1512 ( .A1(n1217), .A2(n1218), .ZN(n1220) );
  NAND2_X4 U1513 ( .A1(n1220), .A2(n1219), .ZN(n2713) );
  INV_X8 U1516 ( .A(n2713), .ZN(n2714) );
  OAI21_X4 U1517 ( .B1(n1463), .B2(n1464), .A(n3383), .ZN(n1542) );
  OAI221_X4 U1518 ( .B1(net256800), .B2(n1471), .C1(n1262), .C2(net253422), 
        .A(net257435), .ZN(net253405) );
  INV_X8 U1519 ( .A(n1896), .ZN(n1260) );
  NAND4_X4 U1520 ( .A1(b[25]), .A2(net257782), .A3(a[0]), .A4(net256087), .ZN(
        n2015) );
  INV_X4 U1521 ( .A(n2041), .ZN(n1363) );
  NAND2_X2 U1522 ( .A1(net253806), .A2(net253804), .ZN(net253776) );
  INV_X2 U1523 ( .A(n2080), .ZN(n1761) );
  INV_X4 U1524 ( .A(n2555), .ZN(n2556) );
  NAND2_X4 U1525 ( .A1(n1348), .A2(n1349), .ZN(n2387) );
  INV_X4 U1526 ( .A(net253659), .ZN(net253657) );
  INV_X4 U1527 ( .A(n1811), .ZN(n2662) );
  AOI211_X4 U1528 ( .C1(net253182), .C2(net253183), .A(n1716), .B(net253185), 
        .ZN(n1715) );
  INV_X4 U1529 ( .A(n2623), .ZN(n2624) );
  INV_X4 U1530 ( .A(n2716), .ZN(n1263) );
  INV_X4 U1531 ( .A(n3851), .ZN(n1472) );
  NAND2_X2 U1532 ( .A1(n2390), .A2(n1819), .ZN(n1225) );
  NAND2_X4 U1533 ( .A1(n1223), .A2(n1224), .ZN(n1226) );
  NAND2_X4 U1534 ( .A1(n1225), .A2(n1226), .ZN(net255504) );
  INV_X4 U1535 ( .A(n2390), .ZN(n1223) );
  INV_X4 U1536 ( .A(n1819), .ZN(n1224) );
  INV_X8 U1537 ( .A(net255504), .ZN(net255507) );
  INV_X8 U1538 ( .A(n3714), .ZN(n3716) );
  INV_X4 U1539 ( .A(n1458), .ZN(n1227) );
  INV_X1 U1540 ( .A(n1458), .ZN(net255878) );
  INV_X2 U1541 ( .A(n3755), .ZN(n1921) );
  INV_X8 U1542 ( .A(n3595), .ZN(n3685) );
  NAND2_X4 U1543 ( .A1(n1338), .A2(n1339), .ZN(n3595) );
  NAND3_X1 U1544 ( .A1(n2116), .A2(n2370), .A3(net255910), .ZN(n2112) );
  NAND2_X2 U1545 ( .A1(n1120), .A2(n3393), .ZN(n1230) );
  NAND2_X4 U1546 ( .A1(n1228), .A2(n1229), .ZN(n1231) );
  NAND2_X4 U1547 ( .A1(n1230), .A2(n1231), .ZN(n1935) );
  INV_X4 U1548 ( .A(n3394), .ZN(n1228) );
  INV_X4 U1549 ( .A(n3393), .ZN(n1229) );
  NAND2_X2 U1550 ( .A1(n2521), .A2(n1794), .ZN(n1276) );
  NAND2_X4 U1551 ( .A1(n1276), .A2(n1277), .ZN(n2523) );
  NOR2_X1 U1552 ( .A1(n2111), .A2(net257772), .ZN(n2109) );
  NAND2_X4 U1553 ( .A1(net256054), .A2(net256055), .ZN(n1232) );
  INV_X32 U1554 ( .A(net257585), .ZN(net257586) );
  INV_X2 U1555 ( .A(net256145), .ZN(net256141) );
  INV_X16 U1556 ( .A(net255721), .ZN(n1460) );
  INV_X1 U1557 ( .A(net257586), .ZN(net255721) );
  NAND2_X2 U1558 ( .A1(n1161), .A2(net253315), .ZN(n1235) );
  NAND2_X4 U1559 ( .A1(n1233), .A2(n1234), .ZN(n1236) );
  NAND2_X4 U1560 ( .A1(n1235), .A2(n1236), .ZN(net253305) );
  INV_X4 U1561 ( .A(net253315), .ZN(n1233) );
  INV_X4 U1562 ( .A(net253316), .ZN(n1234) );
  NAND2_X4 U1563 ( .A1(net256054), .A2(net256055), .ZN(net253246) );
  AOI21_X4 U1564 ( .B1(net253405), .B2(n1442), .A(net253206), .ZN(net253315)
         );
  NAND2_X2 U1565 ( .A1(n2257), .A2(net255705), .ZN(n1239) );
  NAND2_X4 U1566 ( .A1(n1237), .A2(n1238), .ZN(n1240) );
  NAND2_X4 U1567 ( .A1(n1239), .A2(n1240), .ZN(net255702) );
  INV_X4 U1568 ( .A(n2257), .ZN(n1237) );
  INV_X4 U1569 ( .A(net255705), .ZN(n1238) );
  NAND2_X2 U1570 ( .A1(net255427), .A2(net255618), .ZN(net255705) );
  NAND2_X4 U1571 ( .A1(net255702), .A2(net255703), .ZN(net255629) );
  INV_X4 U1572 ( .A(net257296), .ZN(net254306) );
  NAND2_X4 U1573 ( .A1(n1587), .A2(n1241), .ZN(n1589) );
  NAND2_X1 U1574 ( .A1(n2787), .A2(n1800), .ZN(n1242) );
  NAND2_X2 U1575 ( .A1(n1242), .A2(n1243), .ZN(n1946) );
  XNOR2_X2 U1576 ( .A(n3744), .B(n3743), .ZN(n1244) );
  NAND2_X1 U1577 ( .A1(a[23]), .A2(net256125), .ZN(n1245) );
  NAND2_X4 U1578 ( .A1(n1246), .A2(n3747), .ZN(n3939) );
  INV_X4 U1579 ( .A(n1245), .ZN(n1246) );
  NAND2_X4 U1580 ( .A1(n3838), .A2(n3839), .ZN(n3743) );
  INV_X4 U1581 ( .A(n3939), .ZN(n3898) );
  XNOR2_X2 U1582 ( .A(net255040), .B(n1248), .ZN(n1757) );
  NAND2_X4 U1583 ( .A1(n1117), .A2(n2527), .ZN(n2674) );
  NAND4_X2 U1584 ( .A1(b[1]), .A2(control[1]), .A3(a[4]), .A4(control[0]), 
        .ZN(n2100) );
  INV_X4 U1585 ( .A(n1697), .ZN(net256874) );
  INV_X4 U1586 ( .A(net253810), .ZN(n1397) );
  INV_X2 U1587 ( .A(net254695), .ZN(net257266) );
  INV_X8 U1588 ( .A(n2854), .ZN(n2855) );
  INV_X4 U1589 ( .A(n2338), .ZN(n2336) );
  INV_X8 U1590 ( .A(n1506), .ZN(net255324) );
  NAND2_X4 U1591 ( .A1(n2332), .A2(n2331), .ZN(n2334) );
  NAND2_X4 U1592 ( .A1(n3154), .A2(net254411), .ZN(n1477) );
  INV_X8 U1593 ( .A(net254188), .ZN(n1296) );
  NAND2_X4 U1594 ( .A1(n1752), .A2(n1751), .ZN(n1443) );
  NAND2_X2 U1595 ( .A1(n2714), .A2(n2715), .ZN(n1278) );
  NAND2_X4 U1596 ( .A1(n1273), .A2(n2738), .ZN(n2635) );
  INV_X4 U1597 ( .A(n2630), .ZN(n2538) );
  INV_X1 U1598 ( .A(net255548), .ZN(n1249) );
  NAND2_X4 U1599 ( .A1(n3411), .A2(n3412), .ZN(net253797) );
  BUF_X4 U1600 ( .A(net253764), .Z(n1721) );
  NAND2_X4 U1601 ( .A1(net254577), .A2(net254367), .ZN(net254576) );
  NAND3_X4 U1602 ( .A1(n1441), .A2(a[12]), .A3(net256173), .ZN(n3185) );
  NAND2_X4 U1603 ( .A1(n3020), .A2(n1895), .ZN(n3021) );
  NAND2_X2 U1604 ( .A1(net255324), .A2(net255107), .ZN(net256627) );
  NAND2_X2 U1605 ( .A1(n3798), .A2(net253519), .ZN(n3803) );
  INV_X8 U1606 ( .A(n3606), .ZN(n3681) );
  INV_X4 U1607 ( .A(n2952), .ZN(n1904) );
  NAND2_X1 U1608 ( .A1(n1319), .A2(n1916), .ZN(n1252) );
  NAND2_X4 U1609 ( .A1(n1250), .A2(n1251), .ZN(n1253) );
  INV_X4 U1610 ( .A(n1319), .ZN(n1250) );
  INV_X2 U1611 ( .A(n1916), .ZN(n1251) );
  INV_X4 U1612 ( .A(n2671), .ZN(n1319) );
  NAND2_X4 U1613 ( .A1(n2631), .A2(n2632), .ZN(n1273) );
  INV_X4 U1614 ( .A(n2881), .ZN(n2954) );
  INV_X4 U1615 ( .A(n2809), .ZN(n2810) );
  INV_X8 U1616 ( .A(net254696), .ZN(n1585) );
  NAND2_X2 U1617 ( .A1(net254577), .A2(net254364), .ZN(n3112) );
  OAI21_X4 U1618 ( .B1(net254468), .B2(n3112), .A(n3190), .ZN(n3154) );
  NAND2_X4 U1619 ( .A1(n3116), .A2(n2974), .ZN(n3207) );
  AOI21_X4 U1621 ( .B1(net254189), .B2(n1666), .A(net254191), .ZN(net254188)
         );
  NAND2_X1 U1622 ( .A1(net255502), .A2(net255501), .ZN(n1380) );
  NAND2_X4 U1623 ( .A1(n1553), .A2(n1835), .ZN(n2147) );
  NAND2_X4 U1624 ( .A1(n2146), .A2(n2147), .ZN(n2194) );
  NAND2_X2 U1625 ( .A1(net254142), .A2(n1632), .ZN(net254182) );
  INV_X2 U1626 ( .A(n1584), .ZN(n1453) );
  NAND2_X4 U1627 ( .A1(n2233), .A2(n2232), .ZN(n2308) );
  INV_X2 U1628 ( .A(n2234), .ZN(n2235) );
  NAND2_X2 U1629 ( .A1(net254183), .A2(net254182), .ZN(n1256) );
  NAND2_X4 U1630 ( .A1(n1254), .A2(n1255), .ZN(n1257) );
  NAND2_X4 U1631 ( .A1(n1257), .A2(n1256), .ZN(net254180) );
  INV_X4 U1632 ( .A(net254183), .ZN(n1255) );
  INV_X4 U1633 ( .A(n2504), .ZN(n2611) );
  AND2_X4 U1634 ( .A1(net257485), .A2(net257240), .ZN(n1430) );
  NAND2_X2 U1635 ( .A1(n1379), .A2(net255503), .ZN(n1381) );
  NAND2_X2 U1636 ( .A1(n1259), .A2(net254751), .ZN(net256974) );
  NAND2_X4 U1637 ( .A1(n2811), .A2(n1882), .ZN(n2787) );
  INV_X2 U1638 ( .A(net253690), .ZN(n1509) );
  INV_X2 U1639 ( .A(n1585), .ZN(n1483) );
  INV_X32 U1640 ( .A(control[1]), .ZN(net257721) );
  INV_X32 U1641 ( .A(control[1]), .ZN(n1466) );
  NAND2_X4 U1642 ( .A1(n3062), .A2(n3191), .ZN(n3138) );
  INV_X8 U1643 ( .A(n1324), .ZN(n2425) );
  INV_X4 U1644 ( .A(n1260), .ZN(n1261) );
  INV_X4 U1645 ( .A(n2213), .ZN(n2211) );
  INV_X2 U1646 ( .A(n1945), .ZN(n3759) );
  OAI21_X2 U1647 ( .B1(net253380), .B2(n3865), .A(n3934), .ZN(n3908) );
  NAND2_X1 U1648 ( .A1(n2758), .A2(n2890), .ZN(n2764) );
  INV_X4 U1649 ( .A(n2579), .ZN(n2753) );
  NAND2_X4 U1650 ( .A1(net254242), .A2(net254285), .ZN(net254147) );
  NAND2_X2 U1651 ( .A1(net256375), .A2(n3628), .ZN(n1538) );
  INV_X4 U1652 ( .A(n2347), .ZN(n2350) );
  NAND2_X4 U1653 ( .A1(n2277), .A2(n1763), .ZN(n2360) );
  XNOR2_X2 U1654 ( .A(n2275), .B(n2274), .ZN(n1763) );
  NAND2_X4 U1655 ( .A1(n2421), .A2(n2305), .ZN(n2294) );
  NAND2_X2 U1656 ( .A1(n2716), .A2(n1318), .ZN(n1265) );
  NAND2_X4 U1657 ( .A1(n1263), .A2(n1264), .ZN(n1266) );
  NAND2_X4 U1658 ( .A1(n1265), .A2(n1266), .ZN(n2719) );
  INV_X4 U1659 ( .A(n1318), .ZN(n1264) );
  NAND2_X2 U1660 ( .A1(n3267), .A2(n3171), .ZN(n1581) );
  INV_X2 U1661 ( .A(n2949), .ZN(n1318) );
  NAND3_X4 U1662 ( .A1(n2719), .A2(a[8]), .A3(net256173), .ZN(n2871) );
  NAND2_X4 U1663 ( .A1(net253657), .A2(net253656), .ZN(n1471) );
  NOR2_X4 U1664 ( .A1(n3428), .A2(n1138), .ZN(n3435) );
  NAND2_X4 U1665 ( .A1(n3234), .A2(n3430), .ZN(n3427) );
  NOR3_X4 U1666 ( .A1(net255413), .A2(n1411), .A3(n2586), .ZN(n2440) );
  INV_X8 U1667 ( .A(n3538), .ZN(n3539) );
  INV_X4 U1669 ( .A(n2997), .ZN(n1267) );
  OAI21_X4 U1670 ( .B1(n2328), .B2(n2327), .A(n2326), .ZN(n2333) );
  NAND2_X1 U1671 ( .A1(n2090), .A2(n2164), .ZN(net254390) );
  NAND2_X4 U1672 ( .A1(n1599), .A2(n1600), .ZN(n1602) );
  NAND2_X4 U1673 ( .A1(n1303), .A2(n1483), .ZN(n2883) );
  INV_X8 U1674 ( .A(net254684), .ZN(net254681) );
  BUF_X32 U1675 ( .A(n1839), .Z(n1268) );
  NAND2_X4 U1676 ( .A1(n1602), .A2(n1601), .ZN(n2623) );
  INV_X4 U1677 ( .A(net254711), .ZN(n1270) );
  INV_X4 U1678 ( .A(net254711), .ZN(net254695) );
  NOR2_X2 U1679 ( .A1(n1678), .A2(net253643), .ZN(n1674) );
  NAND2_X2 U1680 ( .A1(n2886), .A2(n2890), .ZN(n2007) );
  NAND2_X4 U1681 ( .A1(n3519), .A2(n3520), .ZN(n1271) );
  INV_X4 U1683 ( .A(n1271), .ZN(n1272) );
  NAND2_X4 U1684 ( .A1(n3080), .A2(n3081), .ZN(n3519) );
  INV_X8 U1685 ( .A(n2846), .ZN(n2847) );
  INV_X8 U1686 ( .A(n2516), .ZN(n2584) );
  NAND2_X4 U1687 ( .A1(n1499), .A2(n1500), .ZN(n1886) );
  NAND2_X4 U1688 ( .A1(n2874), .A2(n1498), .ZN(n1500) );
  NAND2_X4 U1689 ( .A1(n1274), .A2(n1275), .ZN(n1277) );
  INV_X4 U1690 ( .A(n2521), .ZN(n1274) );
  INV_X2 U1691 ( .A(n1794), .ZN(n1275) );
  NAND2_X4 U1692 ( .A1(n2592), .A2(n1285), .ZN(n1794) );
  INV_X8 U1693 ( .A(n2461), .ZN(n2462) );
  NAND4_X4 U1694 ( .A1(n2459), .A2(n2458), .A3(n2457), .A4(n2456), .ZN(n2461)
         );
  INV_X8 U1695 ( .A(net255332), .ZN(net255500) );
  INV_X4 U1696 ( .A(n3995), .ZN(n1554) );
  INV_X4 U1697 ( .A(n3351), .ZN(n1464) );
  INV_X4 U1698 ( .A(n1953), .ZN(n1279) );
  NAND2_X1 U1699 ( .A1(n1132), .A2(n3163), .ZN(n1281) );
  NAND2_X4 U1700 ( .A1(n1468), .A2(n1280), .ZN(n1282) );
  NAND2_X4 U1701 ( .A1(n1281), .A2(n1282), .ZN(n3166) );
  INV_X4 U1702 ( .A(n3164), .ZN(n1280) );
  OAI21_X4 U1703 ( .B1(net255429), .B2(net255428), .A(net255430), .ZN(n1953)
         );
  NAND2_X2 U1705 ( .A1(n2445), .A2(n1822), .ZN(n2254) );
  NAND2_X2 U1706 ( .A1(n1545), .A2(net253776), .ZN(n1283) );
  NAND3_X2 U1707 ( .A1(net253775), .A2(net253646), .A3(n1284), .ZN(net253772)
         );
  INV_X4 U1708 ( .A(n1283), .ZN(n1284) );
  NAND2_X2 U1709 ( .A1(net253772), .A2(n3614), .ZN(n3631) );
  INV_X4 U1710 ( .A(n3988), .ZN(n3987) );
  NAND2_X2 U1711 ( .A1(n1295), .A2(net254184), .ZN(net254050) );
  OAI21_X4 U1712 ( .B1(net256145), .B2(n2511), .A(n2590), .ZN(n1285) );
  NAND2_X2 U1713 ( .A1(net254284), .A2(net254239), .ZN(n1288) );
  NAND2_X4 U1714 ( .A1(n1286), .A2(n1287), .ZN(n1289) );
  NAND2_X4 U1715 ( .A1(n1288), .A2(n1289), .ZN(net254255) );
  INV_X1 U1716 ( .A(net254239), .ZN(n1287) );
  NAND2_X4 U1717 ( .A1(net254361), .A2(n1105), .ZN(net254284) );
  INV_X2 U1718 ( .A(net254255), .ZN(net254283) );
  NAND2_X2 U1719 ( .A1(net253449), .A2(net253450), .ZN(n1290) );
  INV_X8 U1720 ( .A(n3324), .ZN(n1291) );
  INV_X2 U1721 ( .A(n3049), .ZN(n2904) );
  OAI21_X4 U1722 ( .B1(n3042), .B2(n1928), .A(n3040), .ZN(n3119) );
  NAND2_X2 U1723 ( .A1(n2141), .A2(n2076), .ZN(n2077) );
  NAND2_X2 U1724 ( .A1(n2461), .A2(n2460), .ZN(n2464) );
  INV_X4 U1725 ( .A(n1291), .ZN(n1292) );
  AOI21_X2 U1726 ( .B1(n3325), .B2(n3455), .A(n3456), .ZN(net254189) );
  NAND2_X2 U1727 ( .A1(n3353), .A2(n1936), .ZN(n1293) );
  NAND3_X2 U1728 ( .A1(n2400), .A2(a[3]), .A3(net256165), .ZN(n2555) );
  INV_X2 U1729 ( .A(n2400), .ZN(n2399) );
  NAND2_X1 U1730 ( .A1(a[17]), .A2(net256105), .ZN(n1294) );
  INV_X4 U1731 ( .A(n1294), .ZN(n1295) );
  NAND2_X2 U1732 ( .A1(net254188), .A2(n3326), .ZN(n1298) );
  NAND2_X4 U1733 ( .A1(n1296), .A2(n1297), .ZN(n1299) );
  NAND2_X4 U1734 ( .A1(n1298), .A2(n1299), .ZN(net254184) );
  INV_X4 U1735 ( .A(n3326), .ZN(n1297) );
  INV_X4 U1736 ( .A(net256362), .ZN(net254084) );
  BUF_X8 U1737 ( .A(net255914), .Z(net257401) );
  INV_X4 U1738 ( .A(n1131), .ZN(n1994) );
  OAI21_X4 U1739 ( .B1(n3111), .B2(n1852), .A(n1799), .ZN(n1300) );
  INV_X8 U1740 ( .A(n2873), .ZN(n1301) );
  NAND2_X1 U1741 ( .A1(n2789), .A2(n2880), .ZN(n1304) );
  NAND2_X4 U1742 ( .A1(n1302), .A2(n1303), .ZN(n1305) );
  NAND2_X4 U1743 ( .A1(n1304), .A2(n1305), .ZN(n1855) );
  INV_X4 U1744 ( .A(n2789), .ZN(n1302) );
  INV_X8 U1745 ( .A(n3179), .ZN(n2873) );
  NAND3_X1 U1746 ( .A1(n2688), .A2(n2687), .A3(n2686), .ZN(n2689) );
  INV_X8 U1747 ( .A(net255431), .ZN(net255430) );
  XNOR2_X2 U1748 ( .A(n2385), .B(n1347), .ZN(n1306) );
  INV_X8 U1749 ( .A(n2690), .ZN(n2696) );
  NAND2_X1 U1750 ( .A1(n2612), .A2(n2465), .ZN(n1309) );
  NAND2_X4 U1751 ( .A1(n1307), .A2(n1308), .ZN(n1310) );
  NAND2_X4 U1752 ( .A1(n1309), .A2(n1310), .ZN(net255225) );
  INV_X4 U1753 ( .A(n2465), .ZN(n1307) );
  INV_X1 U1754 ( .A(n2612), .ZN(n1308) );
  NAND2_X4 U1755 ( .A1(n1377), .A2(n1378), .ZN(n2920) );
  INV_X4 U1756 ( .A(n2040), .ZN(n1387) );
  NAND2_X2 U1757 ( .A1(n3334), .A2(n3333), .ZN(n1312) );
  NAND2_X4 U1758 ( .A1(n1501), .A2(n1311), .ZN(n1313) );
  NAND2_X4 U1759 ( .A1(n1313), .A2(n1312), .ZN(n1943) );
  INV_X4 U1760 ( .A(n3333), .ZN(n1311) );
  AOI22_X2 U1761 ( .A1(n3856), .A2(n3475), .B1(n3477), .B2(n1850), .ZN(n3479)
         );
  INV_X2 U1762 ( .A(net255047), .ZN(n1485) );
  OAI22_X2 U1763 ( .A1(net256099), .A2(n2864), .B1(n3405), .B2(n2864), .ZN(
        n2849) );
  NAND3_X2 U1764 ( .A1(net256402), .A2(net256527), .A3(n1840), .ZN(n2203) );
  OAI21_X4 U1765 ( .B1(n2184), .B2(n2183), .A(n1444), .ZN(n2125) );
  NAND2_X4 U1766 ( .A1(n2124), .A2(n2157), .ZN(n2265) );
  NAND2_X1 U1767 ( .A1(n1669), .A2(n1666), .ZN(n1315) );
  NAND2_X4 U1768 ( .A1(n1314), .A2(net254192), .ZN(n1316) );
  NAND2_X2 U1769 ( .A1(n1315), .A2(n1316), .ZN(n1670) );
  INV_X4 U1770 ( .A(n1669), .ZN(n1314) );
  OAI21_X4 U1771 ( .B1(n3246), .B2(n3323), .A(n3245), .ZN(n1317) );
  NAND2_X2 U1772 ( .A1(n3340), .A2(n3334), .ZN(n1502) );
  NAND2_X4 U1773 ( .A1(n2744), .A2(n2745), .ZN(n2671) );
  INV_X8 U1774 ( .A(n2072), .ZN(n1792) );
  NAND2_X4 U1775 ( .A1(net255507), .A2(net255506), .ZN(n2500) );
  NAND2_X2 U1776 ( .A1(n2749), .A2(n2748), .ZN(n2676) );
  NOR2_X2 U1777 ( .A1(n2184), .A2(n2183), .ZN(n2160) );
  INV_X4 U1778 ( .A(n2091), .ZN(n2184) );
  OAI21_X1 U1779 ( .B1(n3544), .B2(n3543), .A(n3702), .ZN(n3616) );
  INV_X2 U1780 ( .A(n3702), .ZN(n3703) );
  NAND2_X2 U1781 ( .A1(net254297), .A2(n1321), .ZN(n1322) );
  NAND2_X1 U1782 ( .A1(n1320), .A2(net254298), .ZN(n1323) );
  NAND2_X2 U1783 ( .A1(n1322), .A2(n1323), .ZN(net256947) );
  INV_X1 U1784 ( .A(net254297), .ZN(n1320) );
  INV_X1 U1785 ( .A(net254298), .ZN(n1321) );
  NAND2_X4 U1789 ( .A1(n2261), .A2(n2262), .ZN(n1324) );
  NAND2_X2 U1790 ( .A1(n2261), .A2(n2262), .ZN(n2424) );
  NOR2_X4 U1791 ( .A1(n1326), .A2(control[0]), .ZN(n1325) );
  INV_X32 U1792 ( .A(a[3]), .ZN(n1326) );
  NOR2_X4 U1793 ( .A1(n2502), .A2(net255179), .ZN(n2503) );
  INV_X4 U1794 ( .A(n3450), .ZN(n3446) );
  INV_X8 U1795 ( .A(net253414), .ZN(net253424) );
  NAND2_X4 U1797 ( .A1(n3281), .A2(n2942), .ZN(n3027) );
  NAND2_X4 U1798 ( .A1(n1375), .A2(n1376), .ZN(n1378) );
  OAI22_X2 U1799 ( .A1(n2038), .A2(n2039), .B1(n2037), .B2(n1207), .ZN(n1327)
         );
  NAND2_X4 U1800 ( .A1(b[24]), .A2(n1467), .ZN(n2038) );
  NAND2_X2 U1801 ( .A1(n2768), .A2(n2769), .ZN(n2765) );
  INV_X1 U1802 ( .A(n2095), .ZN(n2096) );
  AOI21_X4 U1803 ( .B1(n3459), .B2(n3458), .A(n2006), .ZN(n3460) );
  XNOR2_X2 U1804 ( .A(n3914), .B(n3913), .ZN(net253327) );
  INV_X8 U1805 ( .A(n1461), .ZN(n1712) );
  NOR2_X2 U1806 ( .A1(net254681), .A2(net254682), .ZN(n2955) );
  OAI22_X2 U1807 ( .A1(n2032), .A2(n2033), .B1(net256018), .B2(n2031), .ZN(
        n1872) );
  NAND2_X4 U1808 ( .A1(n3756), .A2(n3755), .ZN(net253386) );
  NAND2_X2 U1809 ( .A1(n1882), .A2(net254932), .ZN(n1330) );
  NAND2_X4 U1810 ( .A1(n1328), .A2(n1329), .ZN(n1331) );
  NAND2_X4 U1811 ( .A1(n1330), .A2(n1331), .ZN(n2809) );
  INV_X4 U1812 ( .A(net254932), .ZN(n1328) );
  AND2_X4 U1813 ( .A1(net254864), .A2(net254688), .ZN(n1882) );
  NAND2_X4 U1814 ( .A1(n2809), .A2(n2788), .ZN(n2812) );
  NOR2_X2 U1815 ( .A1(net254935), .A2(net254689), .ZN(net254934) );
  INV_X32 U1816 ( .A(control[0]), .ZN(n1332) );
  INV_X32 U1817 ( .A(control[0]), .ZN(n1333) );
  XNOR2_X2 U1818 ( .A(n1806), .B(n3646), .ZN(n1901) );
  INV_X4 U1819 ( .A(n3646), .ZN(n3648) );
  INV_X4 U1820 ( .A(n1838), .ZN(n2673) );
  INV_X8 U1821 ( .A(net255428), .ZN(net257752) );
  NAND2_X4 U1822 ( .A1(n2122), .A2(n2121), .ZN(n2152) );
  INV_X4 U1823 ( .A(n3799), .ZN(n3811) );
  INV_X4 U1824 ( .A(n2506), .ZN(n2431) );
  NAND2_X4 U1825 ( .A1(n1306), .A2(n2386), .ZN(n2389) );
  NAND2_X4 U1827 ( .A1(net256795), .A2(n1691), .ZN(net254684) );
  NAND3_X2 U1828 ( .A1(b[25]), .A2(net256089), .A3(net257283), .ZN(n2102) );
  INV_X4 U1829 ( .A(net255380), .ZN(net256742) );
  NAND2_X4 U1830 ( .A1(n2622), .A2(n1789), .ZN(n2745) );
  INV_X4 U1831 ( .A(n2147), .ZN(n2115) );
  INV_X8 U1832 ( .A(net256153), .ZN(net256147) );
  INV_X2 U1833 ( .A(n1334), .ZN(n1335) );
  NAND2_X4 U1834 ( .A1(n1336), .A2(n1337), .ZN(n1339) );
  INV_X4 U1835 ( .A(n3594), .ZN(n1336) );
  INV_X2 U1836 ( .A(net257779), .ZN(n1459) );
  NOR2_X2 U1837 ( .A1(net256153), .A2(n4027), .ZN(n4032) );
  INV_X4 U1838 ( .A(net256153), .ZN(net256151) );
  INV_X1 U1839 ( .A(n2107), .ZN(n2042) );
  INV_X4 U1840 ( .A(n1123), .ZN(n1351) );
  XNOR2_X1 U1841 ( .A(n1810), .B(n3070), .ZN(n3071) );
  NAND2_X2 U1842 ( .A1(net254464), .A2(net254465), .ZN(n3248) );
  NAND2_X1 U1843 ( .A1(net255533), .A2(net255854), .ZN(net255853) );
  INV_X2 U1844 ( .A(n3033), .ZN(n1949) );
  NAND2_X2 U1845 ( .A1(net255852), .A2(net255853), .ZN(n1343) );
  NAND2_X4 U1846 ( .A1(n1341), .A2(n1342), .ZN(n1344) );
  NAND2_X4 U1847 ( .A1(n1344), .A2(n1343), .ZN(net255795) );
  INV_X4 U1848 ( .A(net255852), .ZN(n1341) );
  INV_X2 U1849 ( .A(net255853), .ZN(n1342) );
  INV_X4 U1850 ( .A(net255221), .ZN(net255441) );
  INV_X4 U1851 ( .A(net257564), .ZN(net257565) );
  INV_X4 U1852 ( .A(n1446), .ZN(net256305) );
  AOI21_X2 U1853 ( .B1(net254367), .B2(net254366), .A(net254363), .ZN(
        net254468) );
  INV_X1 U1854 ( .A(net255537), .ZN(n1345) );
  NAND2_X2 U1855 ( .A1(n3320), .A2(n3319), .ZN(n3602) );
  NAND2_X4 U1856 ( .A1(n1398), .A2(n1399), .ZN(n1706) );
  OAI21_X4 U1857 ( .B1(n3288), .B2(n1910), .A(n1777), .ZN(n3411) );
  NAND2_X1 U1858 ( .A1(n2385), .A2(n2584), .ZN(n1348) );
  NAND2_X2 U1859 ( .A1(n1346), .A2(n1347), .ZN(n1349) );
  INV_X32 U1860 ( .A(control[1]), .ZN(n1465) );
  NAND3_X2 U1861 ( .A1(n1952), .A2(n2140), .A3(n2141), .ZN(n2142) );
  INV_X8 U1862 ( .A(net255407), .ZN(net256401) );
  NAND2_X4 U1863 ( .A1(net253444), .A2(net257153), .ZN(net253443) );
  AOI22_X4 U1864 ( .A1(n3979), .A2(n1783), .B1(n3978), .B2(n3992), .ZN(n3980)
         );
  NAND2_X4 U1866 ( .A1(n1351), .A2(n1352), .ZN(n1354) );
  INV_X4 U1868 ( .A(n3072), .ZN(n1352) );
  OAI21_X4 U1869 ( .B1(n1948), .B2(net255232), .A(net255101), .ZN(net257953)
         );
  NAND2_X4 U1870 ( .A1(n2531), .A2(n2530), .ZN(n1896) );
  BUF_X32 U1871 ( .A(n3336), .Z(n1439) );
  NAND2_X4 U1872 ( .A1(n1325), .A2(n1355), .ZN(n1356) );
  NAND2_X4 U1873 ( .A1(n1356), .A2(n2034), .ZN(n2095) );
  INV_X4 U1874 ( .A(n2035), .ZN(n1355) );
  NAND2_X2 U1875 ( .A1(n2210), .A2(n2209), .ZN(n1361) );
  NAND2_X4 U1876 ( .A1(n1359), .A2(n1360), .ZN(n1362) );
  NAND2_X4 U1877 ( .A1(n1362), .A2(n1361), .ZN(n2213) );
  INV_X4 U1878 ( .A(n2210), .ZN(n1359) );
  INV_X4 U1879 ( .A(n2209), .ZN(n1360) );
  NAND2_X2 U1880 ( .A1(n1363), .A2(n1387), .ZN(n1364) );
  NAND2_X2 U1881 ( .A1(n1364), .A2(n1388), .ZN(n1976) );
  INV_X8 U1882 ( .A(n2871), .ZN(n2940) );
  INV_X4 U1883 ( .A(n2066), .ZN(n2070) );
  NAND3_X4 U1884 ( .A1(n2510), .A2(n1792), .A3(net257586), .ZN(n2592) );
  INV_X2 U1885 ( .A(n2307), .ZN(n2312) );
  NAND2_X1 U1886 ( .A1(net255546), .A2(net255583), .ZN(n1371) );
  INV_X8 U1887 ( .A(control[1]), .ZN(n1467) );
  INV_X1 U1888 ( .A(net256402), .ZN(n1391) );
  NAND2_X2 U1891 ( .A1(n1367), .A2(n1368), .ZN(n2168) );
  INV_X4 U1892 ( .A(n2166), .ZN(n1365) );
  INV_X4 U1893 ( .A(n2165), .ZN(n1366) );
  OAI21_X4 U1894 ( .B1(n2026), .B2(n2065), .A(n1940), .ZN(n1862) );
  NAND2_X4 U1895 ( .A1(n2666), .A2(n2665), .ZN(n2721) );
  INV_X2 U1896 ( .A(n3966), .ZN(n3968) );
  NAND2_X4 U1897 ( .A1(n4001), .A2(n4000), .ZN(n3998) );
  NAND2_X2 U1898 ( .A1(n1705), .A2(net253810), .ZN(n1398) );
  INV_X4 U1899 ( .A(n3116), .ZN(n3117) );
  XNOR2_X1 U1900 ( .A(net255852), .B(net255853), .ZN(net257482) );
  NAND2_X4 U1901 ( .A1(n1369), .A2(n1370), .ZN(n1372) );
  NAND2_X4 U1902 ( .A1(n1371), .A2(n1372), .ZN(net255581) );
  INV_X4 U1903 ( .A(net255583), .ZN(n1369) );
  INV_X2 U1904 ( .A(net255546), .ZN(n1370) );
  INV_X2 U1906 ( .A(n2067), .ZN(n1373) );
  INV_X8 U1907 ( .A(n2071), .ZN(n2067) );
  NAND2_X4 U1908 ( .A1(n2070), .A2(net257127), .ZN(n1802) );
  NAND2_X4 U1909 ( .A1(n2545), .A2(n2546), .ZN(n2657) );
  NAND4_X4 U1910 ( .A1(b[9]), .A2(control[1]), .A3(a[4]), .A4(net256089), .ZN(
        net255929) );
  OAI211_X4 U1911 ( .C1(n2664), .C2(n2663), .A(n1432), .B(n1273), .ZN(n2665)
         );
  NAND2_X4 U1912 ( .A1(n3835), .A2(n3836), .ZN(n3744) );
  INV_X2 U1913 ( .A(net254363), .ZN(net257864) );
  NAND2_X2 U1914 ( .A1(net254459), .A2(net254460), .ZN(net254670) );
  NAND2_X4 U1915 ( .A1(a[2]), .A2(net257127), .ZN(n2012) );
  INV_X8 U1916 ( .A(n2164), .ZN(n2266) );
  XNOR2_X2 U1917 ( .A(n2840), .B(net254856), .ZN(n1773) );
  INV_X4 U1918 ( .A(n3120), .ZN(n3043) );
  NAND2_X4 U1919 ( .A1(n2776), .A2(n1853), .ZN(n2778) );
  OAI211_X2 U1920 ( .C1(n2767), .C2(n2772), .A(n2770), .B(n2771), .ZN(n2776)
         );
  OAI211_X2 U1921 ( .C1(n3634), .C2(n1903), .A(n3637), .B(n3443), .ZN(n3451)
         );
  NAND2_X4 U1922 ( .A1(n3263), .A2(n3262), .ZN(n3502) );
  INV_X8 U1923 ( .A(n2500), .ZN(n2749) );
  NAND2_X2 U1924 ( .A1(a[12]), .A2(net256421), .ZN(n2590) );
  INV_X2 U1925 ( .A(n2940), .ZN(n2004) );
  NAND2_X4 U1926 ( .A1(n2366), .A2(net257052), .ZN(n2391) );
  NAND2_X2 U1927 ( .A1(n3271), .A2(n3173), .ZN(n3476) );
  INV_X2 U1928 ( .A(n2215), .ZN(n1518) );
  INV_X8 U1930 ( .A(net256159), .ZN(net256157) );
  NAND2_X4 U1931 ( .A1(n2769), .A2(n2771), .ZN(n2774) );
  OAI21_X2 U1932 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3865) );
  OAI21_X2 U1933 ( .B1(n3446), .B2(n3445), .A(n3448), .ZN(n1817) );
  AND3_X2 U1935 ( .A1(net255910), .A2(n2074), .A3(n2122), .ZN(n2069) );
  NAND2_X4 U1936 ( .A1(n2245), .A2(n2322), .ZN(n2258) );
  NAND2_X4 U1937 ( .A1(n2904), .A2(n3048), .ZN(n2907) );
  NAND2_X4 U1938 ( .A1(net257266), .A2(net257343), .ZN(n2918) );
  NAND2_X2 U1939 ( .A1(n1625), .A2(net254746), .ZN(net257343) );
  NAND2_X2 U1940 ( .A1(net254766), .A2(net254767), .ZN(net256680) );
  NAND2_X1 U1941 ( .A1(n2919), .A2(n2918), .ZN(n1377) );
  INV_X2 U1942 ( .A(n2919), .ZN(n1375) );
  INV_X2 U1943 ( .A(n2918), .ZN(n1376) );
  NAND2_X4 U1944 ( .A1(n1380), .A2(n1381), .ZN(net255332) );
  INV_X2 U1945 ( .A(net255501), .ZN(n1379) );
  NAND2_X2 U1946 ( .A1(net254861), .A2(net254862), .ZN(n1384) );
  NAND2_X4 U1947 ( .A1(n1382), .A2(n1383), .ZN(n1385) );
  NAND2_X4 U1948 ( .A1(n1384), .A2(n1385), .ZN(net254857) );
  INV_X4 U1949 ( .A(net254862), .ZN(n1382) );
  NAND2_X4 U1950 ( .A1(net255332), .A2(net255333), .ZN(net255329) );
  XNOR2_X2 U1951 ( .A(net255374), .B(n1386), .ZN(n1927) );
  NAND2_X2 U1953 ( .A1(n2041), .A2(n2040), .ZN(n1388) );
  NAND2_X4 U1954 ( .A1(n1387), .A2(n1363), .ZN(n1389) );
  NAND2_X4 U1955 ( .A1(n1389), .A2(n1388), .ZN(n2107) );
  BUF_X4 U1956 ( .A(a[2]), .Z(n1390) );
  INV_X4 U1957 ( .A(n3863), .ZN(n1893) );
  INV_X8 U1958 ( .A(n3866), .ZN(n3870) );
  INV_X8 U1959 ( .A(n3258), .ZN(n3917) );
  INV_X8 U1960 ( .A(net255166), .ZN(net255100) );
  NOR2_X4 U1961 ( .A1(n3755), .A2(n1876), .ZN(net253592) );
  NAND2_X4 U1962 ( .A1(n3756), .A2(n3755), .ZN(n3757) );
  NAND2_X2 U1963 ( .A1(n3414), .A2(net253820), .ZN(net253986) );
  NAND2_X1 U1964 ( .A1(n3431), .A2(n3429), .ZN(n3354) );
  NAND2_X1 U1965 ( .A1(n3429), .A2(n3430), .ZN(n3355) );
  NAND2_X4 U1966 ( .A1(n3311), .A2(n3429), .ZN(n3431) );
  OAI21_X4 U1967 ( .B1(n4074), .B2(n4073), .A(net253056), .ZN(net253043) );
  OAI211_X4 U1969 ( .C1(n3695), .C2(net256184), .A(n3694), .B(n3693), .ZN(
        n3765) );
  XNOR2_X2 U1970 ( .A(n1335), .B(n3689), .ZN(n3695) );
  NAND2_X2 U1971 ( .A1(n3688), .A2(n1895), .ZN(n3689) );
  INV_X8 U1972 ( .A(n1650), .ZN(net254942) );
  NAND2_X4 U1973 ( .A1(n3992), .A2(n3996), .ZN(n3911) );
  NAND2_X4 U1974 ( .A1(n3835), .A2(n3836), .ZN(n3837) );
  INV_X8 U1975 ( .A(n1590), .ZN(n1591) );
  AOI22_X4 U1976 ( .A1(n2750), .A2(n2751), .B1(n2749), .B2(n2748), .ZN(n2754)
         );
  NAND2_X2 U1977 ( .A1(n2463), .A2(n2462), .ZN(n1392) );
  NAND2_X4 U1978 ( .A1(n2377), .A2(n1982), .ZN(n2441) );
  INV_X4 U1981 ( .A(n3622), .ZN(n1393) );
  NAND2_X4 U1982 ( .A1(n1397), .A2(n1508), .ZN(n1399) );
  NAND2_X2 U1983 ( .A1(n3053), .A2(n3221), .ZN(n3126) );
  NOR2_X2 U1984 ( .A1(net253780), .A2(net253390), .ZN(n3612) );
  NAND2_X2 U1985 ( .A1(n1881), .A2(n1508), .ZN(n1402) );
  NAND2_X4 U1986 ( .A1(n1400), .A2(n1401), .ZN(n1403) );
  NAND2_X4 U1987 ( .A1(n1402), .A2(n1403), .ZN(net253763) );
  INV_X4 U1988 ( .A(n1508), .ZN(n1401) );
  NOR2_X4 U1989 ( .A1(net253406), .A2(net253407), .ZN(net253206) );
  INV_X4 U1990 ( .A(n1434), .ZN(net254807) );
  NOR2_X4 U1991 ( .A1(n3285), .A2(n3284), .ZN(n1777) );
  NAND4_X4 U1992 ( .A1(n1452), .A2(net254367), .A3(net254364), .A4(n1686), 
        .ZN(net254233) );
  INV_X4 U1993 ( .A(n3805), .ZN(n3802) );
  INV_X4 U1994 ( .A(n3795), .ZN(n3804) );
  NAND2_X4 U1995 ( .A1(n2833), .A2(n2708), .ZN(n2830) );
  NAND2_X2 U1997 ( .A1(n2707), .A2(n2706), .ZN(n2833) );
  NOR2_X1 U1998 ( .A1(n1701), .A2(net253111), .ZN(net253109) );
  NAND3_X2 U1999 ( .A1(n2777), .A2(a[13]), .A3(net256117), .ZN(n2892) );
  INV_X4 U2000 ( .A(n2893), .ZN(n2895) );
  INV_X4 U2001 ( .A(net255106), .ZN(net256583) );
  INV_X8 U2002 ( .A(net254463), .ZN(net254570) );
  AOI21_X2 U2003 ( .B1(n2266), .B2(n2217), .A(n2216), .ZN(n2218) );
  INV_X4 U2004 ( .A(n1877), .ZN(n1878) );
  NAND3_X2 U2005 ( .A1(n2173), .A2(n2172), .A3(n2171), .ZN(net253272) );
  NAND3_X2 U2006 ( .A1(n2244), .A2(n2243), .A3(n2242), .ZN(net253271) );
  NOR2_X2 U2007 ( .A1(n3486), .A2(n3543), .ZN(n3484) );
  OAI211_X2 U2008 ( .C1(net258044), .C2(net256184), .A(net253525), .B(n1641), 
        .ZN(net253302) );
  NOR2_X2 U2009 ( .A1(net256097), .A2(n1724), .ZN(n1723) );
  INV_X4 U2010 ( .A(n1970), .ZN(n2695) );
  INV_X4 U2011 ( .A(net257484), .ZN(net257485) );
  INV_X4 U2012 ( .A(n1857), .ZN(n2505) );
  INV_X4 U2013 ( .A(net255593), .ZN(net255592) );
  NOR2_X2 U2014 ( .A1(n3048), .A2(n3047), .ZN(n3050) );
  INV_X4 U2015 ( .A(net255044), .ZN(n1691) );
  INV_X4 U2016 ( .A(n2837), .ZN(n2838) );
  INV_X1 U2017 ( .A(n3047), .ZN(n1775) );
  INV_X2 U2018 ( .A(net254562), .ZN(net254666) );
  NAND3_X2 U2019 ( .A1(n2914), .A2(a[14]), .A3(net256135), .ZN(n3140) );
  OAI21_X1 U2020 ( .B1(n3431), .B2(n3430), .A(n3429), .ZN(n3434) );
  INV_X4 U2021 ( .A(net254570), .ZN(n1596) );
  INV_X4 U2022 ( .A(n2945), .ZN(n2667) );
  INV_X16 U2023 ( .A(net256139), .ZN(net256137) );
  INV_X4 U2024 ( .A(n3292), .ZN(n3441) );
  INV_X4 U2025 ( .A(n1648), .ZN(net256127) );
  NOR2_X2 U2026 ( .A1(net256179), .A2(n4037), .ZN(n4040) );
  NOR2_X2 U2027 ( .A1(net256111), .A2(n4038), .ZN(n4039) );
  INV_X16 U2028 ( .A(n1698), .ZN(n1701) );
  NAND2_X2 U2029 ( .A1(n2091), .A2(n2186), .ZN(n2082) );
  OAI221_X2 U2030 ( .B1(net254058), .B2(net253764), .C1(n1546), .C2(n1122), 
        .A(n3472), .ZN(n3387) );
  NAND2_X2 U2031 ( .A1(net253396), .A2(net253398), .ZN(n1743) );
  INV_X16 U2032 ( .A(net256179), .ZN(net256173) );
  NOR2_X1 U2033 ( .A1(n2995), .A2(net256184), .ZN(n2996) );
  NOR2_X1 U2034 ( .A1(n3512), .A2(n3762), .ZN(n3087) );
  INV_X4 U2035 ( .A(net253279), .ZN(net253278) );
  NOR2_X2 U2036 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  NAND2_X2 U2037 ( .A1(n2306), .A2(n2169), .ZN(n2170) );
  INV_X4 U2038 ( .A(net253053), .ZN(net256103) );
  INV_X4 U2039 ( .A(net253204), .ZN(net253274) );
  NOR2_X2 U2040 ( .A1(n1639), .A2(net253173), .ZN(n1638) );
  NOR2_X1 U2041 ( .A1(n2488), .A2(n2487), .ZN(n2489) );
  OAI21_X2 U2042 ( .B1(n2934), .B2(n3098), .A(n3094), .ZN(n2935) );
  NOR2_X1 U2043 ( .A1(net253044), .A2(n1656), .ZN(n1655) );
  AND2_X4 U2044 ( .A1(a[17]), .A2(net256125), .ZN(n1404) );
  AND2_X2 U2045 ( .A1(a[14]), .A2(net253103), .ZN(n1405) );
  NAND2_X1 U2046 ( .A1(a[8]), .A2(net256165), .ZN(n2794) );
  INV_X1 U2047 ( .A(net256101), .ZN(net256097) );
  INV_X8 U2048 ( .A(net256097), .ZN(net256095) );
  AND2_X4 U2049 ( .A1(a[13]), .A2(net256125), .ZN(n1406) );
  NAND3_X2 U2050 ( .A1(n2085), .A2(n2084), .A3(n2083), .ZN(net253231) );
  INV_X8 U2051 ( .A(net253231), .ZN(n1648) );
  AND2_X4 U2052 ( .A1(n1425), .A2(n2822), .ZN(n1407) );
  AND2_X4 U2053 ( .A1(product_in[13]), .A2(net256095), .ZN(n1408) );
  AND2_X2 U2054 ( .A1(a[6]), .A2(net256175), .ZN(n1409) );
  AND2_X4 U2055 ( .A1(a[18]), .A2(net256105), .ZN(n1410) );
  NAND2_X1 U2056 ( .A1(a[9]), .A2(net256165), .ZN(n2866) );
  INV_X16 U2057 ( .A(net256115), .ZN(net256105) );
  INV_X4 U2058 ( .A(n2278), .ZN(n1519) );
  AND3_X4 U2059 ( .A1(net256420), .A2(net257586), .A3(net255872), .ZN(n1411)
         );
  AND2_X4 U2060 ( .A1(n1390), .A2(net256137), .ZN(n1412) );
  AND2_X4 U2061 ( .A1(a[3]), .A2(a[4]), .ZN(n1413) );
  AND2_X2 U2062 ( .A1(a[7]), .A2(net256119), .ZN(n1414) );
  NAND2_X2 U2063 ( .A1(net255629), .A2(n2322), .ZN(net255627) );
  INV_X4 U2064 ( .A(net255627), .ZN(net257456) );
  XOR2_X2 U2065 ( .A(n4003), .B(n4073), .Z(n1415) );
  AND2_X4 U2066 ( .A1(a[11]), .A2(net256175), .ZN(n1416) );
  INV_X2 U2067 ( .A(net256183), .ZN(net256184) );
  INV_X4 U2068 ( .A(net253064), .ZN(net256183) );
  AND2_X4 U2069 ( .A1(a[20]), .A2(net256165), .ZN(n1417) );
  AND2_X4 U2070 ( .A1(product_in[18]), .A2(net256095), .ZN(n1418) );
  AND2_X2 U2071 ( .A1(net254467), .A2(net254464), .ZN(n1419) );
  AND2_X4 U2072 ( .A1(n2674), .A2(n2675), .ZN(n1420) );
  AND2_X4 U2073 ( .A1(net253647), .A2(net257109), .ZN(n1421) );
  AND2_X4 U2074 ( .A1(net253398), .A2(net253401), .ZN(n1422) );
  CLKBUF_X3 U2075 ( .A(n1828), .Z(n1784) );
  AND2_X4 U2076 ( .A1(a[13]), .A2(n1865), .ZN(n1423) );
  AND2_X2 U2077 ( .A1(a[0]), .A2(net256165), .ZN(n1424) );
  AND2_X4 U2078 ( .A1(a[14]), .A2(net256143), .ZN(n1425) );
  AND2_X4 U2079 ( .A1(a[16]), .A2(n1460), .ZN(n1426) );
  AND2_X4 U2080 ( .A1(a[18]), .A2(n1460), .ZN(n1427) );
  AND2_X4 U2081 ( .A1(a[22]), .A2(n1460), .ZN(n1428) );
  AND2_X4 U2082 ( .A1(a[28]), .A2(net256143), .ZN(n1429) );
  NAND2_X1 U2083 ( .A1(a[18]), .A2(net256165), .ZN(n3628) );
  INV_X4 U2084 ( .A(net255587), .ZN(net256747) );
  NAND2_X1 U2085 ( .A1(a[16]), .A2(net256165), .ZN(n3395) );
  INV_X4 U2086 ( .A(n3447), .ZN(n3444) );
  NAND2_X2 U2087 ( .A1(product_in[22]), .A2(net256095), .ZN(n3340) );
  INV_X1 U2088 ( .A(net253103), .ZN(net256111) );
  INV_X16 U2089 ( .A(net253272), .ZN(net256179) );
  INV_X8 U2090 ( .A(net256179), .ZN(net256175) );
  INV_X2 U2092 ( .A(n1431), .ZN(n1432) );
  NAND2_X4 U2093 ( .A1(n2651), .A2(n2650), .ZN(n2850) );
  XNOR2_X2 U2094 ( .A(n3079), .B(n3078), .ZN(n1433) );
  NAND2_X2 U2095 ( .A1(n3174), .A2(n1787), .ZN(n3078) );
  XNOR2_X2 U2096 ( .A(n3090), .B(n1885), .ZN(product_out[19]) );
  OAI21_X4 U2097 ( .B1(n3268), .B2(n1845), .A(n3337), .ZN(n3269) );
  XNOR2_X2 U2098 ( .A(n3270), .B(n3269), .ZN(product_out[21]) );
  INV_X4 U2100 ( .A(n3335), .ZN(n3338) );
  NAND2_X1 U2101 ( .A1(n2047), .A2(n2192), .ZN(n2048) );
  AOI21_X2 U2102 ( .B1(n2476), .B2(n2558), .A(n2556), .ZN(n2477) );
  NAND2_X2 U2104 ( .A1(n1741), .A2(n1740), .ZN(net254709) );
  INV_X4 U2106 ( .A(n2938), .ZN(n2939) );
  INV_X4 U2107 ( .A(n2738), .ZN(n2660) );
  NOR2_X2 U2108 ( .A1(n2324), .A2(n2323), .ZN(n2328) );
  BUF_X4 U2109 ( .A(n3113), .Z(n1505) );
  NAND2_X4 U2110 ( .A1(n1589), .A2(n1588), .ZN(n2813) );
  NAND2_X2 U2111 ( .A1(n1697), .A2(net256823), .ZN(net254933) );
  INV_X4 U2112 ( .A(net256823), .ZN(net254948) );
  NAND2_X2 U2113 ( .A1(n1800), .A2(n2787), .ZN(n1588) );
  INV_X4 U2114 ( .A(n3774), .ZN(n3768) );
  XNOR2_X2 U2115 ( .A(n3404), .B(n3505), .ZN(product_out[23]) );
  OAI21_X2 U2116 ( .B1(n4101), .B2(n4092), .A(n3493), .ZN(n3404) );
  AOI21_X2 U2117 ( .B1(n3509), .B2(net257630), .A(net253535), .ZN(n3518) );
  INV_X4 U2118 ( .A(n1244), .ZN(n3745) );
  INV_X4 U2119 ( .A(net254767), .ZN(net256678) );
  NAND2_X4 U2120 ( .A1(n2850), .A2(n1527), .ZN(n2857) );
  NAND2_X2 U2121 ( .A1(net254086), .A2(net254051), .ZN(n1562) );
  INV_X2 U2122 ( .A(n3516), .ZN(n3514) );
  NAND2_X4 U2123 ( .A1(n3517), .A2(n3516), .ZN(n3790) );
  OAI221_X4 U2124 ( .B1(n1139), .B2(net256184), .C1(n1889), .C2(n3512), .A(
        n3511), .ZN(n3516) );
  NOR2_X2 U2125 ( .A1(n1717), .A2(net253187), .ZN(n1716) );
  CLKBUF_X3 U2126 ( .A(n3198), .Z(n1437) );
  NAND2_X1 U2127 ( .A1(n1922), .A2(n4067), .ZN(n4070) );
  NAND2_X4 U2128 ( .A1(n1502), .A2(n1503), .ZN(n1828) );
  INV_X4 U2129 ( .A(net254291), .ZN(net254302) );
  NAND2_X4 U2130 ( .A1(n3263), .A2(n3262), .ZN(n1440) );
  INV_X8 U2131 ( .A(n3261), .ZN(n3263) );
  NAND2_X4 U2132 ( .A1(n1761), .A2(n2079), .ZN(n2091) );
  NAND2_X4 U2133 ( .A1(n1512), .A2(n1511), .ZN(net253685) );
  INV_X2 U2134 ( .A(n1974), .ZN(net255105) );
  INV_X8 U2135 ( .A(n2872), .ZN(n3024) );
  XNOR2_X2 U2138 ( .A(net254631), .B(n2984), .ZN(n1441) );
  NAND2_X4 U2139 ( .A1(n1505), .A2(n3455), .ZN(n3070) );
  NAND2_X2 U2140 ( .A1(net255165), .A2(net255164), .ZN(n1601) );
  NAND2_X4 U2141 ( .A1(n3159), .A2(n3158), .ZN(n3278) );
  XNOR2_X1 U2142 ( .A(n3853), .B(n1783), .ZN(n1442) );
  INV_X2 U2143 ( .A(n1787), .ZN(n3162) );
  NAND2_X4 U2145 ( .A1(n1597), .A2(net254751), .ZN(net254748) );
  NAND2_X2 U2146 ( .A1(n1848), .A2(n3175), .ZN(n3178) );
  INV_X4 U2147 ( .A(n2446), .ZN(n2256) );
  NAND2_X2 U2148 ( .A1(n1751), .A2(n1752), .ZN(net254140) );
  INV_X4 U2149 ( .A(n1856), .ZN(n1444) );
  INV_X4 U2150 ( .A(n2186), .ZN(n1856) );
  INV_X1 U2151 ( .A(n3003), .ZN(n1445) );
  CLKBUF_X3 U2153 ( .A(n3185), .Z(n1776) );
  INV_X2 U2154 ( .A(n2967), .ZN(n2910) );
  NAND2_X2 U2155 ( .A1(n2711), .A2(n1823), .ZN(n1446) );
  NAND2_X4 U2156 ( .A1(n3534), .A2(n3535), .ZN(n3537) );
  NAND2_X2 U2157 ( .A1(n2843), .A2(n2844), .ZN(n1848) );
  INV_X2 U2158 ( .A(n2314), .ZN(n2272) );
  NAND2_X4 U2159 ( .A1(n3470), .A2(n3469), .ZN(n3623) );
  INV_X8 U2160 ( .A(net254708), .ZN(net254367) );
  NAND2_X2 U2162 ( .A1(n3923), .A2(net253296), .ZN(n1515) );
  NAND2_X4 U2163 ( .A1(n1452), .A2(net254367), .ZN(net254631) );
  INV_X2 U2164 ( .A(n3350), .ZN(n1463) );
  NAND2_X4 U2165 ( .A1(n3685), .A2(n3686), .ZN(n1876) );
  NAND2_X4 U2166 ( .A1(n3685), .A2(n3686), .ZN(net253391) );
  OAI21_X4 U2167 ( .B1(net254695), .B2(net254709), .A(n1624), .ZN(net254708)
         );
  INV_X4 U2168 ( .A(n2758), .ZN(n1836) );
  OAI21_X4 U2169 ( .B1(n1942), .B2(net254363), .A(net254364), .ZN(net254234)
         );
  INV_X1 U2170 ( .A(net256135), .ZN(n1448) );
  NAND2_X2 U2171 ( .A1(n2837), .A2(n1450), .ZN(n1449) );
  INV_X2 U2172 ( .A(n1449), .ZN(n1447) );
  NOR2_X1 U2173 ( .A1(n2839), .A2(n1448), .ZN(n1450) );
  NAND2_X2 U2174 ( .A1(net254760), .A2(n1739), .ZN(n1736) );
  NAND2_X4 U2175 ( .A1(a[11]), .A2(net256125), .ZN(net254760) );
  NOR2_X4 U2176 ( .A1(n1974), .A2(net256583), .ZN(net256582) );
  OAI21_X4 U2177 ( .B1(n3347), .B2(net257239), .A(n1544), .ZN(n3351) );
  NOR2_X4 U2178 ( .A1(n3250), .A2(n1404), .ZN(net257239) );
  NOR2_X4 U2179 ( .A1(net253457), .A2(n1421), .ZN(n1451) );
  NAND2_X2 U2180 ( .A1(n1108), .A2(net253646), .ZN(net253457) );
  NAND2_X4 U2181 ( .A1(a[11]), .A2(net256135), .ZN(n2710) );
  OAI21_X4 U2182 ( .B1(n2953), .B2(n1453), .A(net254693), .ZN(n1452) );
  OAI21_X2 U2183 ( .B1(n2953), .B2(n1453), .A(net254693), .ZN(net254366) );
  INV_X4 U2184 ( .A(n3107), .ZN(n2990) );
  NAND2_X4 U2185 ( .A1(a[6]), .A2(net256125), .ZN(net255333) );
  NAND2_X2 U2186 ( .A1(n1430), .A2(n1457), .ZN(net255542) );
  NAND2_X2 U2187 ( .A1(n1457), .A2(net255427), .ZN(net255590) );
  NAND2_X2 U2188 ( .A1(n3185), .A2(n3281), .ZN(n2987) );
  INV_X2 U2189 ( .A(n1676), .ZN(n1677) );
  NOR3_X4 U2190 ( .A1(net253643), .A2(n1671), .A3(n1676), .ZN(n1673) );
  NAND2_X1 U2191 ( .A1(n2266), .A2(n2264), .ZN(n2269) );
  AND2_X4 U2192 ( .A1(net254235), .A2(net254238), .ZN(n1454) );
  INV_X4 U2193 ( .A(n1454), .ZN(net254411) );
  OAI21_X1 U2194 ( .B1(n3922), .B2(n3921), .A(n3920), .ZN(n1456) );
  NAND2_X4 U2195 ( .A1(net255090), .A2(n1649), .ZN(net255436) );
  NAND2_X4 U2196 ( .A1(n1501), .A2(n3333), .ZN(n1503) );
  INV_X2 U2197 ( .A(n3207), .ZN(n3123) );
  NAND2_X2 U2198 ( .A1(net255167), .A2(net255166), .ZN(n1718) );
  NOR2_X4 U2199 ( .A1(net253805), .A2(net253804), .ZN(n1703) );
  NAND3_X2 U2200 ( .A1(net253553), .A2(net253187), .A3(n3774), .ZN(n3775) );
  NAND2_X1 U2201 ( .A1(n3508), .A2(n3507), .ZN(net253187) );
  INV_X4 U2202 ( .A(net254058), .ZN(n1545) );
  OAI21_X2 U2203 ( .B1(n1456), .B2(net253296), .A(n1515), .ZN(product_out[29])
         );
  NAND2_X2 U2204 ( .A1(net255618), .A2(net255619), .ZN(n1457) );
  NAND2_X4 U2205 ( .A1(net255624), .A2(n1713), .ZN(net255618) );
  AOI21_X2 U2206 ( .B1(n1786), .B2(n1446), .A(net255044), .ZN(n1696) );
  NAND2_X4 U2207 ( .A1(a[10]), .A2(net256125), .ZN(net255044) );
  NAND3_X2 U2208 ( .A1(net253246), .A2(net256420), .A3(n1413), .ZN(n1458) );
  NAND3_X1 U2209 ( .A1(net255613), .A2(net256420), .A3(n1413), .ZN(net257778)
         );
  NAND2_X1 U2210 ( .A1(n3519), .A2(n3523), .ZN(n3084) );
  XNOR2_X2 U2211 ( .A(n1709), .B(net253580), .ZN(n1461) );
  INV_X1 U2212 ( .A(net253764), .ZN(n1462) );
  INV_X8 U2213 ( .A(n3110), .ZN(n1860) );
  AOI21_X4 U2214 ( .B1(n2916), .B2(n2917), .A(n1592), .ZN(net254767) );
  INV_X1 U2215 ( .A(n2961), .ZN(n1592) );
  NOR2_X4 U2216 ( .A1(n1993), .A2(n1788), .ZN(n3933) );
  XNOR2_X2 U2217 ( .A(n2335), .B(net255458), .ZN(n2338) );
  NAND2_X4 U2218 ( .A1(net254094), .A2(net254085), .ZN(net257109) );
  INV_X8 U2219 ( .A(net253804), .ZN(net254094) );
  AOI21_X4 U2221 ( .B1(net257456), .B2(net255322), .A(net255443), .ZN(
        net255583) );
  NAND3_X4 U2222 ( .A1(net257677), .A2(net257721), .A3(b[24]), .ZN(n1685) );
  NAND4_X4 U2223 ( .A1(n1466), .A2(b[17]), .A3(control[0]), .A4(a[4]), .ZN(
        n2101) );
  NAND3_X2 U2224 ( .A1(n2699), .A2(n2698), .A3(n2700), .ZN(n2768) );
  XNOR2_X2 U2225 ( .A(n3900), .B(n3800), .ZN(n3805) );
  NAND3_X1 U2226 ( .A1(n1976), .A2(n2027), .A3(n1862), .ZN(n2044) );
  NAND3_X4 U2227 ( .A1(net257678), .A2(net257721), .A3(b[25]), .ZN(net256063)
         );
  INV_X8 U2228 ( .A(n1898), .ZN(n2948) );
  OAI21_X2 U2229 ( .B1(n1447), .B2(net254666), .A(n1834), .ZN(n2962) );
  NOR2_X2 U2230 ( .A1(n1447), .A2(net254666), .ZN(n2917) );
  NAND2_X4 U2231 ( .A1(n3852), .A2(net253398), .ZN(n3995) );
  INV_X8 U2232 ( .A(net253651), .ZN(net257031) );
  NOR2_X2 U2233 ( .A1(net254085), .A2(net254086), .ZN(net254082) );
  INV_X8 U2234 ( .A(n3109), .ZN(n3111) );
  NAND2_X4 U2235 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND2_X4 U2236 ( .A1(n1540), .A2(n1541), .ZN(n1543) );
  NAND2_X4 U2237 ( .A1(n3138), .A2(n3193), .ZN(n3148) );
  NAND2_X1 U2238 ( .A1(n1280), .A2(n3163), .ZN(n1469) );
  NAND2_X2 U2239 ( .A1(n1468), .A2(n1132), .ZN(n1470) );
  NAND2_X2 U2240 ( .A1(n1469), .A2(n1470), .ZN(n1759) );
  OAI211_X4 U2241 ( .C1(n1859), .C2(n1909), .A(net253588), .B(n3757), .ZN(
        n3795) );
  INV_X4 U2244 ( .A(net253386), .ZN(n1676) );
  NAND2_X2 U2245 ( .A1(n1594), .A2(n3680), .ZN(n3712) );
  INV_X8 U2246 ( .A(n3767), .ZN(n3776) );
  NAND2_X4 U2247 ( .A1(n1509), .A2(n1510), .ZN(n1512) );
  NAND2_X2 U2249 ( .A1(n3851), .A2(net253407), .ZN(n1474) );
  NAND2_X4 U2250 ( .A1(n1472), .A2(n1473), .ZN(n1475) );
  NAND2_X4 U2251 ( .A1(n1474), .A2(n1475), .ZN(n3853) );
  INV_X8 U2252 ( .A(net253407), .ZN(n1473) );
  NAND2_X1 U2253 ( .A1(a[21]), .A2(net256165), .ZN(net253407) );
  NAND2_X2 U2255 ( .A1(net254696), .A2(n1434), .ZN(net254856) );
  NAND2_X4 U2256 ( .A1(n1476), .A2(n1454), .ZN(n1478) );
  NAND2_X4 U2257 ( .A1(n1477), .A2(n1478), .ZN(n3157) );
  INV_X4 U2258 ( .A(n3154), .ZN(n1476) );
  NAND2_X1 U2259 ( .A1(n3031), .A2(n2786), .ZN(n1481) );
  NAND2_X2 U2260 ( .A1(n1480), .A2(n1479), .ZN(n1482) );
  NAND2_X4 U2261 ( .A1(n1481), .A2(n1482), .ZN(net254682) );
  INV_X2 U2262 ( .A(n2786), .ZN(n1480) );
  NAND2_X1 U2263 ( .A1(net256376), .A2(net255047), .ZN(n1486) );
  INV_X2 U2264 ( .A(net256376), .ZN(n1484) );
  NAND2_X4 U2265 ( .A1(n1690), .A2(n1689), .ZN(n1686) );
  AOI21_X4 U2266 ( .B1(n2540), .B2(n2539), .A(n2538), .ZN(n2541) );
  NAND2_X4 U2267 ( .A1(n3176), .A2(n3175), .ZN(n2872) );
  AND2_X4 U2268 ( .A1(n3124), .A2(n3210), .ZN(n1961) );
  NAND2_X4 U2269 ( .A1(n3137), .A2(n1960), .ZN(n3203) );
  INV_X4 U2270 ( .A(n1646), .ZN(net257052) );
  NAND2_X4 U2271 ( .A1(n1645), .A2(net255331), .ZN(n1506) );
  INV_X4 U2272 ( .A(net255335), .ZN(n1646) );
  INV_X8 U2273 ( .A(net253390), .ZN(net253588) );
  INV_X8 U2274 ( .A(net254145), .ZN(net254237) );
  NOR2_X1 U2275 ( .A1(n2516), .A2(n2588), .ZN(n2518) );
  INV_X2 U2276 ( .A(n2697), .ZN(n2587) );
  NAND2_X4 U2277 ( .A1(net254577), .A2(net254470), .ZN(n2984) );
  INV_X8 U2278 ( .A(n1630), .ZN(net253805) );
  NAND2_X4 U2279 ( .A1(n3184), .A2(n3185), .ZN(n1910) );
  NAND2_X2 U2280 ( .A1(n2155), .A2(n2154), .ZN(n1490) );
  NAND2_X2 U2281 ( .A1(n1998), .A2(n1489), .ZN(n1491) );
  NAND2_X2 U2282 ( .A1(n1490), .A2(n1491), .ZN(n2156) );
  INV_X2 U2283 ( .A(n2154), .ZN(n1489) );
  NAND3_X4 U2284 ( .A1(n2639), .A2(a[6]), .A3(net256165), .ZN(n2734) );
  NAND2_X4 U2285 ( .A1(n1539), .A2(n1538), .ZN(n3622) );
  NAND2_X4 U2286 ( .A1(n1536), .A2(n1537), .ZN(n1539) );
  NAND2_X4 U2287 ( .A1(n1834), .A2(net254669), .ZN(n3034) );
  OAI21_X4 U2288 ( .B1(n1911), .B2(n3107), .A(n3106), .ZN(n3520) );
  INV_X8 U2290 ( .A(net254470), .ZN(net254363) );
  NAND2_X4 U2291 ( .A1(n1612), .A2(n1613), .ZN(n1492) );
  NAND2_X2 U2292 ( .A1(n3452), .A2(n3608), .ZN(n1495) );
  NAND2_X4 U2293 ( .A1(n1493), .A2(n1494), .ZN(n1496) );
  NAND2_X4 U2294 ( .A1(n1495), .A2(n1496), .ZN(n3465) );
  INV_X4 U2295 ( .A(n3452), .ZN(n1493) );
  INV_X4 U2296 ( .A(n3608), .ZN(n1494) );
  NAND2_X2 U2297 ( .A1(n1612), .A2(n1613), .ZN(net253819) );
  OAI21_X4 U2298 ( .B1(net255547), .B2(net255548), .A(net255440), .ZN(
        net255546) );
  NAND2_X4 U2299 ( .A1(n3537), .A2(n3536), .ZN(n3541) );
  NAND2_X4 U2300 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  NOR2_X2 U2301 ( .A1(n1422), .A2(n1745), .ZN(net253320) );
  NOR2_X2 U2302 ( .A1(n3758), .A2(net253522), .ZN(n1603) );
  INV_X8 U2303 ( .A(net253391), .ZN(net253522) );
  NOR2_X4 U2304 ( .A1(net255456), .A2(net255457), .ZN(net255445) );
  NAND2_X2 U2305 ( .A1(n1566), .A2(n1567), .ZN(net255440) );
  NAND2_X4 U2306 ( .A1(net253460), .A2(n3850), .ZN(n3993) );
  INV_X4 U2307 ( .A(net253411), .ZN(net253425) );
  NOR2_X4 U2308 ( .A1(n2668), .A2(n2667), .ZN(n2670) );
  NAND2_X4 U2309 ( .A1(n3864), .A2(n3863), .ZN(n3934) );
  NAND2_X4 U2310 ( .A1(n3632), .A2(n1537), .ZN(n3701) );
  INV_X4 U2311 ( .A(net255874), .ZN(net255916) );
  XNOR2_X2 U2312 ( .A(n3073), .B(n3072), .ZN(n3075) );
  AOI21_X2 U2313 ( .B1(n3769), .B2(net253553), .A(n3768), .ZN(n3773) );
  INV_X8 U2314 ( .A(net254296), .ZN(net254293) );
  OAI211_X4 U2315 ( .C1(net256153), .C2(n1373), .A(n2105), .B(n1862), .ZN(
        n2073) );
  NAND2_X4 U2316 ( .A1(n2074), .A2(n2073), .ZN(n2075) );
  NAND2_X4 U2317 ( .A1(n1571), .A2(n1570), .ZN(n2845) );
  NAND2_X1 U2318 ( .A1(n3181), .A2(n2792), .ZN(n1499) );
  INV_X2 U2319 ( .A(n2792), .ZN(n1498) );
  NAND2_X4 U2320 ( .A1(net255506), .A2(net255507), .ZN(net256296) );
  NAND2_X4 U2321 ( .A1(n2201), .A2(n2252), .ZN(n2253) );
  INV_X8 U2322 ( .A(n1851), .ZN(n1852) );
  AOI211_X4 U2323 ( .C1(net253385), .C2(n1677), .A(n1671), .B(net253388), .ZN(
        net253380) );
  OAI21_X2 U2324 ( .B1(net257838), .B2(n1705), .A(net253391), .ZN(net253385)
         );
  INV_X2 U2325 ( .A(net255543), .ZN(net255616) );
  INV_X2 U2326 ( .A(net253274), .ZN(net257023) );
  NAND2_X4 U2327 ( .A1(n1620), .A2(n1621), .ZN(n1623) );
  AOI21_X2 U2328 ( .B1(net253205), .B2(net257023), .A(n1788), .ZN(n3990) );
  INV_X1 U2329 ( .A(n2875), .ZN(n1504) );
  NAND3_X2 U2330 ( .A1(net254234), .A2(net254233), .A3(net254235), .ZN(
        net254361) );
  INV_X4 U2331 ( .A(n3253), .ZN(n1507) );
  XNOR2_X2 U2332 ( .A(n3344), .B(n3388), .ZN(n1779) );
  INV_X2 U2333 ( .A(net253553), .ZN(net253557) );
  NAND2_X4 U2334 ( .A1(n1687), .A2(n1688), .ZN(net254238) );
  INV_X8 U2335 ( .A(n2185), .ZN(n2189) );
  NAND2_X2 U2336 ( .A1(n1976), .A2(n1802), .ZN(n2074) );
  NOR2_X4 U2337 ( .A1(net257469), .A2(net255868), .ZN(net257693) );
  NOR2_X2 U2338 ( .A1(net254689), .A2(net254690), .ZN(net254687) );
  INV_X32 U2339 ( .A(a[4]), .ZN(net255488) );
  NAND2_X4 U2340 ( .A1(n3217), .A2(n3218), .ZN(n3304) );
  NAND2_X4 U2341 ( .A1(n3362), .A2(n3363), .ZN(n3416) );
  NAND2_X2 U2342 ( .A1(n3676), .A2(n3675), .ZN(n3809) );
  AOI21_X2 U2343 ( .B1(n1870), .B2(n3799), .A(n3801), .ZN(n3752) );
  NAND4_X4 U2344 ( .A1(b[8]), .A2(n1332), .A3(a[1]), .A4(control[1]), .ZN(
        n2022) );
  NAND2_X4 U2345 ( .A1(b[9]), .A2(control[1]), .ZN(n2029) );
  NAND2_X4 U2346 ( .A1(b[8]), .A2(control[1]), .ZN(n2035) );
  INV_X8 U2347 ( .A(net253588), .ZN(n1705) );
  NAND2_X2 U2348 ( .A1(net253690), .A2(net253691), .ZN(n1511) );
  INV_X4 U2349 ( .A(net253691), .ZN(n1510) );
  INV_X4 U2350 ( .A(net253448), .ZN(net253446) );
  NAND2_X4 U2351 ( .A1(n1513), .A2(n3006), .ZN(n1514) );
  NAND2_X4 U2352 ( .A1(n1514), .A2(n3336), .ZN(n3500) );
  NAND2_X4 U2353 ( .A1(n3336), .A2(n3337), .ZN(n3497) );
  NAND3_X2 U2354 ( .A1(net256402), .A2(n1840), .A3(net256527), .ZN(n2369) );
  NAND2_X4 U2355 ( .A1(n3051), .A2(n3217), .ZN(n3053) );
  INV_X4 U2356 ( .A(n2826), .ZN(n2827) );
  INV_X4 U2357 ( .A(n1779), .ZN(n3254) );
  OR2_X4 U2358 ( .A1(net256179), .A2(net254628), .ZN(n1516) );
  NAND2_X4 U2359 ( .A1(n2986), .A2(n1516), .ZN(n3281) );
  INV_X32 U2360 ( .A(a[12]), .ZN(net254628) );
  XNOR2_X2 U2361 ( .A(net254631), .B(n2984), .ZN(n2985) );
  NAND2_X2 U2362 ( .A1(net256135), .A2(a[13]), .ZN(n1517) );
  NAND2_X4 U2363 ( .A1(n2838), .A2(n1517), .ZN(n2961) );
  INV_X16 U2364 ( .A(net253237), .ZN(net256139) );
  INV_X32 U2365 ( .A(a[13]), .ZN(n2839) );
  NAND2_X2 U2366 ( .A1(n1518), .A2(n1519), .ZN(n1521) );
  NAND2_X4 U2367 ( .A1(n1520), .A2(n1521), .ZN(n2219) );
  NAND2_X1 U2368 ( .A1(n2219), .A2(n1824), .ZN(n1524) );
  NAND2_X4 U2369 ( .A1(n1522), .A2(n1523), .ZN(n1525) );
  NAND2_X2 U2370 ( .A1(n1524), .A2(n1525), .ZN(n1951) );
  INV_X4 U2371 ( .A(n2219), .ZN(n1522) );
  INV_X2 U2372 ( .A(n1824), .ZN(n1523) );
  NAND2_X1 U2373 ( .A1(n2851), .A2(n2852), .ZN(n1526) );
  INV_X4 U2374 ( .A(n1526), .ZN(n1527) );
  NAND2_X4 U2375 ( .A1(n1390), .A2(net253103), .ZN(n2278) );
  NAND2_X4 U2376 ( .A1(n2728), .A2(n2727), .ZN(n2852) );
  NAND2_X4 U2377 ( .A1(n2938), .A2(n2004), .ZN(n3181) );
  INV_X4 U2378 ( .A(net254675), .ZN(net254939) );
  NAND2_X1 U2379 ( .A1(n3702), .A2(n3623), .ZN(n3543) );
  OAI21_X4 U2380 ( .B1(net255437), .B2(net255438), .A(n1249), .ZN(net255090)
         );
  OAI21_X4 U2381 ( .B1(n2870), .B2(n1994), .A(n1455), .ZN(n2936) );
  NAND2_X2 U2382 ( .A1(n3007), .A2(n3008), .ZN(n2735) );
  OAI21_X2 U2383 ( .B1(n3044), .B2(n3207), .A(n3116), .ZN(n3061) );
  NAND2_X2 U2384 ( .A1(n2865), .A2(n2849), .ZN(n1529) );
  NAND2_X4 U2385 ( .A1(n1528), .A2(n2863), .ZN(n1530) );
  NAND2_X4 U2386 ( .A1(n1529), .A2(n1530), .ZN(n1839) );
  INV_X4 U2387 ( .A(n2849), .ZN(n1528) );
  NAND2_X2 U2388 ( .A1(n2472), .A2(n2471), .ZN(n1533) );
  NAND2_X4 U2389 ( .A1(n1531), .A2(n1532), .ZN(n1534) );
  NAND2_X4 U2390 ( .A1(n1533), .A2(n1534), .ZN(n2494) );
  INV_X4 U2391 ( .A(n2472), .ZN(n1531) );
  INV_X4 U2392 ( .A(n2471), .ZN(n1532) );
  OAI22_X4 U2393 ( .A1(n2475), .A2(n2474), .B1(n2559), .B2(n2560), .ZN(n1535)
         );
  NAND2_X2 U2394 ( .A1(n2630), .A2(n2533), .ZN(n2471) );
  OAI22_X2 U2395 ( .A1(n2475), .A2(n2474), .B1(n2559), .B2(n2560), .ZN(n2654)
         );
  NAND2_X4 U2396 ( .A1(n1633), .A2(net254871), .ZN(net254673) );
  INV_X4 U2397 ( .A(net256375), .ZN(n1536) );
  INV_X2 U2398 ( .A(n3628), .ZN(n1537) );
  NAND2_X4 U2399 ( .A1(n1542), .A2(n1543), .ZN(n3385) );
  INV_X4 U2400 ( .A(n3383), .ZN(n1541) );
  NAND2_X2 U2401 ( .A1(n2628), .A2(n1897), .ZN(n2539) );
  NAND2_X4 U2402 ( .A1(n3845), .A2(n3844), .ZN(n3897) );
  INV_X4 U2403 ( .A(n3897), .ZN(n3941) );
  NAND2_X4 U2404 ( .A1(n1893), .A2(n3848), .ZN(n3938) );
  OAI221_X1 U2405 ( .B1(n3618), .B2(n1133), .C1(n4102), .C2(n3616), .A(
        net256099), .ZN(n3619) );
  NAND2_X2 U2406 ( .A1(n2259), .A2(n1755), .ZN(n2316) );
  NAND2_X1 U2407 ( .A1(n2285), .A2(n2284), .ZN(n1549) );
  NAND2_X2 U2408 ( .A1(n1547), .A2(n1548), .ZN(n1550) );
  NAND2_X2 U2409 ( .A1(n1549), .A2(n1550), .ZN(n1831) );
  INV_X1 U2410 ( .A(n2285), .ZN(n1547) );
  INV_X2 U2411 ( .A(n2284), .ZN(n1548) );
  NAND2_X2 U2412 ( .A1(n1840), .A2(net256402), .ZN(n2204) );
  NOR2_X4 U2413 ( .A1(n1497), .A2(n3160), .ZN(n3164) );
  NAND2_X4 U2414 ( .A1(n2239), .A2(n2238), .ZN(n2291) );
  INV_X2 U2415 ( .A(n2659), .ZN(n2661) );
  NAND2_X2 U2416 ( .A1(n1551), .A2(n1552), .ZN(n1553) );
  INV_X1 U2417 ( .A(n2110), .ZN(n1552) );
  INV_X4 U2418 ( .A(n3677), .ZN(n1937) );
  NAND2_X2 U2419 ( .A1(n3995), .A2(n1930), .ZN(n1556) );
  NAND2_X4 U2420 ( .A1(n1554), .A2(n1555), .ZN(n1557) );
  NAND2_X4 U2421 ( .A1(n1556), .A2(n1557), .ZN(net253406) );
  INV_X4 U2422 ( .A(n1930), .ZN(n1555) );
  NAND2_X4 U2423 ( .A1(n1559), .A2(net253443), .ZN(n3852) );
  NAND2_X4 U2424 ( .A1(n1563), .A2(n1562), .ZN(net253804) );
  INV_X4 U2425 ( .A(net254086), .ZN(n1560) );
  INV_X1 U2426 ( .A(net254051), .ZN(n1561) );
  NOR2_X4 U2427 ( .A1(net253406), .A2(net253407), .ZN(n1788) );
  NAND2_X4 U2428 ( .A1(n2139), .A2(n2152), .ZN(n2195) );
  INV_X4 U2429 ( .A(net253650), .ZN(net253445) );
  INV_X4 U2430 ( .A(n3053), .ZN(n3055) );
  NAND2_X4 U2431 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  NAND2_X1 U2432 ( .A1(net255585), .A2(net255584), .ZN(n1566) );
  NAND2_X4 U2433 ( .A1(n1564), .A2(n1565), .ZN(n1567) );
  INV_X4 U2434 ( .A(net255584), .ZN(n1564) );
  INV_X2 U2435 ( .A(net255585), .ZN(n1565) );
  INV_X2 U2436 ( .A(net253547), .ZN(net253289) );
  NAND2_X4 U2437 ( .A1(n1569), .A2(n2869), .ZN(n1571) );
  INV_X4 U2438 ( .A(n2807), .ZN(n1569) );
  NAND2_X1 U2439 ( .A1(n2082), .A2(n2183), .ZN(n1574) );
  NAND2_X2 U2440 ( .A1(n1572), .A2(n1573), .ZN(n1575) );
  NAND2_X2 U2441 ( .A1(n1574), .A2(n1575), .ZN(n2087) );
  INV_X1 U2442 ( .A(n2183), .ZN(n1573) );
  INV_X4 U2443 ( .A(n2087), .ZN(n2088) );
  NAND2_X1 U2444 ( .A1(n1153), .A2(n2640), .ZN(n1578) );
  NAND2_X4 U2445 ( .A1(n1576), .A2(n1577), .ZN(n1579) );
  NAND2_X2 U2446 ( .A1(n1578), .A2(n1579), .ZN(n1944) );
  INV_X4 U2448 ( .A(n2640), .ZN(n1577) );
  INV_X1 U2449 ( .A(n3020), .ZN(n2937) );
  NAND2_X4 U2450 ( .A1(n1639), .A2(net256095), .ZN(net253176) );
  INV_X4 U2452 ( .A(n3171), .ZN(n1580) );
  OAI21_X2 U2453 ( .B1(n3761), .B2(net256095), .A(n3088), .ZN(n1939) );
  XNOR2_X2 U2454 ( .A(n2922), .B(n2921), .ZN(n2926) );
  INV_X4 U2455 ( .A(net253442), .ZN(net253449) );
  NAND2_X4 U2456 ( .A1(n1805), .A2(n2315), .ZN(n2166) );
  INV_X4 U2457 ( .A(n3524), .ZN(n1583) );
  NOR2_X4 U2459 ( .A1(n1586), .A2(net254807), .ZN(n2882) );
  NAND2_X4 U2460 ( .A1(n1507), .A2(n3255), .ZN(n1593) );
  INV_X4 U2461 ( .A(n2195), .ZN(n2143) );
  INV_X4 U2462 ( .A(n1800), .ZN(n1587) );
  NAND3_X4 U2463 ( .A1(control[0]), .A2(control[1]), .A3(a[2]), .ZN(n1590) );
  NAND2_X4 U2464 ( .A1(n1591), .A2(b[1]), .ZN(n2028) );
  INV_X4 U2465 ( .A(n2961), .ZN(n3032) );
  OAI21_X4 U2466 ( .B1(n3811), .B2(n3810), .A(n3899), .ZN(n3847) );
  NAND2_X4 U2467 ( .A1(n2197), .A2(net257778), .ZN(net255915) );
  INV_X4 U2468 ( .A(n2491), .ZN(n1932) );
  NAND2_X2 U2469 ( .A1(net253038), .A2(net253039), .ZN(n1622) );
  NAND2_X4 U2470 ( .A1(n3254), .A2(n3255), .ZN(n1769) );
  CLKBUF_X3 U2471 ( .A(n3344), .Z(n1774) );
  CLKBUF_X3 U2472 ( .A(n3536), .Z(n1992) );
  NAND2_X4 U2473 ( .A1(n1455), .A2(n3015), .ZN(n3016) );
  NOR2_X2 U2474 ( .A1(n2664), .A2(n2548), .ZN(n2549) );
  NAND2_X4 U2475 ( .A1(n2572), .A2(n2548), .ZN(n2499) );
  CLKBUF_X3 U2476 ( .A(n3708), .Z(n1619) );
  INV_X8 U2477 ( .A(n3279), .ZN(n3412) );
  INV_X2 U2478 ( .A(n1937), .ZN(n1594) );
  INV_X4 U2479 ( .A(n2609), .ZN(n2502) );
  INV_X2 U2480 ( .A(net254571), .ZN(n1595) );
  NAND2_X4 U2481 ( .A1(n2289), .A2(n2288), .ZN(n2305) );
  OAI211_X4 U2482 ( .C1(n4111), .C2(net256095), .A(n2726), .B(n2725), .ZN(
        n2729) );
  AOI21_X4 U2483 ( .B1(n2540), .B2(n2539), .A(n2538), .ZN(n1867) );
  NOR2_X4 U2484 ( .A1(net255442), .A2(net257363), .ZN(net255545) );
  XNOR2_X2 U2485 ( .A(n2671), .B(n2747), .ZN(n2633) );
  NAND2_X2 U2486 ( .A1(n2718), .A2(n2717), .ZN(n1598) );
  INV_X2 U2487 ( .A(net255164), .ZN(n1599) );
  INV_X1 U2488 ( .A(net255165), .ZN(n1600) );
  XNOR2_X2 U2489 ( .A(net255164), .B(net255165), .ZN(n1789) );
  NAND2_X4 U2490 ( .A1(net253286), .A2(net253194), .ZN(n3928) );
  NAND2_X4 U2491 ( .A1(net253697), .A2(n1605), .ZN(net253693) );
  INV_X4 U2492 ( .A(n3685), .ZN(n1604) );
  NAND2_X2 U2493 ( .A1(net253429), .A2(n1742), .ZN(n1608) );
  NAND2_X4 U2494 ( .A1(n1606), .A2(n1607), .ZN(n1609) );
  NAND2_X4 U2495 ( .A1(n1608), .A2(n1609), .ZN(net253427) );
  INV_X4 U2496 ( .A(net253429), .ZN(n1606) );
  INV_X4 U2497 ( .A(n1742), .ZN(n1607) );
  NAND2_X2 U2498 ( .A1(n3465), .A2(n3464), .ZN(n1612) );
  NAND2_X4 U2499 ( .A1(n1610), .A2(n1611), .ZN(n1613) );
  INV_X4 U2500 ( .A(n3465), .ZN(n1610) );
  INV_X4 U2501 ( .A(n3464), .ZN(n1611) );
  NAND2_X2 U2502 ( .A1(n3463), .A2(n1878), .ZN(n3464) );
  NAND2_X4 U2504 ( .A1(n3307), .A2(n3306), .ZN(n3358) );
  NAND2_X4 U2505 ( .A1(n3754), .A2(n3753), .ZN(net253452) );
  INV_X4 U2506 ( .A(n3271), .ZN(n3272) );
  NAND2_X4 U2507 ( .A1(n2148), .A2(n1815), .ZN(n2149) );
  CLKBUF_X3 U2508 ( .A(n3208), .Z(n1614) );
  NAND2_X2 U2509 ( .A1(n3683), .A2(n3684), .ZN(n1617) );
  NAND2_X4 U2510 ( .A1(n1615), .A2(n1616), .ZN(n1618) );
  NAND2_X4 U2511 ( .A1(n1617), .A2(n1618), .ZN(n3797) );
  INV_X4 U2512 ( .A(n3683), .ZN(n1615) );
  INV_X4 U2513 ( .A(n3684), .ZN(n1616) );
  NAND2_X4 U2514 ( .A1(n3796), .A2(n3797), .ZN(net253519) );
  INV_X8 U2515 ( .A(n3797), .ZN(n3755) );
  NAND4_X4 U2516 ( .A1(a[17]), .A2(n3126), .A3(n3056), .A4(net256117), .ZN(
        n3205) );
  NAND2_X4 U2517 ( .A1(n1733), .A2(net255706), .ZN(net257240) );
  NAND2_X4 U2518 ( .A1(n2295), .A2(n2296), .ZN(n2347) );
  NAND2_X2 U2519 ( .A1(n1623), .A2(n1622), .ZN(product_out[31]) );
  INV_X4 U2520 ( .A(net253038), .ZN(n1620) );
  INV_X2 U2521 ( .A(net253039), .ZN(n1621) );
  NAND2_X4 U2522 ( .A1(n1653), .A2(n1654), .ZN(net253039) );
  NAND2_X4 U2523 ( .A1(net254746), .A2(n1625), .ZN(n1624) );
  INV_X4 U2524 ( .A(net254744), .ZN(n1625) );
  INV_X4 U2525 ( .A(net256700), .ZN(net254746) );
  XNOR2_X2 U2526 ( .A(net256974), .B(net254747), .ZN(net256700) );
  INV_X8 U2527 ( .A(net254462), .ZN(net254571) );
  NAND2_X2 U2528 ( .A1(a[12]), .A2(net256105), .ZN(net254744) );
  NAND2_X4 U2529 ( .A1(net254743), .A2(net254744), .ZN(net254711) );
  NAND2_X4 U2530 ( .A1(net257880), .A2(net254460), .ZN(net254747) );
  XNOR2_X2 U2531 ( .A(net254748), .B(net254747), .ZN(net254743) );
  INV_X8 U2532 ( .A(net257703), .ZN(net254460) );
  NAND2_X2 U2533 ( .A1(net254460), .A2(net254467), .ZN(net254566) );
  NAND3_X4 U2534 ( .A1(net254459), .A2(net254460), .A3(net254461), .ZN(
        net254296) );
  NOR2_X4 U2535 ( .A1(n1627), .A2(n1406), .ZN(net257703) );
  INV_X8 U2536 ( .A(n1626), .ZN(n1627) );
  NAND2_X4 U2537 ( .A1(n1406), .A2(n1627), .ZN(net257880) );
  NAND2_X4 U2538 ( .A1(n1406), .A2(n1627), .ZN(net254465) );
  NAND2_X4 U2539 ( .A1(net256680), .A2(n1629), .ZN(n1626) );
  NAND2_X4 U2540 ( .A1(net256678), .A2(n1628), .ZN(n1629) );
  INV_X4 U2541 ( .A(net254766), .ZN(n1628) );
  NAND2_X4 U2542 ( .A1(n1104), .A2(net254149), .ZN(n1630) );
  INV_X4 U2543 ( .A(net254181), .ZN(net254149) );
  NAND2_X4 U2544 ( .A1(net254150), .A2(net254149), .ZN(net257069) );
  NAND2_X2 U2545 ( .A1(net254149), .A2(net254150), .ZN(net257068) );
  NAND2_X2 U2546 ( .A1(a[16]), .A2(net256173), .ZN(net254181) );
  NAND2_X2 U2547 ( .A1(net254140), .A2(net254050), .ZN(net254183) );
  NAND3_X4 U2548 ( .A1(net254142), .A2(n1443), .A3(n1631), .ZN(net253820) );
  INV_X4 U2549 ( .A(net254050), .ZN(net253815) );
  OAI21_X4 U2550 ( .B1(net256947), .B2(net254143), .A(n1488), .ZN(n1631) );
  NAND3_X4 U2551 ( .A1(net254573), .A2(net256953), .A3(net254752), .ZN(
        net254751) );
  INV_X4 U2552 ( .A(net254574), .ZN(net254752) );
  NAND2_X4 U2553 ( .A1(net254753), .A2(net254941), .ZN(net254573) );
  NAND3_X2 U2554 ( .A1(net254572), .A2(net254573), .A3(net254465), .ZN(
        net254567) );
  INV_X2 U2555 ( .A(net254755), .ZN(net254753) );
  NAND2_X4 U2556 ( .A1(net254870), .A2(net254690), .ZN(net256953) );
  INV_X4 U2557 ( .A(net254871), .ZN(net254690) );
  NAND2_X4 U2558 ( .A1(net254870), .A2(net254690), .ZN(net254463) );
  XNOR2_X2 U2559 ( .A(net254872), .B(net254873), .ZN(net254680) );
  NAND2_X2 U2560 ( .A1(net257064), .A2(net254688), .ZN(net254574) );
  NOR2_X2 U2561 ( .A1(net254570), .A2(net254574), .ZN(net254572) );
  INV_X4 U2562 ( .A(net254689), .ZN(net257064) );
  AOI22_X2 U2563 ( .A1(net254933), .A2(net257064), .B1(net254934), .B2(
        net254868), .ZN(net254932) );
  NAND3_X2 U2564 ( .A1(net254755), .A2(net254688), .A3(net257064), .ZN(
        net254865) );
  INV_X8 U2565 ( .A(net254756), .ZN(net254689) );
  OAI211_X2 U2566 ( .C1(net254863), .C2(net254941), .A(net254865), .B(
        net254864), .ZN(net254862) );
  NAND2_X4 U2567 ( .A1(net254940), .A2(net254941), .ZN(net254675) );
  XNOR2_X2 U2568 ( .A(net254872), .B(net254873), .ZN(n1633) );
  XNOR2_X1 U2569 ( .A(net254872), .B(net254873), .ZN(net257979) );
  NAND2_X1 U2570 ( .A1(net254688), .A2(net254756), .ZN(net254863) );
  NAND2_X4 U2571 ( .A1(net256063), .A2(net256062), .ZN(net256061) );
  NAND2_X4 U2572 ( .A1(net255796), .A2(net255795), .ZN(net255622) );
  OAI21_X1 U2573 ( .B1(net255626), .B2(net255622), .A(n1258), .ZN(net255773)
         );
  NAND3_X2 U2574 ( .A1(net255622), .A2(n1258), .A3(net255434), .ZN(net255619)
         );
  NAND2_X4 U2575 ( .A1(net255867), .A2(net255868), .ZN(net255796) );
  NAND2_X2 U2576 ( .A1(net255796), .A2(net257482), .ZN(net255725) );
  INV_X1 U2577 ( .A(net255796), .ZN(net257589) );
  XNOR2_X2 U2578 ( .A(net255870), .B(net255871), .ZN(net255867) );
  INV_X1 U2579 ( .A(net255533), .ZN(net255871) );
  XNOR2_X2 U2580 ( .A(net255870), .B(net255871), .ZN(net257469) );
  AOI21_X1 U2581 ( .B1(net255779), .B2(net255915), .A(n1391), .ZN(net255785)
         );
  NOR2_X4 U2582 ( .A1(n1227), .A2(net256401), .ZN(net255875) );
  NAND3_X2 U2583 ( .A1(n1999), .A2(net255613), .A3(n1635), .ZN(net255407) );
  NOR2_X4 U2584 ( .A1(net255488), .A2(n1634), .ZN(n1635) );
  INV_X4 U2585 ( .A(a[5]), .ZN(n1634) );
  OAI22_X4 U2586 ( .A1(net257585), .A2(n1634), .B1(net256159), .B2(net255718), 
        .ZN(net255855) );
  NOR2_X4 U2587 ( .A1(n1634), .A2(net255718), .ZN(net255872) );
  OAI21_X4 U2588 ( .B1(net256179), .B2(net255488), .A(net255489), .ZN(
        net257702) );
  OAI21_X2 U2589 ( .B1(net256179), .B2(net255488), .A(net255489), .ZN(
        net255341) );
  NOR2_X4 U2590 ( .A1(net255488), .A2(control[1]), .ZN(net257283) );
  INV_X8 U2591 ( .A(net255613), .ZN(net257585) );
  NAND2_X4 U2592 ( .A1(net256054), .A2(net256055), .ZN(net255613) );
  OAI21_X4 U2594 ( .B1(net253164), .B2(net253165), .A(net253166), .ZN(
        net253161) );
  NOR2_X4 U2595 ( .A1(n1637), .A2(n1638), .ZN(n1636) );
  INV_X4 U2596 ( .A(net253302), .ZN(n1639) );
  NAND2_X2 U2597 ( .A1(n1639), .A2(net253274), .ZN(net253419) );
  OAI21_X2 U2598 ( .B1(n1639), .B2(net253173), .A(net253177), .ZN(net253165)
         );
  AOI21_X4 U2599 ( .B1(n1640), .B2(net253173), .A(n1140), .ZN(n1637) );
  OAI21_X4 U2600 ( .B1(net253572), .B2(net256095), .A(n1140), .ZN(net253547)
         );
  INV_X1 U2601 ( .A(net253570), .ZN(n1643) );
  INV_X4 U2602 ( .A(net253176), .ZN(n1640) );
  INV_X32 U2604 ( .A(net256103), .ZN(net256101) );
  INV_X32 U2605 ( .A(net256101), .ZN(net256099) );
  NAND2_X4 U2606 ( .A1(control[0]), .A2(control[1]), .ZN(net253053) );
  NOR2_X4 U2607 ( .A1(net253274), .A2(net253302), .ZN(net253421) );
  NAND2_X2 U2608 ( .A1(n1642), .A2(net253067), .ZN(n1641) );
  INV_X8 U2609 ( .A(net253308), .ZN(net253067) );
  INV_X4 U2610 ( .A(net254390), .ZN(n1642) );
  MUX2_X2 U2611 ( .A(product_in[4]), .B(n1642), .S(net256099), .Z(
        product_out[4]) );
  NAND2_X2 U2612 ( .A1(n1642), .A2(net256183), .ZN(net255247) );
  NAND2_X4 U2613 ( .A1(net255966), .A2(net255967), .ZN(net255914) );
  NAND2_X4 U2614 ( .A1(net255914), .A2(net255964), .ZN(net255877) );
  NAND2_X2 U2615 ( .A1(a[3]), .A2(n1232), .ZN(net255966) );
  NAND2_X2 U2616 ( .A1(net255967), .A2(net255966), .ZN(net255936) );
  NAND2_X4 U2617 ( .A1(n1865), .A2(a[4]), .ZN(net255967) );
  NAND3_X2 U2618 ( .A1(net255720), .A2(net255613), .A3(net255611), .ZN(
        net255409) );
  OAI21_X4 U2619 ( .B1(net256870), .B2(net255333), .A(n1646), .ZN(n1645) );
  INV_X4 U2620 ( .A(net255500), .ZN(net256870) );
  NAND2_X4 U2621 ( .A1(net255500), .A2(net255499), .ZN(net255327) );
  NAND2_X4 U2622 ( .A1(n1647), .A2(net255376), .ZN(net255331) );
  INV_X4 U2623 ( .A(net255378), .ZN(n1647) );
  INV_X4 U2624 ( .A(net255333), .ZN(net255499) );
  INV_X32 U2625 ( .A(n1648), .ZN(net256125) );
  NAND2_X2 U2626 ( .A1(net255582), .A2(net255581), .ZN(net255335) );
  NAND2_X2 U2627 ( .A1(net255335), .A2(net255459), .ZN(net255458) );
  INV_X8 U2628 ( .A(n1644), .ZN(n1649) );
  NAND4_X2 U2629 ( .A1(net255089), .A2(net255091), .A3(net256907), .A4(n1649), 
        .ZN(net254992) );
  NAND3_X2 U2630 ( .A1(net255320), .A2(n1649), .A3(net256907), .ZN(net255318)
         );
  INV_X8 U2631 ( .A(net255092), .ZN(n1644) );
  NOR2_X1 U2632 ( .A1(n1644), .A2(net255225), .ZN(net255223) );
  AOI22_X2 U2633 ( .A1(net255545), .A2(net255221), .B1(net255546), .B2(
        net257522), .ZN(net255501) );
  INV_X8 U2634 ( .A(net256061), .ZN(net256054) );
  NAND3_X4 U2635 ( .A1(net257782), .A2(control[0]), .A3(b[17]), .ZN(net256062)
         );
  INV_X32 U2636 ( .A(control[1]), .ZN(net257782) );
  NAND2_X4 U2637 ( .A1(net255324), .A2(net255107), .ZN(n1650) );
  OAI21_X4 U2638 ( .B1(n1651), .B2(net255325), .A(net255327), .ZN(net255107)
         );
  INV_X4 U2639 ( .A(net255329), .ZN(net255325) );
  INV_X4 U2640 ( .A(net255328), .ZN(n1651) );
  OAI21_X4 U2642 ( .B1(net255445), .B2(n1652), .A(net255327), .ZN(net255374)
         );
  NAND2_X2 U2643 ( .A1(net255329), .A2(net255328), .ZN(n1652) );
  NAND2_X2 U2644 ( .A1(n1655), .A2(net253043), .ZN(n1654) );
  AOI22_X2 U2646 ( .A1(net253049), .A2(net253050), .B1(n1660), .B2(n1661), 
        .ZN(n1659) );
  NAND2_X2 U2647 ( .A1(net253050), .A2(net256095), .ZN(n1661) );
  INV_X4 U2648 ( .A(net253049), .ZN(n1660) );
  NAND2_X2 U2649 ( .A1(n1660), .A2(net253050), .ZN(n1656) );
  NOR2_X4 U2651 ( .A1(n1662), .A2(n1656), .ZN(n1657) );
  INV_X4 U2652 ( .A(net253044), .ZN(n1662) );
  AOI22_X4 U2653 ( .A1(net253161), .A2(net253160), .B1(net253162), .B2(
        net253163), .ZN(net253038) );
  XNOR2_X2 U2654 ( .A(n1663), .B(net253193), .ZN(net253162) );
  NAND3_X2 U2655 ( .A1(n1664), .A2(net253198), .A3(net253192), .ZN(n1663) );
  NAND3_X2 U2656 ( .A1(net253059), .A2(net253058), .A3(net253208), .ZN(n1664)
         );
  INV_X4 U2657 ( .A(net256927), .ZN(net253058) );
  NOR2_X4 U2658 ( .A1(net253189), .A2(net253190), .ZN(net253160) );
  INV_X4 U2659 ( .A(net253163), .ZN(net253190) );
  INV_X4 U2660 ( .A(net253194), .ZN(net253189) );
  NAND2_X4 U2661 ( .A1(net254232), .A2(net254231), .ZN(net254142) );
  NOR2_X4 U2662 ( .A1(n1667), .A2(net254237), .ZN(net254231) );
  INV_X4 U2663 ( .A(net254238), .ZN(n1667) );
  NAND3_X2 U2664 ( .A1(net254233), .A2(net254234), .A3(net254235), .ZN(
        net254232) );
  NAND2_X4 U2665 ( .A1(net254147), .A2(n1665), .ZN(net254239) );
  XNOR2_X2 U2666 ( .A(net254298), .B(net254297), .ZN(n1665) );
  NAND2_X4 U2667 ( .A1(n1670), .A2(n1668), .ZN(net254145) );
  INV_X4 U2668 ( .A(net254285), .ZN(n1668) );
  INV_X8 U2669 ( .A(net254192), .ZN(n1666) );
  OAI21_X4 U2670 ( .B1(net254289), .B2(net254290), .A(net257254), .ZN(n1669)
         );
  OAI21_X2 U2671 ( .B1(net254289), .B2(net254290), .A(net257254), .ZN(
        net258069) );
  INV_X4 U2672 ( .A(net254147), .ZN(net254143) );
  NAND2_X4 U2673 ( .A1(n1672), .A2(net253685), .ZN(net253433) );
  NAND3_X2 U2674 ( .A1(net256741), .A2(net257980), .A3(net256982), .ZN(
        net253322) );
  AOI21_X2 U2675 ( .B1(net253688), .B2(net253689), .A(net253662), .ZN(
        net253690) );
  NAND2_X4 U2676 ( .A1(net253687), .A2(net253662), .ZN(n1672) );
  XNOR2_X2 U2677 ( .A(net253660), .B(net257981), .ZN(net253687) );
  XNOR2_X2 U2678 ( .A(net253660), .B(net257981), .ZN(net253659) );
  NAND2_X2 U2679 ( .A1(a[19]), .A2(net256165), .ZN(net253662) );
  INV_X4 U2680 ( .A(net253662), .ZN(net253656) );
  NAND2_X4 U2681 ( .A1(net253458), .A2(n1680), .ZN(n1679) );
  XNOR2_X2 U2682 ( .A(n1674), .B(n1673), .ZN(n1680) );
  INV_X4 U2683 ( .A(net253519), .ZN(n1671) );
  NOR3_X4 U2684 ( .A1(n1671), .A2(net253592), .A3(net253591), .ZN(net253584)
         );
  AND2_X2 U2685 ( .A1(n1603), .A2(n1675), .ZN(n1678) );
  NAND2_X4 U2686 ( .A1(net253701), .A2(n1675), .ZN(net253697) );
  NOR2_X4 U2687 ( .A1(net253756), .A2(net253445), .ZN(net253688) );
  INV_X2 U2688 ( .A(net255877), .ZN(net257564) );
  AOI222_X4 U2689 ( .A1(net255874), .A2(net256402), .B1(net255875), .B2(
        net257772), .C1(net255877), .C2(net257779), .ZN(net255870) );
  NAND3_X1 U2690 ( .A1(net256421), .A2(n1413), .A3(n1232), .ZN(net255964) );
  NAND3_X2 U2691 ( .A1(net253246), .A2(net256420), .A3(n1413), .ZN(net257779)
         );
  NAND3_X2 U2692 ( .A1(net253246), .A2(net256420), .A3(n1413), .ZN(net255540)
         );
  NAND2_X4 U2693 ( .A1(net256032), .A2(net256033), .ZN(net256421) );
  INV_X8 U2694 ( .A(net256421), .ZN(net256159) );
  INV_X8 U2695 ( .A(n1681), .ZN(net256033) );
  NAND2_X4 U2696 ( .A1(n1683), .A2(n1682), .ZN(n1681) );
  NAND3_X4 U2697 ( .A1(n1357), .A2(b[8]), .A3(control[1]), .ZN(n1683) );
  INV_X32 U2698 ( .A(control[0]), .ZN(net257678) );
  NAND3_X4 U2699 ( .A1(control[1]), .A2(control[0]), .A3(b[0]), .ZN(n1682) );
  INV_X8 U2700 ( .A(n1684), .ZN(net256032) );
  NAND2_X4 U2701 ( .A1(n1685), .A2(net256069), .ZN(n1684) );
  NAND3_X4 U2702 ( .A1(net257720), .A2(control[0]), .A3(b[16]), .ZN(net256069)
         );
  NAND2_X4 U2703 ( .A1(a[2]), .A2(n1466), .ZN(net256018) );
  NAND3_X4 U2704 ( .A1(n1467), .A2(b[18]), .A3(control[0]), .ZN(net256042) );
  NAND2_X4 U2705 ( .A1(net256054), .A2(net256055), .ZN(net256388) );
  INV_X8 U2706 ( .A(net256058), .ZN(net256055) );
  INV_X4 U2707 ( .A(net254414), .ZN(n1688) );
  INV_X4 U2708 ( .A(net254415), .ZN(n1687) );
  INV_X4 U2709 ( .A(net254634), .ZN(n1689) );
  NAND2_X4 U2710 ( .A1(n1690), .A2(n1689), .ZN(net254577) );
  INV_X4 U2711 ( .A(net256879), .ZN(n1690) );
  NAND2_X4 U2712 ( .A1(net254868), .A2(net257918), .ZN(net254941) );
  INV_X4 U2713 ( .A(net254935), .ZN(net257918) );
  INV_X4 U2714 ( .A(n1119), .ZN(net254935) );
  OAI21_X4 U2715 ( .B1(net255096), .B2(net254935), .A(net255097), .ZN(
        net255040) );
  NAND2_X4 U2716 ( .A1(n1697), .A2(net254867), .ZN(net254755) );
  NAND3_X2 U2717 ( .A1(net257953), .A2(n1118), .A3(net256555), .ZN(net254867)
         );
  NAND3_X2 U2718 ( .A1(net257953), .A2(net254869), .A3(net256555), .ZN(
        net256823) );
  NAND2_X4 U2719 ( .A1(net256555), .A2(net257392), .ZN(net256584) );
  INV_X8 U2720 ( .A(n1693), .ZN(n1697) );
  OAI21_X4 U2721 ( .B1(n1692), .B2(n1691), .A(n1694), .ZN(n1693) );
  XNOR2_X2 U2722 ( .A(n1695), .B(n1696), .ZN(n1694) );
  AOI21_X2 U2723 ( .B1(net255046), .B2(net255045), .A(net255044), .ZN(n1695)
         );
  NAND2_X4 U2724 ( .A1(net256796), .A2(n1691), .ZN(net254756) );
  XNOR2_X2 U2725 ( .A(net255047), .B(net256376), .ZN(n1692) );
  NAND2_X4 U2726 ( .A1(a[4]), .A2(net256119), .ZN(net255868) );
  INV_X32 U2727 ( .A(n1701), .ZN(net256119) );
  INV_X32 U2728 ( .A(n1701), .ZN(net256117) );
  INV_X4 U2729 ( .A(n1699), .ZN(n1698) );
  NOR3_X4 U2730 ( .A1(net256039), .A2(net256040), .A3(net256041), .ZN(n1699)
         );
  INV_X4 U2731 ( .A(net256042), .ZN(net256041) );
  NOR3_X4 U2732 ( .A1(n1700), .A2(control[0]), .A3(control[1]), .ZN(net256040)
         );
  INV_X4 U2733 ( .A(b[26]), .ZN(n1700) );
  NAND2_X2 U2734 ( .A1(net256044), .A2(net256045), .ZN(net256039) );
  NAND3_X4 U2735 ( .A1(control[1]), .A2(n1222), .A3(b[10]), .ZN(net256045) );
  NAND4_X4 U2736 ( .A1(n1333), .A2(control[1]), .A3(a[0]), .A4(b[9]), .ZN(
        net256050) );
  NAND3_X4 U2737 ( .A1(n1333), .A2(b[9]), .A3(control[1]), .ZN(net256060) );
  NAND3_X4 U2738 ( .A1(control[1]), .A2(control[0]), .A3(b[2]), .ZN(net256044)
         );
  NAND2_X4 U2739 ( .A1(net253688), .A2(net253689), .ZN(net253660) );
  INV_X4 U2740 ( .A(net253758), .ZN(net253756) );
  NAND3_X2 U2741 ( .A1(net253775), .A2(net253652), .A3(net253447), .ZN(
        net253758) );
  NAND2_X4 U2742 ( .A1(net253652), .A2(net253653), .ZN(net253448) );
  OAI21_X4 U2743 ( .B1(n1703), .B2(n1702), .A(net253800), .ZN(net253761) );
  NAND3_X2 U2744 ( .A1(net257439), .A2(n1704), .A3(net253801), .ZN(net253800)
         );
  INV_X4 U2745 ( .A(net253983), .ZN(n1704) );
  NAND3_X2 U2746 ( .A1(net253802), .A2(net253801), .A3(n1704), .ZN(net253646)
         );
  NOR2_X4 U2747 ( .A1(net253805), .A2(net253806), .ZN(n1702) );
  INV_X4 U2748 ( .A(net254085), .ZN(net253806) );
  OAI21_X1 U2749 ( .B1(net253824), .B2(net256362), .A(net253806), .ZN(
        net254083) );
  NAND2_X4 U2750 ( .A1(n1706), .A2(net253780), .ZN(net253650) );
  NAND2_X4 U2751 ( .A1(net253808), .A2(net253650), .ZN(net256375) );
  NAND3_X2 U2752 ( .A1(net253986), .A2(net253987), .A3(n1707), .ZN(net253801)
         );
  INV_X4 U2753 ( .A(net253801), .ZN(net253985) );
  NAND2_X4 U2754 ( .A1(net253824), .A2(n1707), .ZN(net253823) );
  OAI21_X4 U2755 ( .B1(n1708), .B2(net253988), .A(n1492), .ZN(net257439) );
  OAI21_X2 U2756 ( .B1(n1708), .B2(net253988), .A(n1492), .ZN(net253802) );
  INV_X4 U2757 ( .A(net253987), .ZN(net253988) );
  INV_X4 U2758 ( .A(net253986), .ZN(n1708) );
  NAND2_X2 U2759 ( .A1(a[18]), .A2(net256173), .ZN(net253983) );
  OAI21_X4 U2760 ( .B1(net253984), .B2(net253985), .A(net253983), .ZN(
        net253647) );
  OAI21_X4 U2761 ( .B1(n1262), .B2(net253422), .A(net253423), .ZN(net253205)
         );
  OAI22_X4 U2762 ( .A1(net253424), .A2(net253425), .B1(net253424), .B2(n1712), 
        .ZN(net253423) );
  INV_X4 U2763 ( .A(n1712), .ZN(net256800) );
  FA_X1 U2764 ( .A(net253582), .B(net253583), .CI(net253451), .S(n1709) );
  XOR2_X2 U2765 ( .A(net253441), .B(n1417), .Z(net253583) );
  NAND2_X4 U2766 ( .A1(net253427), .A2(n1417), .ZN(net253414) );
  INV_X4 U2767 ( .A(net253450), .ZN(net253441) );
  NAND2_X4 U2768 ( .A1(net253442), .A2(net253441), .ZN(net253398) );
  INV_X4 U2769 ( .A(net253452), .ZN(net253582) );
  OAI21_X2 U2770 ( .B1(n1711), .B2(n1710), .A(net257442), .ZN(net253580) );
  INV_X4 U2771 ( .A(net257796), .ZN(net253641) );
  NAND2_X4 U2772 ( .A1(net253640), .A2(net253641), .ZN(net253323) );
  XNOR2_X2 U2773 ( .A(n1167), .B(net253694), .ZN(net257796) );
  INV_X4 U2774 ( .A(net253643), .ZN(net253640) );
  OAI21_X2 U2775 ( .B1(n1421), .B2(net253457), .A(net253458), .ZN(n1711) );
  AOI21_X2 U2776 ( .B1(net257828), .B2(net253448), .A(net253651), .ZN(n1710)
         );
  INV_X4 U2777 ( .A(n1108), .ZN(net253651) );
  NOR2_X2 U2778 ( .A1(net253651), .A2(net253445), .ZN(net253770) );
  NAND2_X4 U2779 ( .A1(net255619), .A2(net255618), .ZN(net255431) );
  NAND2_X2 U2780 ( .A1(net257240), .A2(net255431), .ZN(net255617) );
  XNOR2_X2 U2781 ( .A(net255708), .B(n1345), .ZN(n1713) );
  NAND3_X4 U2782 ( .A1(net255726), .A2(net255727), .A3(n1714), .ZN(net255434)
         );
  INV_X4 U2783 ( .A(net255775), .ZN(n1714) );
  INV_X8 U2784 ( .A(net256990), .ZN(net257363) );
  NOR3_X4 U2785 ( .A1(net255441), .A2(net255442), .A3(net257363), .ZN(
        net255435) );
  INV_X8 U2786 ( .A(net255443), .ZN(net256990) );
  NAND3_X2 U2787 ( .A1(net255221), .A2(net256990), .A3(net257522), .ZN(
        net255089) );
  NAND3_X2 U2788 ( .A1(net255221), .A2(net257522), .A3(net256990), .ZN(
        net255320) );
  AOI211_X4 U2789 ( .C1(net253179), .C2(net253178), .A(net253180), .B(n1715), 
        .ZN(net253164) );
  INV_X4 U2790 ( .A(net253183), .ZN(n1717) );
  INV_X8 U2791 ( .A(net253291), .ZN(net253180) );
  INV_X4 U2792 ( .A(net253180), .ZN(net257211) );
  OR2_X4 U2793 ( .A1(net253180), .A2(net257159), .ZN(net253553) );
  NAND2_X4 U2794 ( .A1(net253564), .A2(net253533), .ZN(net253291) );
  NOR2_X4 U2795 ( .A1(net253185), .A2(net253188), .ZN(net253178) );
  OAI21_X4 U2796 ( .B1(net254942), .B2(net256584), .A(n1718), .ZN(net254868)
         );
  OAI22_X4 U2797 ( .A1(net255226), .A2(net256556), .B1(net254942), .B2(
        net256584), .ZN(net255164) );
  NAND2_X4 U2798 ( .A1(net255100), .A2(net255099), .ZN(net254869) );
  OAI21_X2 U2799 ( .B1(net255099), .B2(net255100), .A(net255101), .ZN(
        net255098) );
  INV_X4 U2800 ( .A(net255167), .ZN(net255099) );
  NAND2_X2 U2801 ( .A1(n1718), .A2(net254869), .ZN(net255165) );
  NAND3_X2 U2802 ( .A1(net253765), .A2(n1721), .A3(n1719), .ZN(net253775) );
  INV_X8 U2803 ( .A(n1720), .ZN(n1719) );
  NAND3_X2 U2804 ( .A1(n1122), .A2(n1719), .A3(n1721), .ZN(net254054) );
  INV_X1 U2805 ( .A(n1719), .ZN(net256334) );
  NAND3_X2 U2806 ( .A1(net253797), .A2(n1719), .A3(n1721), .ZN(net253653) );
  NAND2_X4 U2807 ( .A1(net257069), .A2(net254057), .ZN(n1720) );
  NAND2_X4 U2808 ( .A1(net253765), .A2(n1721), .ZN(net254179) );
  OAI21_X4 U2809 ( .B1(net253305), .B2(net256095), .A(net253306), .ZN(
        net253169) );
  NAND2_X2 U2810 ( .A1(net253169), .A2(net253194), .ZN(net253286) );
  INV_X4 U2811 ( .A(product_in[29]), .ZN(n1724) );
  OAI21_X4 U2812 ( .B1(n1722), .B2(net253278), .A(n1725), .ZN(net253316) );
  XNOR2_X2 U2813 ( .A(n1726), .B(n1727), .ZN(n1725) );
  OAI21_X2 U2814 ( .B1(n1728), .B2(net253320), .A(n1722), .ZN(n1727) );
  INV_X4 U2815 ( .A(net253280), .ZN(n1722) );
  NOR2_X4 U2816 ( .A1(net253278), .A2(n1722), .ZN(net256927) );
  NAND2_X2 U2817 ( .A1(n1722), .A2(net253327), .ZN(n1726) );
  AOI21_X1 U2818 ( .B1(net253322), .B2(net257153), .A(net253324), .ZN(n1728)
         );
  INV_X4 U2819 ( .A(net253396), .ZN(net253324) );
  NOR2_X2 U2820 ( .A1(net253322), .A2(net253324), .ZN(net253392) );
  INV_X8 U2821 ( .A(net257442), .ZN(net253395) );
  NAND2_X2 U2822 ( .A1(net253395), .A2(n1290), .ZN(net253394) );
  OAI21_X4 U2823 ( .B1(net256982), .B2(net253395), .A(net253431), .ZN(
        net253429) );
  INV_X8 U2824 ( .A(net255439), .ZN(net255548) );
  NAND2_X4 U2825 ( .A1(net255547), .A2(net255548), .ZN(net255220) );
  NAND2_X4 U2826 ( .A1(net255548), .A2(net255547), .ZN(net257522) );
  INV_X4 U2827 ( .A(net255438), .ZN(net255547) );
  NAND2_X4 U2828 ( .A1(net256747), .A2(net255547), .ZN(net255585) );
  OAI21_X4 U2829 ( .B1(net255588), .B2(net255589), .A(net255590), .ZN(
        net255584) );
  XNOR2_X2 U2830 ( .A(net255584), .B(net255585), .ZN(net257481) );
  NOR3_X2 U2831 ( .A1(n1729), .A2(net255438), .A3(n1732), .ZN(net255589) );
  INV_X8 U2832 ( .A(n1730), .ZN(n1732) );
  NOR2_X4 U2833 ( .A1(n1729), .A2(n1732), .ZN(net255429) );
  INV_X8 U2834 ( .A(net255433), .ZN(n1730) );
  NAND2_X2 U2835 ( .A1(n1730), .A2(net255591), .ZN(net255543) );
  XNOR2_X2 U2836 ( .A(net255773), .B(n1730), .ZN(net256290) );
  INV_X4 U2837 ( .A(net255591), .ZN(n1729) );
  NAND2_X4 U2838 ( .A1(n1731), .A2(net256748), .ZN(net255439) );
  CLKBUF_X3 U2839 ( .A(net255439), .Z(net257560) );
  NAND2_X4 U2840 ( .A1(net256746), .A2(net256747), .ZN(n1731) );
  INV_X4 U2841 ( .A(net255594), .ZN(net256746) );
  NAND2_X2 U2842 ( .A1(net255594), .A2(net255587), .ZN(net256748) );
  NAND2_X2 U2843 ( .A1(a[6]), .A2(net256137), .ZN(net255438) );
  NAND2_X4 U2844 ( .A1(net256060), .A2(net256059), .ZN(net256058) );
  NAND3_X4 U2845 ( .A1(control[1]), .A2(control[0]), .A3(b[1]), .ZN(net256059)
         );
  NAND2_X4 U2846 ( .A1(net255706), .A2(n1733), .ZN(net255427) );
  NAND2_X4 U2847 ( .A1(net257485), .A2(net255427), .ZN(net255179) );
  INV_X4 U2848 ( .A(n1734), .ZN(n1733) );
  XNOR2_X2 U2849 ( .A(net255708), .B(n1345), .ZN(n1734) );
  INV_X4 U2850 ( .A(net255624), .ZN(net255706) );
  XNOR2_X2 U2851 ( .A(net254635), .B(n1419), .ZN(net256879) );
  XNOR2_X2 U2852 ( .A(net254635), .B(n1419), .ZN(net254633) );
  NOR2_X4 U2853 ( .A1(n1585), .A2(n1270), .ZN(net254693) );
  INV_X4 U2854 ( .A(net254947), .ZN(net257392) );
  NAND2_X4 U2855 ( .A1(net256627), .A2(net257392), .ZN(net255284) );
  INV_X8 U2856 ( .A(net255229), .ZN(net254947) );
  OAI22_X4 U2857 ( .A1(net255105), .A2(net254947), .B1(net255106), .B2(
        net254947), .ZN(net255104) );
  NAND2_X2 U2858 ( .A1(net254051), .A2(net256541), .ZN(net253987) );
  NAND2_X2 U2859 ( .A1(net254463), .A2(net254462), .ZN(net254461) );
  NAND2_X4 U2860 ( .A1(net254673), .A2(n1735), .ZN(net254462) );
  XNOR2_X2 U2861 ( .A(n1736), .B(n1737), .ZN(n1735) );
  NAND3_X1 U2862 ( .A1(net254562), .A2(n1111), .A3(net254760), .ZN(n1737) );
  INV_X2 U2863 ( .A(n1738), .ZN(n1739) );
  INV_X1 U2864 ( .A(net254761), .ZN(n1738) );
  NAND2_X2 U2865 ( .A1(net254952), .A2(net254760), .ZN(net254864) );
  INV_X4 U2866 ( .A(net254760), .ZN(net254683) );
  INV_X4 U2867 ( .A(net254858), .ZN(n1740) );
  NAND2_X2 U2868 ( .A1(net255433), .A2(net257752), .ZN(net255724) );
  OAI21_X4 U2869 ( .B1(net255616), .B2(net255593), .A(net255617), .ZN(
        net255594) );
  INV_X8 U2870 ( .A(net255910), .ZN(net257772) );
  INV_X2 U2871 ( .A(net253424), .ZN(net257435) );
  INV_X4 U2872 ( .A(n1743), .ZN(n1742) );
  XNOR2_X2 U2873 ( .A(net253579), .B(net256800), .ZN(net253572) );
  NAND3_X2 U2874 ( .A1(net257031), .A2(net258007), .A3(n1744), .ZN(net253689)
         );
  NAND2_X1 U2875 ( .A1(net253647), .A2(net257109), .ZN(n1744) );
  OAI21_X4 U2876 ( .B1(net253446), .B2(net253445), .A(net257031), .ZN(
        net256982) );
  OAI21_X2 U2877 ( .B1(net253445), .B2(net253446), .A(net257031), .ZN(
        net253402) );
  OAI21_X4 U2878 ( .B1(n1422), .B2(n1745), .A(net253394), .ZN(net253393) );
  NAND2_X4 U2880 ( .A1(n1747), .A2(net253401), .ZN(net253156) );
  XNOR2_X2 U2881 ( .A(net253462), .B(net253463), .ZN(n1748) );
  INV_X4 U2882 ( .A(net255538), .ZN(net255537) );
  NAND2_X2 U2883 ( .A1(net255538), .A2(net256909), .ZN(net255606) );
  OAI21_X4 U2884 ( .B1(net256958), .B2(net255624), .A(net257752), .ZN(
        net255593) );
  INV_X8 U2885 ( .A(net255533), .ZN(net255714) );
  INV_X8 U2886 ( .A(net255219), .ZN(net255443) );
  INV_X8 U2887 ( .A(net255220), .ZN(net255442) );
  NAND2_X4 U2888 ( .A1(net255322), .A2(net257456), .ZN(net255221) );
  NAND2_X4 U2889 ( .A1(n1750), .A2(n1749), .ZN(net255219) );
  NAND2_X4 U2890 ( .A1(net255219), .A2(net255629), .ZN(net255699) );
  INV_X4 U2891 ( .A(net255703), .ZN(n1749) );
  INV_X2 U2892 ( .A(net255702), .ZN(n1750) );
  INV_X4 U2893 ( .A(net254184), .ZN(n1752) );
  NAND2_X2 U2894 ( .A1(a[17]), .A2(net256105), .ZN(n1751) );
  INV_X16 U2895 ( .A(net253103), .ZN(net256115) );
  OAI21_X4 U2896 ( .B1(net255435), .B2(net255436), .A(net256296), .ZN(
        net255380) );
  XNOR2_X2 U2897 ( .A(n1415), .B(n3998), .ZN(n3981) );
  INV_X2 U2898 ( .A(n3177), .ZN(n1995) );
  NAND2_X2 U2899 ( .A1(net254669), .A2(n1834), .ZN(n1753) );
  CLKBUF_X2 U2900 ( .A(n3547), .Z(n1754) );
  NAND2_X2 U2901 ( .A1(n3348), .A2(n3453), .ZN(n3547) );
  INV_X2 U2902 ( .A(n2848), .ZN(n2870) );
  INV_X4 U2903 ( .A(n1247), .ZN(n2743) );
  NAND2_X4 U2904 ( .A1(n2543), .A2(n1409), .ZN(n2659) );
  XNOR2_X2 U2905 ( .A(net255699), .B(n2258), .ZN(n1755) );
  CLKBUF_X3 U2906 ( .A(n3899), .Z(n1756) );
  NAND2_X4 U2907 ( .A1(n2498), .A2(n1926), .ZN(n2548) );
  XNOR2_X1 U2909 ( .A(n3998), .B(n4003), .ZN(n3999) );
  NOR3_X2 U2910 ( .A1(n4003), .A2(n4002), .A3(n4008), .ZN(n4064) );
  OAI21_X2 U2911 ( .B1(net257239), .B2(n3453), .A(net257296), .ZN(net254191)
         );
  NAND2_X2 U2912 ( .A1(n3455), .A2(n3249), .ZN(net254290) );
  INV_X2 U2913 ( .A(n4001), .ZN(n4008) );
  INV_X1 U2915 ( .A(n3498), .ZN(n1758) );
  NAND3_X2 U2917 ( .A1(n3462), .A2(n3461), .A3(n3460), .ZN(n1760) );
  XNOR2_X1 U2918 ( .A(n4088), .B(n1892), .ZN(net258044) );
  OAI21_X4 U2919 ( .B1(n2372), .B2(net255714), .A(n2371), .ZN(n2373) );
  INV_X8 U2920 ( .A(n3507), .ZN(n3786) );
  INV_X4 U2921 ( .A(n2325), .ZN(n2376) );
  INV_X4 U2922 ( .A(n3278), .ZN(n3160) );
  XNOR2_X2 U2923 ( .A(n2709), .B(n2758), .ZN(n1762) );
  NAND2_X4 U2924 ( .A1(n2342), .A2(n2343), .ZN(n2496) );
  AOI21_X4 U2926 ( .B1(n2273), .B2(n2426), .A(n2272), .ZN(n2274) );
  NAND2_X4 U2927 ( .A1(n3603), .A2(n1790), .ZN(n3605) );
  INV_X4 U2928 ( .A(n4103), .ZN(n1764) );
  NAND2_X4 U2929 ( .A1(n2624), .A2(n2625), .ZN(n2744) );
  NAND2_X2 U2930 ( .A1(n2625), .A2(n2624), .ZN(n1894) );
  INV_X8 U2931 ( .A(n2448), .ZN(n2513) );
  NAND2_X2 U2932 ( .A1(a[11]), .A2(n3955), .ZN(n2448) );
  NAND2_X2 U2933 ( .A1(n1903), .A2(n3377), .ZN(n1765) );
  INV_X4 U2934 ( .A(n1920), .ZN(n1859) );
  NAND2_X4 U2935 ( .A1(n2923), .A2(n2924), .ZN(n1766) );
  XNOR2_X2 U2936 ( .A(n2980), .B(n1966), .ZN(n1767) );
  NAND2_X4 U2937 ( .A1(n2963), .A2(n3196), .ZN(n2980) );
  NAND2_X2 U2938 ( .A1(n1449), .A2(n1834), .ZN(net254873) );
  XNOR2_X1 U2939 ( .A(n2376), .B(n2435), .ZN(n1768) );
  NAND2_X2 U2940 ( .A1(n3919), .A2(net253177), .ZN(n3861) );
  OAI21_X2 U2941 ( .B1(net255790), .B2(n2199), .A(net256402), .ZN(n1770) );
  INV_X8 U2943 ( .A(n3551), .ZN(n3677) );
  NAND2_X4 U2944 ( .A1(n4087), .A2(n1593), .ZN(n3342) );
  NAND2_X4 U2945 ( .A1(n3938), .A2(n3934), .ZN(net253463) );
  XNOR2_X2 U2946 ( .A(n3904), .B(n3903), .ZN(n1871) );
  NAND2_X2 U2947 ( .A1(n1844), .A2(n3437), .ZN(n3322) );
  NAND2_X4 U2948 ( .A1(n3442), .A2(n3635), .ZN(n3321) );
  INV_X2 U2949 ( .A(net255089), .ZN(net255218) );
  NAND2_X4 U2950 ( .A1(n2629), .A2(n2535), .ZN(n2396) );
  XNOR2_X2 U2951 ( .A(n3945), .B(n3903), .ZN(n1772) );
  NAND2_X4 U2952 ( .A1(n3896), .A2(n3944), .ZN(n3945) );
  INV_X4 U2953 ( .A(n2393), .ZN(n1890) );
  NOR2_X2 U2954 ( .A1(n3596), .A2(n3598), .ZN(n3600) );
  OAI221_X4 U2955 ( .B1(n3512), .B2(n3918), .C1(n3917), .C2(net256095), .A(
        n3259), .ZN(n1832) );
  INV_X2 U2956 ( .A(n1317), .ZN(n3546) );
  INV_X4 U2957 ( .A(n3093), .ZN(n3099) );
  NOR2_X4 U2958 ( .A1(n3758), .A2(n1909), .ZN(net253810) );
  INV_X2 U2959 ( .A(n2989), .ZN(n1911) );
  XNOR2_X1 U2960 ( .A(n2971), .B(n1775), .ZN(n1837) );
  NAND2_X2 U2961 ( .A1(n3243), .A2(n1791), .ZN(n3249) );
  NOR2_X2 U2962 ( .A1(n2222), .A2(n2221), .ZN(n2233) );
  NAND2_X4 U2963 ( .A1(n2138), .A2(n2221), .ZN(n3918) );
  NAND2_X4 U2964 ( .A1(n2137), .A2(n2136), .ZN(n2221) );
  OAI22_X2 U2965 ( .A1(n1619), .A2(n3707), .B1(net253656), .B2(net253657), 
        .ZN(net253579) );
  NAND2_X4 U2966 ( .A1(n2157), .A2(n1795), .ZN(n2158) );
  NAND2_X1 U2967 ( .A1(n1895), .A2(n3019), .ZN(n1778) );
  NAND2_X4 U2968 ( .A1(net253764), .A2(n3252), .ZN(n3388) );
  INV_X8 U2969 ( .A(n3155), .ZN(n3285) );
  OAI221_X4 U2970 ( .B1(net253308), .B2(n3410), .C1(n3409), .C2(net256184), 
        .A(n3408), .ZN(n3507) );
  INV_X2 U2971 ( .A(n2706), .ZN(n2704) );
  INV_X1 U2972 ( .A(n4096), .ZN(n1780) );
  NAND3_X1 U2974 ( .A1(net256420), .A2(net253246), .A3(net255872), .ZN(n1781)
         );
  NAND3_X2 U2975 ( .A1(net256420), .A2(net253246), .A3(net255872), .ZN(n2442)
         );
  BUF_X32 U2976 ( .A(n3625), .Z(n1782) );
  NAND2_X4 U2977 ( .A1(n1825), .A2(n3252), .ZN(n3279) );
  NAND2_X4 U2978 ( .A1(n1350), .A2(net253398), .ZN(n1783) );
  NAND2_X4 U2979 ( .A1(n3075), .A2(n3074), .ZN(n3174) );
  NAND3_X2 U2980 ( .A1(n3503), .A2(n3502), .A3(n3501), .ZN(n1785) );
  NAND2_X4 U2981 ( .A1(n1956), .A2(n3337), .ZN(n3503) );
  OAI221_X4 U2982 ( .B1(n3512), .B2(n3918), .C1(n3917), .C2(net256095), .A(
        n3259), .ZN(n3261) );
  NOR2_X4 U2983 ( .A1(n3758), .A2(net253586), .ZN(net257838) );
  NAND2_X4 U2984 ( .A1(n1762), .A2(n2710), .ZN(n1786) );
  NAND2_X2 U2985 ( .A1(n3077), .A2(n3076), .ZN(n1787) );
  NAND2_X1 U2986 ( .A1(net253287), .A2(net253177), .ZN(n3921) );
  NAND2_X4 U2987 ( .A1(b[25]), .A2(net257720), .ZN(n2032) );
  INV_X8 U2988 ( .A(n3552), .ZN(n1790) );
  INV_X8 U2989 ( .A(n3602), .ZN(n3552) );
  XNOR2_X1 U2990 ( .A(n3149), .B(n3150), .ZN(n1791) );
  NAND2_X4 U2991 ( .A1(n3291), .A2(n3203), .ZN(n3150) );
  NAND3_X2 U2992 ( .A1(n3196), .A2(n3197), .A3(n3193), .ZN(n3036) );
  NAND2_X2 U2993 ( .A1(net253386), .A2(net253519), .ZN(net253694) );
  NAND2_X4 U2994 ( .A1(b[16]), .A2(control[0]), .ZN(n2036) );
  XNOR2_X2 U2995 ( .A(n2075), .B(net257565), .ZN(n1793) );
  INV_X1 U2996 ( .A(n2765), .ZN(n2767) );
  NAND2_X4 U2997 ( .A1(n2439), .A2(net255409), .ZN(net255538) );
  NAND2_X4 U2998 ( .A1(n3157), .A2(n3156), .ZN(n3155) );
  INV_X4 U2999 ( .A(n1874), .ZN(n2450) );
  NAND2_X4 U3000 ( .A1(a[3]), .A2(net256371), .ZN(n2039) );
  INV_X16 U3001 ( .A(control[0]), .ZN(net256371) );
  INV_X2 U3002 ( .A(n2189), .ZN(n1795) );
  NAND4_X4 U3003 ( .A1(b[9]), .A2(n1221), .A3(a[2]), .A4(control[1]), .ZN(
        n2061) );
  NAND2_X2 U3004 ( .A1(n3630), .A2(net253646), .ZN(n3614) );
  NAND2_X4 U3005 ( .A1(n3578), .A2(n3577), .ZN(n3660) );
  INV_X4 U3006 ( .A(n3993), .ZN(n3994) );
  NAND2_X4 U3007 ( .A1(n2463), .A2(n2462), .ZN(n1796) );
  NAND2_X2 U3008 ( .A1(n2463), .A2(n2462), .ZN(n2613) );
  INV_X8 U3009 ( .A(n2119), .ZN(n2122) );
  NAND2_X4 U3010 ( .A1(n1981), .A2(control[1]), .ZN(n2034) );
  NAND2_X4 U3011 ( .A1(a[2]), .A2(n1332), .ZN(n2033) );
  INV_X16 U3012 ( .A(control[0]), .ZN(net256087) );
  INV_X8 U3013 ( .A(n3235), .ZN(n3428) );
  XNOR2_X2 U3014 ( .A(n3589), .B(n3588), .ZN(n1797) );
  NAND2_X4 U3015 ( .A1(n2519), .A2(n2520), .ZN(n2521) );
  NOR2_X2 U3016 ( .A1(net256334), .A2(n3532), .ZN(n3528) );
  INV_X8 U3017 ( .A(n1860), .ZN(n1799) );
  NAND2_X4 U3018 ( .A1(n1943), .A2(n3493), .ZN(n3506) );
  OAI21_X2 U3019 ( .B1(n3147), .B2(n3148), .A(n1206), .ZN(n1801) );
  INV_X8 U3020 ( .A(n3505), .ZN(n3787) );
  INV_X4 U3021 ( .A(n1804), .ZN(n1805) );
  INV_X4 U3022 ( .A(n2056), .ZN(n2057) );
  XNOR2_X1 U3023 ( .A(n3005), .B(n3003), .ZN(product_out[18]) );
  AND4_X4 U3024 ( .A1(n2443), .A2(net256402), .A3(n1840), .A4(net255409), .ZN(
        n2444) );
  NAND3_X2 U3025 ( .A1(n2420), .A2(n2421), .A3(n2419), .ZN(n2495) );
  INV_X2 U3026 ( .A(n3584), .ZN(n1806) );
  NAND2_X1 U3027 ( .A1(net256306), .A2(net254761), .ZN(n1866) );
  XNOR2_X2 U3028 ( .A(n2123), .B(n1998), .ZN(n1807) );
  NAND2_X4 U3030 ( .A1(n2564), .A2(n2644), .ZN(n2645) );
  OAI211_X4 U3031 ( .C1(n3169), .C2(net256095), .A(net255247), .B(n2562), .ZN(
        n2564) );
  NAND4_X4 U3032 ( .A1(b[1]), .A2(control[1]), .A3(a[2]), .A4(control[0]), 
        .ZN(n1808) );
  NAND2_X4 U3033 ( .A1(b[17]), .A2(control[0]), .ZN(n2031) );
  NOR3_X2 U3034 ( .A1(n3771), .A2(net253557), .A3(n3774), .ZN(n3772) );
  NAND2_X4 U3035 ( .A1(n3563), .A2(n3637), .ZN(n3379) );
  NAND2_X4 U3036 ( .A1(n3377), .A2(n1903), .ZN(n3378) );
  OAI21_X4 U3037 ( .B1(n3030), .B2(net254566), .A(n1374), .ZN(n1810) );
  NAND2_X4 U3038 ( .A1(n1965), .A2(n2981), .ZN(net254464) );
  INV_X4 U3039 ( .A(net257211), .ZN(net257672) );
  INV_X2 U3040 ( .A(net253402), .ZN(net253444) );
  NOR2_X2 U3041 ( .A1(net253913), .A2(n3532), .ZN(n3527) );
  NAND2_X4 U3042 ( .A1(net254255), .A2(n3277), .ZN(n3252) );
  NOR2_X4 U3043 ( .A1(n1812), .A2(n1409), .ZN(n1811) );
  XNOR2_X2 U3044 ( .A(n2542), .B(n2541), .ZN(n1812) );
  NOR2_X2 U3045 ( .A1(n3100), .A2(n3101), .ZN(n3103) );
  NOR2_X4 U3046 ( .A1(net253209), .A2(n1924), .ZN(net253208) );
  NAND2_X2 U3047 ( .A1(n1756), .A2(n3900), .ZN(n3940) );
  NOR2_X2 U3048 ( .A1(n3941), .A2(n3898), .ZN(n3902) );
  INV_X4 U3049 ( .A(net253220), .ZN(net257650) );
  INV_X4 U3050 ( .A(net253156), .ZN(net253220) );
  INV_X4 U3051 ( .A(n1960), .ZN(n3136) );
  CLKBUF_X2 U3052 ( .A(n2194), .Z(n1815) );
  OAI21_X4 U3053 ( .B1(net253273), .B2(net253274), .A(n3933), .ZN(net253059)
         );
  INV_X4 U3054 ( .A(net253936), .ZN(net257630) );
  INV_X2 U3055 ( .A(net253182), .ZN(net253936) );
  NAND2_X4 U3056 ( .A1(n1390), .A2(net256127), .ZN(n2224) );
  INV_X2 U3057 ( .A(n2265), .ZN(n2127) );
  INV_X2 U3058 ( .A(n3520), .ZN(n3521) );
  INV_X8 U3059 ( .A(n2860), .ZN(n2861) );
  NOR3_X1 U3060 ( .A1(n4090), .A2(n3767), .A3(n3769), .ZN(n3779) );
  NAND2_X4 U3061 ( .A1(n2191), .A2(n2190), .ZN(n1818) );
  INV_X4 U3062 ( .A(net257481), .ZN(net255437) );
  NAND2_X1 U3063 ( .A1(n2018), .A2(n2059), .ZN(n2019) );
  NAND2_X2 U3064 ( .A1(n3008), .A2(n3007), .ZN(n3009) );
  INV_X2 U3065 ( .A(n2344), .ZN(n2342) );
  INV_X1 U3066 ( .A(n2431), .ZN(n1819) );
  INV_X2 U3067 ( .A(net257589), .ZN(net257590) );
  NAND3_X2 U3068 ( .A1(net255725), .A2(net257752), .A3(n1258), .ZN(n2247) );
  NAND2_X4 U3069 ( .A1(n3593), .A2(n3592), .ZN(n3680) );
  NAND2_X2 U3070 ( .A1(n2122), .A2(n2121), .ZN(n1820) );
  INV_X4 U3071 ( .A(n1793), .ZN(n2121) );
  NAND2_X4 U3072 ( .A1(n2867), .A2(n1301), .ZN(n2807) );
  OAI21_X2 U3073 ( .B1(n2059), .B2(n2060), .A(n2190), .ZN(n2078) );
  NAND2_X2 U3074 ( .A1(net256527), .A2(net256843), .ZN(n2110) );
  INV_X4 U3075 ( .A(net256843), .ZN(net255779) );
  INV_X2 U3076 ( .A(n1455), .ZN(n3018) );
  AOI21_X2 U3077 ( .B1(n3484), .B2(n3485), .A(n3483), .ZN(n3491) );
  INV_X4 U3078 ( .A(net255231), .ZN(n1947) );
  NAND2_X4 U3079 ( .A1(net255231), .A2(net255232), .ZN(net255101) );
  INV_X8 U3080 ( .A(net255434), .ZN(net255428) );
  NAND2_X4 U3081 ( .A1(n3661), .A2(n3660), .ZN(n3722) );
  XNOR2_X2 U3082 ( .A(n2709), .B(n1836), .ZN(n1823) );
  INV_X4 U3083 ( .A(n2964), .ZN(n2965) );
  CLKBUF_X3 U3084 ( .A(n2279), .Z(n1824) );
  NOR2_X2 U3085 ( .A1(n1768), .A2(n2329), .ZN(n2332) );
  AND2_X4 U3086 ( .A1(net255606), .A2(n1768), .ZN(n2326) );
  OAI211_X2 U3087 ( .C1(n2370), .C2(n2369), .A(n1982), .B(net255537), .ZN(
        n2374) );
  NAND2_X4 U3088 ( .A1(n2178), .A2(n2292), .ZN(n2179) );
  NAND2_X4 U3089 ( .A1(n2177), .A2(n2176), .ZN(n2292) );
  NAND2_X4 U3090 ( .A1(n3159), .A2(n3158), .ZN(n1825) );
  XOR2_X1 U3091 ( .A(n3876), .B(n3825), .Z(n1826) );
  INV_X1 U3092 ( .A(n1327), .ZN(n2097) );
  INV_X2 U3093 ( .A(n3894), .ZN(n3892) );
  INV_X8 U3094 ( .A(net253205), .ZN(net253273) );
  NAND2_X2 U3095 ( .A1(n2125), .A2(n1863), .ZN(n2129) );
  OAI221_X4 U3096 ( .B1(n1807), .B2(n2189), .C1(n2188), .C2(n2159), .A(n2187), 
        .ZN(n1829) );
  OAI221_X2 U3097 ( .B1(n1807), .B2(n2189), .C1(n2188), .C2(n2159), .A(n2187), 
        .ZN(n2321) );
  NAND2_X4 U3098 ( .A1(n1444), .A2(n2185), .ZN(n2159) );
  NAND3_X2 U3099 ( .A1(a[22]), .A2(n3425), .A3(net256117), .ZN(n1830) );
  CLKBUF_X3 U3100 ( .A(net254057), .Z(net257407) );
  NAND2_X4 U3101 ( .A1(n2283), .A2(n2282), .ZN(n2284) );
  NAND2_X2 U3102 ( .A1(net255425), .A2(n1873), .ZN(n2433) );
  INV_X2 U3103 ( .A(net255179), .ZN(net255425) );
  NAND2_X2 U3104 ( .A1(net254562), .A2(n1111), .ZN(n2786) );
  NAND2_X4 U3105 ( .A1(n2782), .A2(n2783), .ZN(net254562) );
  INV_X4 U3106 ( .A(net255426), .ZN(net257484) );
  OAI22_X4 U3107 ( .A1(n2281), .A2(n2235), .B1(n1827), .B2(n2234), .ZN(n2237)
         );
  OAI22_X4 U3108 ( .A1(net256145), .A2(n2248), .B1(n2072), .B2(n2434), .ZN(
        n2439) );
  NAND3_X2 U3109 ( .A1(n2321), .A2(n2320), .A3(n2319), .ZN(n2245) );
  INV_X1 U3110 ( .A(n3898), .ZN(n1833) );
  OAI21_X4 U3111 ( .B1(net256139), .B2(n2839), .A(n2838), .ZN(n1834) );
  NAND3_X2 U3112 ( .A1(net255916), .A2(net257401), .A3(net255915), .ZN(n1835)
         );
  NAND2_X4 U3113 ( .A1(n2318), .A2(n1764), .ZN(n2365) );
  NAND2_X4 U3114 ( .A1(n2967), .A2(n3046), .ZN(n2971) );
  OAI21_X2 U3115 ( .B1(n2970), .B2(n2969), .A(n3045), .ZN(n3047) );
  XNOR2_X1 U3116 ( .A(n1153), .B(n2640), .ZN(n3915) );
  NOR2_X4 U3117 ( .A1(n2750), .A2(n2751), .ZN(n1838) );
  NAND2_X1 U3118 ( .A1(a[10]), .A2(net256135), .ZN(n2618) );
  NAND4_X1 U3119 ( .A1(n2699), .A2(n2449), .A3(n2700), .A4(n2452), .ZN(n2459)
         );
  NAND2_X4 U3120 ( .A1(n2303), .A2(n2302), .ZN(n2416) );
  XNOR2_X1 U3121 ( .A(n2301), .B(n2302), .ZN(product_out[8]) );
  OAI22_X4 U3122 ( .A1(net256184), .A2(n3410), .B1(n3406), .B2(net256095), 
        .ZN(n2302) );
  INV_X2 U3123 ( .A(net253815), .ZN(net257171) );
  XNOR2_X2 U3124 ( .A(n3700), .B(net256966), .ZN(product_out[26]) );
  INV_X8 U3125 ( .A(n2372), .ZN(n1840) );
  INV_X8 U3126 ( .A(n2442), .ZN(n2372) );
  NAND2_X1 U3128 ( .A1(n2415), .A2(n2414), .ZN(n2356) );
  INV_X1 U3129 ( .A(n2929), .ZN(n2927) );
  INV_X1 U3130 ( .A(n2995), .ZN(n1841) );
  OAI22_X4 U3132 ( .A1(n4102), .A2(n3705), .B1(n4089), .B2(n3703), .ZN(n3706)
         );
  INV_X4 U3133 ( .A(n3157), .ZN(n3158) );
  NAND2_X4 U3134 ( .A1(n3236), .A2(n3237), .ZN(n1844) );
  INV_X2 U3135 ( .A(n3238), .ZN(n3236) );
  INV_X4 U3136 ( .A(n3177), .ZN(n1991) );
  NAND2_X4 U3137 ( .A1(n2656), .A2(n2657), .ZN(n2732) );
  NAND2_X1 U3138 ( .A1(n2851), .A2(n2850), .ZN(n2730) );
  NAND2_X1 U3139 ( .A1(n3193), .A2(n3142), .ZN(n3035) );
  NAND2_X4 U3140 ( .A1(n2554), .A2(n2553), .ZN(n2557) );
  XNOR2_X2 U3142 ( .A(n1847), .B(n1892), .ZN(n1846) );
  AND2_X4 U3143 ( .A1(net255581), .A2(n2424), .ZN(n2430) );
  NAND2_X1 U3144 ( .A1(n3271), .A2(n3173), .ZN(n1849) );
  NAND2_X4 U3145 ( .A1(n2926), .A2(n2925), .ZN(n3105) );
  XNOR2_X2 U3146 ( .A(n2922), .B(n2921), .ZN(n1950) );
  INV_X1 U3147 ( .A(n3102), .ZN(n1885) );
  NAND2_X2 U3148 ( .A1(n2560), .A2(n1891), .ZN(n2653) );
  INV_X1 U3149 ( .A(n2899), .ZN(n1853) );
  INV_X8 U3150 ( .A(n2821), .ZN(n2899) );
  INV_X1 U3151 ( .A(n2855), .ZN(n1854) );
  NAND2_X4 U3152 ( .A1(n2801), .A2(n2859), .ZN(n2854) );
  NAND3_X2 U3153 ( .A1(n3129), .A2(a[19]), .A3(n1460), .ZN(n3297) );
  INV_X2 U3154 ( .A(n2425), .ZN(n1990) );
  NAND2_X4 U3155 ( .A1(n3426), .A2(n3569), .ZN(n3570) );
  NAND3_X2 U3156 ( .A1(a[13]), .A2(n2701), .A3(net256143), .ZN(n2771) );
  AOI21_X2 U3157 ( .B1(n2333), .B2(n2334), .A(n1414), .ZN(n1857) );
  NAND2_X4 U3158 ( .A1(n1770), .A2(net255714), .ZN(n1858) );
  OAI21_X2 U3159 ( .B1(net253816), .B2(net253815), .A(n3610), .ZN(n1920) );
  NAND3_X2 U3160 ( .A1(a[15]), .A2(n2819), .A3(n1460), .ZN(n2900) );
  NAND3_X2 U3161 ( .A1(n3421), .A2(a[23]), .A3(net256143), .ZN(n3574) );
  NAND2_X1 U3162 ( .A1(a[24]), .A2(net256143), .ZN(n3571) );
  NAND3_X2 U3163 ( .A1(n2970), .A2(a[17]), .A3(n1460), .ZN(n3045) );
  NAND3_X2 U3164 ( .A1(a[21]), .A2(n3295), .A3(n1460), .ZN(n3359) );
  NAND3_X2 U3165 ( .A1(n3656), .A2(a[25]), .A3(net256143), .ZN(n3723) );
  NAND2_X4 U3166 ( .A1(n3120), .A2(n3121), .ZN(n3209) );
  NAND2_X4 U3167 ( .A1(n3038), .A2(n3039), .ZN(n3120) );
  NAND3_X1 U3168 ( .A1(n2044), .A2(n2045), .A3(n2058), .ZN(n2047) );
  NAND2_X1 U3169 ( .A1(n2148), .A2(n2182), .ZN(n2144) );
  INV_X1 U3170 ( .A(n2157), .ZN(n1863) );
  NAND2_X4 U3171 ( .A1(net254567), .A2(n3029), .ZN(n3030) );
  XNOR2_X2 U3172 ( .A(n2223), .B(n2226), .ZN(n1864) );
  NAND2_X4 U3173 ( .A1(net256032), .A2(net256033), .ZN(n1865) );
  NAND2_X4 U3174 ( .A1(n2816), .A2(net254669), .ZN(net254872) );
  NAND2_X2 U3175 ( .A1(n3678), .A2(n1937), .ZN(n3556) );
  INV_X4 U3176 ( .A(net257295), .ZN(net257296) );
  NOR2_X4 U3177 ( .A1(n3565), .A2(n3566), .ZN(n3589) );
  NAND2_X4 U3178 ( .A1(n2685), .A2(n1929), .ZN(n2709) );
  INV_X4 U3179 ( .A(n1459), .ZN(net256527) );
  INV_X1 U3180 ( .A(n3406), .ZN(n3407) );
  OAI21_X2 U3181 ( .B1(n3406), .B2(net256184), .A(n2804), .ZN(n2864) );
  NOR2_X2 U3182 ( .A1(n3681), .A2(n3682), .ZN(n3607) );
  NAND2_X4 U3183 ( .A1(n2402), .A2(n2401), .ZN(n2553) );
  NAND2_X1 U3184 ( .A1(n2347), .A2(n2348), .ZN(n2300) );
  NOR2_X4 U3185 ( .A1(n2627), .A2(n2626), .ZN(n2540) );
  INV_X4 U3186 ( .A(n3604), .ZN(n1877) );
  XNOR2_X2 U3187 ( .A(n2154), .B(n1412), .ZN(n1868) );
  AND2_X2 U3188 ( .A1(net255092), .A2(n2466), .ZN(n2574) );
  NAND2_X1 U3189 ( .A1(a[8]), .A2(net256135), .ZN(n2578) );
  INV_X2 U3190 ( .A(n2578), .ZN(n2466) );
  NAND2_X4 U3191 ( .A1(n1869), .A2(n3843), .ZN(n3942) );
  XNOR2_X2 U3192 ( .A(n3842), .B(n3870), .ZN(n1869) );
  NAND2_X4 U3193 ( .A1(n3867), .A2(n3868), .ZN(n3842) );
  NAND2_X4 U3194 ( .A1(n3899), .A2(n3939), .ZN(n3800) );
  NAND2_X4 U3195 ( .A1(n2054), .A2(n2053), .ZN(n2183) );
  OAI21_X2 U3196 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n4010) );
  NAND2_X4 U3197 ( .A1(n2061), .A2(n1808), .ZN(n2065) );
  BUF_X4 U3198 ( .A(n3809), .Z(n1870) );
  OAI221_X1 U3199 ( .B1(net253308), .B2(n3762), .C1(n3761), .C2(net256184), 
        .A(n3760), .ZN(net253570) );
  INV_X1 U3200 ( .A(n4012), .ZN(n4013) );
  INV_X1 U3201 ( .A(n4011), .ZN(n4018) );
  NOR3_X2 U3202 ( .A1(n4014), .A2(n4018), .A3(n4013), .ZN(n4058) );
  NOR3_X2 U3203 ( .A1(n4100), .A2(net255790), .A3(net255878), .ZN(n2068) );
  AOI21_X4 U3204 ( .B1(n3902), .B2(n3940), .A(n3901), .ZN(n3903) );
  NOR2_X2 U3205 ( .A1(net254059), .A2(net254058), .ZN(n3413) );
  NAND2_X1 U3207 ( .A1(n2612), .A2(n2578), .ZN(n2748) );
  NAND2_X4 U3208 ( .A1(n3802), .A2(n3801), .ZN(n3862) );
  NAND2_X4 U3209 ( .A1(n3479), .A2(n3478), .ZN(n3485) );
  XNOR2_X1 U3210 ( .A(n2514), .B(n2513), .ZN(n1874) );
  INV_X4 U3211 ( .A(n2324), .ZN(n1875) );
  NAND2_X2 U3212 ( .A1(n2467), .A2(net255380), .ZN(n1984) );
  NAND3_X2 U3213 ( .A1(n3244), .A2(net254296), .A3(n3455), .ZN(n3114) );
  NAND2_X4 U3214 ( .A1(n3350), .A2(n3351), .ZN(n3384) );
  XNOR2_X2 U3215 ( .A(n3387), .B(n1880), .ZN(n1879) );
  NOR2_X4 U3216 ( .A1(n1859), .A2(n1909), .ZN(n1881) );
  NAND2_X4 U3217 ( .A1(n3567), .A2(n3568), .ZN(n3558) );
  XNOR2_X2 U3218 ( .A(n3861), .B(n1972), .ZN(product_out[28]) );
  NAND2_X4 U3219 ( .A1(net253820), .A2(net257171), .ZN(net254086) );
  OAI21_X2 U3220 ( .B1(net253182), .B2(net253535), .A(n3789), .ZN(n3791) );
  INV_X1 U3221 ( .A(net253209), .ZN(net257044) );
  XNOR2_X2 U3222 ( .A(n1884), .B(net253191), .ZN(n1973) );
  AND3_X4 U3223 ( .A1(net257661), .A2(net253198), .A3(net253192), .ZN(n1884)
         );
  NOR2_X2 U3224 ( .A1(n3546), .A2(n1754), .ZN(n3555) );
  OAI21_X2 U3225 ( .B1(n1921), .B2(n3796), .A(net253522), .ZN(n3798) );
  AOI21_X4 U3226 ( .B1(n3278), .B2(n3284), .A(n3285), .ZN(n3189) );
  XNOR2_X2 U3227 ( .A(n3842), .B(n3870), .ZN(n1887) );
  INV_X4 U3228 ( .A(n1887), .ZN(n3844) );
  OAI21_X4 U3229 ( .B1(n3499), .B2(n3500), .A(n3498), .ZN(n3501) );
  NAND2_X2 U3230 ( .A1(n2319), .A2(n1829), .ZN(n2210) );
  NOR2_X2 U3231 ( .A1(n3801), .A2(n3800), .ZN(n3751) );
  INV_X1 U3232 ( .A(n4108), .ZN(n1888) );
  INV_X2 U3233 ( .A(n1888), .ZN(n1889) );
  AND2_X2 U3234 ( .A1(net253533), .A2(n3790), .ZN(net257159) );
  XNOR2_X2 U3235 ( .A(n2573), .B(n2473), .ZN(n1891) );
  OAI21_X2 U3236 ( .B1(n3977), .B2(n3997), .A(n3996), .ZN(n4071) );
  NAND2_X4 U3237 ( .A1(n3244), .A2(net254296), .ZN(n3323) );
  NAND2_X4 U3238 ( .A1(n3176), .A2(n2941), .ZN(n2875) );
  NAND2_X4 U3239 ( .A1(n4087), .A2(n3168), .ZN(n1892) );
  NAND2_X4 U3240 ( .A1(n1759), .A2(n3165), .ZN(n3168) );
  NAND2_X2 U3241 ( .A1(n3273), .A2(n3168), .ZN(n3530) );
  NAND2_X4 U3242 ( .A1(n2923), .A2(n2924), .ZN(n1895) );
  OAI21_X4 U3243 ( .B1(n2363), .B2(n2364), .A(n2362), .ZN(n1897) );
  OAI21_X4 U3244 ( .B1(n1932), .B2(n2493), .A(n2572), .ZN(n2473) );
  NAND2_X4 U3245 ( .A1(n2744), .A2(n2745), .ZN(n1898) );
  OAI21_X4 U3246 ( .B1(net255790), .B2(n2199), .A(net256402), .ZN(n2251) );
  NAND2_X4 U3247 ( .A1(n3795), .A2(net253584), .ZN(net253451) );
  NAND2_X2 U3248 ( .A1(n2683), .A2(n2682), .ZN(n2615) );
  XNOR2_X2 U3249 ( .A(net255284), .B(net255226), .ZN(n1902) );
  NAND2_X4 U3250 ( .A1(n1832), .A2(n3260), .ZN(n3492) );
  NAND2_X4 U3251 ( .A1(net255855), .A2(n1781), .ZN(net255533) );
  NOR2_X4 U3252 ( .A1(n1900), .A2(n1416), .ZN(n1899) );
  INV_X8 U3253 ( .A(n1899), .ZN(n3180) );
  XNOR2_X2 U3254 ( .A(n2919), .B(n2918), .ZN(n1900) );
  NAND2_X4 U3255 ( .A1(n3583), .A2(n3651), .ZN(n3646) );
  NAND2_X4 U3256 ( .A1(net256032), .A2(net256033), .ZN(net257127) );
  XNOR2_X1 U3257 ( .A(n3418), .B(n3423), .ZN(n1913) );
  INV_X8 U3258 ( .A(n3418), .ZN(n3576) );
  NAND2_X4 U3259 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  NAND2_X4 U3260 ( .A1(n3318), .A2(n3317), .ZN(n1903) );
  INV_X4 U3261 ( .A(n3316), .ZN(n3317) );
  NAND2_X2 U3262 ( .A1(n3318), .A2(n3317), .ZN(n3635) );
  XNOR2_X1 U3263 ( .A(n2643), .B(n1408), .ZN(n1907) );
  INV_X1 U3264 ( .A(n1872), .ZN(n2099) );
  XNOR2_X2 U3265 ( .A(n3329), .B(n3328), .ZN(n1905) );
  OAI22_X4 U3266 ( .A1(n2351), .A2(net256184), .B1(n3513), .B2(net256095), 
        .ZN(n2353) );
  BUF_X4 U3267 ( .A(n3442), .Z(n1908) );
  INV_X4 U3268 ( .A(n3287), .ZN(n3186) );
  OAI21_X4 U3269 ( .B1(n3609), .B2(n3608), .A(net253823), .ZN(n1909) );
  XNOR2_X2 U3270 ( .A(n2215), .B(n2278), .ZN(n1912) );
  INV_X2 U3271 ( .A(n3575), .ZN(n3423) );
  INV_X1 U3272 ( .A(n1941), .ZN(n3003) );
  NAND2_X4 U3273 ( .A1(net254633), .A2(net254634), .ZN(net254470) );
  INV_X2 U3274 ( .A(n3284), .ZN(n1914) );
  INV_X8 U3275 ( .A(n3174), .ZN(n3284) );
  INV_X4 U3276 ( .A(n2719), .ZN(n2717) );
  NAND2_X4 U3277 ( .A1(n1975), .A2(n1404), .ZN(net254004) );
  INV_X2 U3278 ( .A(n2290), .ZN(n2293) );
  NAND2_X1 U3279 ( .A1(n2290), .A2(n2291), .ZN(n2240) );
  INV_X8 U3280 ( .A(n3634), .ZN(n1915) );
  OAI21_X4 U3281 ( .B1(n2947), .B2(n2946), .A(n1261), .ZN(n1916) );
  BUF_X8 U3282 ( .A(n3975), .Z(n1917) );
  NAND2_X4 U3283 ( .A1(n3906), .A2(n1772), .ZN(n3975) );
  INV_X4 U3284 ( .A(n2941), .ZN(n3026) );
  NAND2_X4 U3285 ( .A1(n2070), .A2(n3955), .ZN(n2105) );
  NAND2_X2 U3286 ( .A1(n1598), .A2(n2871), .ZN(n2720) );
  XNOR2_X2 U3287 ( .A(net255047), .B(net256376), .ZN(net256795) );
  XNOR2_X1 U3288 ( .A(net256375), .B(n3628), .ZN(n3615) );
  INV_X2 U3289 ( .A(net255324), .ZN(net256303) );
  NAND2_X4 U3290 ( .A1(net255714), .A2(n2251), .ZN(n2201) );
  NAND2_X4 U3291 ( .A1(n2153), .A2(n1820), .ZN(n2155) );
  AND2_X4 U3292 ( .A1(control[0]), .A2(n1466), .ZN(n1922) );
  INV_X4 U3293 ( .A(n1922), .ZN(n3512) );
  INV_X4 U3294 ( .A(n1999), .ZN(n2072) );
  INV_X1 U3295 ( .A(n2088), .ZN(n1923) );
  INV_X4 U3296 ( .A(n3987), .ZN(n1924) );
  INV_X4 U3297 ( .A(n2497), .ZN(n1925) );
  NAND3_X4 U3298 ( .A1(n1317), .A2(n1544), .A3(n3349), .ZN(n3350) );
  CLKBUF_X3 U3299 ( .A(n3041), .Z(n1928) );
  NAND2_X4 U3300 ( .A1(n2607), .A2(n2606), .ZN(n1929) );
  NAND2_X4 U3301 ( .A1(n2607), .A2(n2606), .ZN(n2834) );
  INV_X8 U3302 ( .A(n2604), .ZN(n2607) );
  AND2_X2 U3303 ( .A1(n3993), .A2(net253156), .ZN(n1930) );
  INV_X2 U3304 ( .A(n1963), .ZN(n3641) );
  INV_X4 U3305 ( .A(n2494), .ZN(n2491) );
  NAND2_X4 U3306 ( .A1(net256077), .A2(a[3]), .ZN(n2037) );
  XNOR2_X2 U3307 ( .A(n2636), .B(n2635), .ZN(n1934) );
  XNOR2_X1 U3308 ( .A(n1907), .B(n2650), .ZN(product_out[13]) );
  NAND3_X2 U3309 ( .A1(n3390), .A2(n3389), .A3(net257407), .ZN(n3394) );
  NAND2_X4 U3310 ( .A1(n2494), .A2(n2493), .ZN(n2572) );
  INV_X2 U3311 ( .A(n2978), .ZN(n2976) );
  INV_X2 U3312 ( .A(net256290), .ZN(net255770) );
  NAND2_X2 U3313 ( .A1(n2207), .A2(net256290), .ZN(n2322) );
  BUF_X8 U3314 ( .A(n3352), .Z(n1936) );
  XNOR2_X2 U3315 ( .A(n3908), .B(n3907), .ZN(n1938) );
  NAND2_X4 U3316 ( .A1(n3937), .A2(n3975), .ZN(n3907) );
  AOI21_X2 U3317 ( .B1(n3024), .B2(n3023), .A(n1899), .ZN(n3028) );
  NAND2_X1 U3318 ( .A1(n1440), .A2(n3492), .ZN(n3270) );
  NAND2_X4 U3319 ( .A1(n3353), .A2(n1936), .ZN(n3235) );
  NAND4_X2 U3320 ( .A1(n2024), .A2(n2023), .A3(n2022), .A4(n2021), .ZN(n1940)
         );
  NAND4_X4 U3321 ( .A1(b[0]), .A2(control[1]), .A3(a[1]), .A4(control[0]), 
        .ZN(n2021) );
  NOR2_X4 U3322 ( .A1(n3071), .A2(n1405), .ZN(n1942) );
  NAND2_X4 U3323 ( .A1(n1390), .A2(net256119), .ZN(n2119) );
  XNOR2_X2 U3324 ( .A(n1535), .B(n2477), .ZN(n1945) );
  INV_X4 U3325 ( .A(n2467), .ZN(n1983) );
  NAND2_X2 U3326 ( .A1(n2579), .A2(net255091), .ZN(n2467) );
  XNOR2_X2 U3327 ( .A(n1774), .B(n3345), .ZN(n3346) );
  INV_X8 U3328 ( .A(n3146), .ZN(n3033) );
  NAND2_X4 U3330 ( .A1(net253449), .A2(net253450), .ZN(net253396) );
  INV_X1 U3331 ( .A(net253286), .ZN(net253296) );
  INV_X8 U3332 ( .A(n1822), .ZN(n2371) );
  INV_X8 U3333 ( .A(n2060), .ZN(n1952) );
  CLKBUF_X3 U3334 ( .A(net255409), .Z(net256909) );
  OAI21_X4 U3335 ( .B1(net255437), .B2(net255438), .A(net257560), .ZN(
        net256907) );
  OAI21_X4 U3336 ( .B1(n1948), .B2(net255232), .A(net255101), .ZN(net254949)
         );
  CLKBUF_X3 U3337 ( .A(n3042), .Z(n1955) );
  NAND2_X4 U3338 ( .A1(n3040), .A2(n2911), .ZN(n3042) );
  NAND4_X4 U3339 ( .A1(n1465), .A2(n1358), .A3(a[2]), .A4(b[25]), .ZN(n2062)
         );
  NOR2_X2 U3340 ( .A1(n1876), .A2(n3756), .ZN(net253591) );
  NAND4_X4 U3341 ( .A1(b[17]), .A2(control[0]), .A3(a[0]), .A4(net257782), 
        .ZN(n2014) );
  INV_X4 U3342 ( .A(n2790), .ZN(n1957) );
  NAND2_X2 U3343 ( .A1(n1995), .A2(n3026), .ZN(n3282) );
  OAI21_X4 U3344 ( .B1(n3990), .B2(net256927), .A(n3989), .ZN(net253198) );
  INV_X2 U3345 ( .A(net256907), .ZN(net255217) );
  NAND2_X4 U3346 ( .A1(n2120), .A2(n4100), .ZN(n2141) );
  XNOR2_X2 U3347 ( .A(n3860), .B(net253173), .ZN(n1958) );
  OAI211_X4 U3348 ( .C1(net256839), .C2(net253419), .A(n3859), .B(net253176), 
        .ZN(n3860) );
  NAND2_X4 U3349 ( .A1(n1959), .A2(n1405), .ZN(net254364) );
  XNOR2_X2 U3350 ( .A(n1810), .B(n3070), .ZN(n1959) );
  XNOR2_X2 U3351 ( .A(n1961), .B(n3204), .ZN(n1960) );
  XNOR2_X2 U3352 ( .A(n3065), .B(n3064), .ZN(n1962) );
  NAND2_X4 U3353 ( .A1(n3036), .A2(n3035), .ZN(n3065) );
  NAND2_X4 U3354 ( .A1(n3548), .A2(n3348), .ZN(net254192) );
  XNOR2_X1 U3355 ( .A(n3436), .B(n3558), .ZN(n1963) );
  XNOR2_X2 U3356 ( .A(n2103), .B(n2001), .ZN(net256843) );
  NAND2_X2 U3357 ( .A1(n2027), .A2(n1862), .ZN(n2043) );
  NAND2_X2 U3358 ( .A1(n2711), .A2(n1823), .ZN(net254770) );
  XNOR2_X2 U3359 ( .A(n3372), .B(n3432), .ZN(n1964) );
  XNOR2_X2 U3360 ( .A(n2980), .B(n1966), .ZN(n1965) );
  INV_X4 U3361 ( .A(n1767), .ZN(n2983) );
  AND2_X2 U3362 ( .A1(n3193), .A2(n1202), .ZN(n1966) );
  NAND2_X1 U3363 ( .A1(n2577), .A2(n2576), .ZN(n2580) );
  NAND4_X2 U3364 ( .A1(n2677), .A2(n2755), .A3(net254992), .A4(n2676), .ZN(
        net255046) );
  XNOR2_X2 U3366 ( .A(n2012), .B(n2011), .ZN(n1967) );
  XNOR2_X2 U3367 ( .A(n2154), .B(n1412), .ZN(n2123) );
  XNOR2_X2 U3368 ( .A(n1124), .B(n3911), .ZN(n1969) );
  XNOR2_X2 U3369 ( .A(n2589), .B(n1423), .ZN(n1970) );
  INV_X2 U3370 ( .A(n2589), .ZN(n2691) );
  INV_X2 U3371 ( .A(n1436), .ZN(n1971) );
  NAND2_X2 U3372 ( .A1(net257702), .A2(n2497), .ZN(n2397) );
  NAND3_X2 U3373 ( .A1(net257702), .A2(n2496), .A3(n2495), .ZN(n2422) );
  NAND3_X2 U3374 ( .A1(n2496), .A2(net255341), .A3(n2495), .ZN(n2498) );
  NAND3_X2 U3375 ( .A1(n2129), .A2(n2265), .A3(n2264), .ZN(n2268) );
  INV_X2 U3376 ( .A(n2129), .ZN(n2126) );
  XNOR2_X2 U3377 ( .A(n2529), .B(n1420), .ZN(n1974) );
  OAI22_X4 U3378 ( .A1(n1162), .A2(n3018), .B1(n3017), .B2(n3016), .ZN(n3019)
         );
  XNOR2_X2 U3379 ( .A(n3241), .B(n3240), .ZN(n1975) );
  NAND2_X4 U3380 ( .A1(n3533), .A2(n3532), .ZN(n3535) );
  OAI21_X4 U3381 ( .B1(n1838), .B2(n2756), .A(n2755), .ZN(net255045) );
  INV_X2 U3382 ( .A(n3624), .ZN(n1977) );
  XNOR2_X2 U3383 ( .A(n1801), .B(n3150), .ZN(n1978) );
  XNOR2_X2 U3384 ( .A(n1868), .B(n1998), .ZN(n1979) );
  NAND2_X4 U3385 ( .A1(n2612), .A2(n1392), .ZN(n2681) );
  NAND3_X4 U3386 ( .A1(control[0]), .A2(a[3]), .A3(b[0]), .ZN(n1980) );
  NAND2_X1 U3387 ( .A1(net257069), .A2(net254057), .ZN(n3629) );
  XNOR2_X2 U3388 ( .A(n2376), .B(n2435), .ZN(n1982) );
  OAI21_X4 U3389 ( .B1(n3195), .B2(n3194), .A(n3198), .ZN(n3202) );
  AOI21_X4 U3390 ( .B1(n3014), .B2(n3013), .A(n2005), .ZN(n3017) );
  NAND2_X2 U3391 ( .A1(n2621), .A2(n2620), .ZN(n1988) );
  NAND2_X2 U3392 ( .A1(net255098), .A2(n1118), .ZN(net255097) );
  NAND2_X1 U3393 ( .A1(n3455), .A2(n3247), .ZN(n3115) );
  INV_X8 U3394 ( .A(n3247), .ZN(n3324) );
  INV_X4 U3395 ( .A(n3068), .ZN(n3066) );
  INV_X1 U3396 ( .A(n1451), .ZN(net256741) );
  NAND2_X4 U3397 ( .A1(net256742), .A2(n1983), .ZN(n1985) );
  NAND2_X4 U3398 ( .A1(n1984), .A2(n1985), .ZN(net255378) );
  NAND2_X2 U3399 ( .A1(n2505), .A2(net257485), .ZN(net255587) );
  OAI21_X4 U3400 ( .B1(net255776), .B2(net255777), .A(net255775), .ZN(n2206)
         );
  AND2_X4 U3401 ( .A1(n1786), .A2(net254770), .ZN(net256376) );
  INV_X4 U3402 ( .A(n3086), .ZN(n3761) );
  NAND2_X1 U3403 ( .A1(n1929), .A2(n2833), .ZN(n2835) );
  NAND2_X4 U3404 ( .A1(n3605), .A2(n1878), .ZN(n3606) );
  NOR2_X2 U3405 ( .A1(n1411), .A2(n2371), .ZN(n2200) );
  INV_X4 U3406 ( .A(n3140), .ZN(n2915) );
  NAND2_X4 U3407 ( .A1(n3596), .A2(n3556), .ZN(n3594) );
  NAND2_X1 U3408 ( .A1(n2436), .A2(n1137), .ZN(n2437) );
  NAND2_X2 U3409 ( .A1(a[10]), .A2(n1999), .ZN(n2382) );
  NAND3_X2 U3410 ( .A1(n3140), .A2(n3139), .A3(n2962), .ZN(n2963) );
  NAND2_X2 U3411 ( .A1(a[8]), .A2(n1232), .ZN(n2325) );
  INV_X1 U3412 ( .A(net253797), .ZN(net253913) );
  NAND4_X4 U3413 ( .A1(b[1]), .A2(control[1]), .A3(a[0]), .A4(control[0]), 
        .ZN(n2013) );
  NAND2_X4 U3414 ( .A1(n3066), .A2(n3067), .ZN(n3113) );
  AOI21_X4 U3415 ( .B1(n1291), .B2(n3455), .A(net254302), .ZN(n3245) );
  NAND2_X4 U3416 ( .A1(n2785), .A2(n2784), .ZN(net254669) );
  NOR2_X4 U3417 ( .A1(net256874), .A2(net254948), .ZN(net254940) );
  AOI21_X1 U3418 ( .B1(n1783), .B2(net257650), .A(n3994), .ZN(n3997) );
  NAND3_X4 U3419 ( .A1(n3089), .A2(product_in[19]), .A3(net256095), .ZN(n3336)
         );
  NOR2_X1 U3420 ( .A1(net256145), .A2(n4028), .ZN(n4031) );
  NAND2_X1 U3421 ( .A1(n2892), .A2(n2885), .ZN(n2780) );
  NAND3_X2 U3422 ( .A1(n2889), .A2(n2885), .A3(n2835), .ZN(n2893) );
  INV_X2 U3423 ( .A(n2778), .ZN(n2777) );
  NAND2_X4 U3424 ( .A1(n2779), .A2(n2778), .ZN(n2885) );
  NOR2_X1 U3425 ( .A1(net256145), .A2(net254656), .ZN(n2969) );
  OAI21_X1 U3426 ( .B1(net255721), .B2(n2839), .A(n2702), .ZN(n2703) );
  NAND3_X2 U3427 ( .A1(a[1]), .A2(n2168), .A3(net256105), .ZN(n2306) );
  INV_X1 U3428 ( .A(n2168), .ZN(n2167) );
  NOR2_X2 U3429 ( .A1(n3143), .A2(n2915), .ZN(net254766) );
  INV_X1 U3430 ( .A(n3192), .ZN(n3062) );
  NOR2_X2 U3431 ( .A1(n3063), .A2(n3192), .ZN(n3195) );
  NOR2_X1 U3432 ( .A1(net256095), .A2(n1895), .ZN(n2998) );
  NAND2_X1 U3433 ( .A1(net256099), .A2(n1895), .ZN(n2993) );
  NAND2_X4 U3434 ( .A1(n2656), .A2(n2734), .ZN(n2640) );
  XNOR2_X1 U3435 ( .A(n2646), .B(n2565), .ZN(product_out[12]) );
  NAND3_X2 U3436 ( .A1(net255543), .A2(net257240), .A3(n2367), .ZN(n2368) );
  NAND2_X4 U3437 ( .A1(n1986), .A2(n1987), .ZN(n1989) );
  NAND2_X4 U3438 ( .A1(n1988), .A2(n1989), .ZN(net255166) );
  INV_X4 U3439 ( .A(n2621), .ZN(n1986) );
  INV_X4 U3440 ( .A(n2620), .ZN(n1987) );
  NAND2_X4 U3441 ( .A1(n2658), .A2(n2734), .ZN(n3010) );
  INV_X8 U3442 ( .A(n2533), .ZN(n2627) );
  NAND3_X2 U3443 ( .A1(n2365), .A2(n1990), .A3(net255459), .ZN(n2366) );
  NAND2_X1 U3444 ( .A1(n2859), .A2(n2860), .ZN(n2858) );
  NAND2_X4 U3445 ( .A1(n2336), .A2(n2337), .ZN(n2362) );
  NAND2_X4 U3446 ( .A1(n2944), .A2(n2945), .ZN(n2946) );
  NAND2_X4 U3447 ( .A1(n3559), .A2(n3560), .ZN(n3640) );
  NAND2_X4 U3448 ( .A1(n2608), .A2(n2834), .ZN(n2759) );
  OAI211_X4 U3449 ( .C1(n1129), .C2(net256095), .A(n2798), .B(n2797), .ZN(
        n2801) );
  INV_X8 U3450 ( .A(n2944), .ZN(n2668) );
  OAI21_X4 U3451 ( .B1(net255102), .B2(net256303), .A(net255104), .ZN(
        net255096) );
  NAND2_X4 U3452 ( .A1(n2469), .A2(n2470), .ZN(n2630) );
  NAND2_X4 U3453 ( .A1(net255454), .A2(net255453), .ZN(net255459) );
  NAND2_X4 U3454 ( .A1(n2163), .A2(n2162), .ZN(n2315) );
  NAND2_X4 U3455 ( .A1(n2413), .A2(n2481), .ZN(n2482) );
  OAI211_X4 U3456 ( .C1(n2995), .C2(net256095), .A(n2409), .B(n2410), .ZN(
        n2413) );
  NAND2_X4 U3457 ( .A1(n1247), .A2(n2742), .ZN(n2746) );
  NOR2_X2 U3458 ( .A1(n2574), .A2(net255223), .ZN(n2575) );
  NAND2_X4 U3459 ( .A1(n2426), .A2(n2314), .ZN(n2215) );
  NAND2_X2 U3460 ( .A1(a[7]), .A2(net257127), .ZN(n2436) );
  INV_X8 U3461 ( .A(n2537), .ZN(n2628) );
  XNOR2_X2 U3462 ( .A(n2848), .B(n1994), .ZN(n3405) );
  NAND3_X4 U3463 ( .A1(n2446), .A2(n2445), .A3(n2444), .ZN(n2700) );
  NAND2_X4 U3464 ( .A1(net255915), .A2(net255779), .ZN(n2446) );
  NAND2_X2 U3465 ( .A1(n3456), .A2(n3457), .ZN(n3461) );
  NAND2_X4 U3466 ( .A1(n2422), .A2(n1926), .ZN(n2573) );
  NAND2_X1 U3467 ( .A1(a[0]), .A2(n1460), .ZN(n2010) );
  NAND3_X1 U3468 ( .A1(a[27]), .A2(n3823), .A3(net256143), .ZN(n3874) );
  NAND2_X1 U3469 ( .A1(a[27]), .A2(net256143), .ZN(n3821) );
  NAND2_X1 U3470 ( .A1(a[26]), .A2(net256143), .ZN(n3726) );
  NAND3_X1 U3471 ( .A1(n2695), .A2(n2686), .A3(n2687), .ZN(n2602) );
  NOR2_X1 U3472 ( .A1(n2696), .A2(n2695), .ZN(n2600) );
  NAND3_X2 U3473 ( .A1(a[11]), .A2(net256141), .A3(n2591), .ZN(n2686) );
  NAND2_X2 U3474 ( .A1(a[1]), .A2(net256388), .ZN(n2011) );
  NAND2_X2 U3475 ( .A1(n2534), .A2(n2536), .ZN(n2395) );
  AOI211_X2 U3476 ( .C1(n2598), .C2(n2688), .A(n1794), .B(n2588), .ZN(n2603)
         );
  NOR2_X4 U3477 ( .A1(n2831), .A2(n2887), .ZN(n2832) );
  NAND2_X4 U3478 ( .A1(n2431), .A2(n2505), .ZN(n2432) );
  XNOR2_X1 U3479 ( .A(n2486), .B(n1126), .ZN(product_out[11]) );
  XNOR2_X1 U3480 ( .A(n2482), .B(n4109), .ZN(product_out[10]) );
  NAND2_X4 U3481 ( .A1(n2355), .A2(n2354), .ZN(n2414) );
  INV_X2 U3482 ( .A(n2223), .ZN(n2225) );
  NAND2_X4 U3483 ( .A1(n3179), .A2(n3175), .ZN(n2792) );
  NAND2_X2 U3484 ( .A1(n2952), .A2(n2881), .ZN(n2815) );
  XNOR2_X2 U3485 ( .A(n2867), .B(n2875), .ZN(n2868) );
  NOR2_X2 U3486 ( .A1(net254683), .A2(net254681), .ZN(n2956) );
  NAND2_X2 U3487 ( .A1(n3026), .A2(n4093), .ZN(n2942) );
  INV_X2 U3488 ( .A(net256555), .ZN(net256556) );
  NOR2_X4 U3489 ( .A1(n1969), .A2(net253280), .ZN(n1993) );
  NAND2_X1 U3490 ( .A1(a[22]), .A2(net256165), .ZN(net253280) );
  NAND2_X4 U3491 ( .A1(n1927), .A2(n2468), .ZN(n2533) );
  INV_X2 U3492 ( .A(net255409), .ZN(net255413) );
  INV_X1 U3493 ( .A(net253824), .ZN(net256541) );
  OAI211_X4 U3494 ( .C1(n2256), .C2(n2255), .A(n2254), .B(n2253), .ZN(
        net255708) );
  NAND2_X4 U3495 ( .A1(n3069), .A2(n1962), .ZN(n3455) );
  NAND2_X4 U3496 ( .A1(n3467), .A2(n3468), .ZN(n3702) );
  NAND2_X4 U3497 ( .A1(n3808), .A2(n3807), .ZN(n3799) );
  OAI21_X4 U3498 ( .B1(n3685), .B2(n3686), .A(n3601), .ZN(net253390) );
  INV_X4 U3499 ( .A(n2000), .ZN(n1997) );
  NAND2_X4 U3500 ( .A1(n2180), .A2(n2150), .ZN(n2187) );
  INV_X1 U3501 ( .A(n1782), .ZN(n3544) );
  NAND3_X1 U3502 ( .A1(net253270), .A2(n3934), .A3(n3935), .ZN(n3936) );
  NAND2_X4 U3503 ( .A1(n3955), .A2(a[9]), .ZN(n2435) );
  INV_X4 U3504 ( .A(n3530), .ZN(n3173) );
  INV_X4 U3505 ( .A(n3181), .ZN(n2874) );
  NAND2_X4 U3506 ( .A1(net255611), .A2(a[5]), .ZN(n2103) );
  INV_X2 U3507 ( .A(n2700), .ZN(n2451) );
  NAND2_X4 U3508 ( .A1(n2287), .A2(n2286), .ZN(n2421) );
  NAND2_X4 U3509 ( .A1(n2553), .A2(n2554), .ZN(n2476) );
  INV_X1 U3510 ( .A(n3405), .ZN(n3409) );
  NAND2_X4 U3511 ( .A1(net255045), .A2(net255046), .ZN(net255047) );
  NAND2_X4 U3512 ( .A1(n3139), .A2(n3200), .ZN(n3145) );
  NAND3_X2 U3513 ( .A1(n2943), .A2(n3180), .A3(n2942), .ZN(n2988) );
  NAND3_X2 U3514 ( .A1(n3023), .A2(n1991), .A3(n3024), .ZN(n2943) );
  OAI211_X4 U3515 ( .C1(n2311), .C2(n2312), .A(n2310), .B(n2309), .ZN(n2361)
         );
  NAND2_X4 U3516 ( .A1(n1188), .A2(n2276), .ZN(n2309) );
  INV_X2 U3517 ( .A(net255459), .ZN(net255456) );
  NOR3_X4 U3518 ( .A1(n2697), .A2(n2696), .A3(n2695), .ZN(n2698) );
  AND4_X4 U3519 ( .A1(n2102), .A2(net255929), .A3(n2101), .A4(n2100), .ZN(
        n2001) );
  NAND2_X4 U3520 ( .A1(n3022), .A2(n1861), .ZN(n3085) );
  OAI21_X4 U3521 ( .B1(n2939), .B2(n2940), .A(n3179), .ZN(n3023) );
  NAND2_X4 U3522 ( .A1(n3200), .A2(n3143), .ZN(n3144) );
  INV_X8 U3523 ( .A(n3142), .ZN(n3200) );
  NAND4_X4 U3524 ( .A1(n1465), .A2(control[0]), .A3(a[2]), .A4(b[17]), .ZN(
        n2063) );
  NAND2_X4 U3525 ( .A1(n3211), .A2(n3210), .ZN(n3212) );
  NAND3_X2 U3526 ( .A1(n3549), .A2(n3604), .A3(n3548), .ZN(n3554) );
  NAND2_X4 U3528 ( .A1(net255378), .A2(net255379), .ZN(net255229) );
  NAND2_X4 U3529 ( .A1(n2576), .A2(n2577), .ZN(n2675) );
  AOI21_X4 U3530 ( .B1(n3697), .B2(net256097), .A(n3696), .ZN(net253564) );
  NAND2_X4 U3531 ( .A1(n3914), .A2(n3910), .ZN(n3996) );
  NAND2_X4 U3532 ( .A1(n2688), .A2(n2384), .ZN(n2516) );
  NAND2_X1 U3533 ( .A1(n2383), .A2(n2382), .ZN(n2384) );
  NAND2_X4 U3534 ( .A1(n2976), .A2(n2977), .ZN(n3193) );
  NAND2_X4 U3535 ( .A1(n3289), .A2(n3291), .ZN(n3241) );
  NAND2_X4 U3536 ( .A1(n2718), .A2(n2717), .ZN(n2741) );
  AOI22_X4 U3537 ( .A1(n3986), .A2(n3332), .B1(n3332), .B2(net256095), .ZN(
        n3334) );
  NOR2_X4 U3538 ( .A1(n3758), .A2(net253522), .ZN(net253701) );
  NAND2_X4 U3539 ( .A1(n3076), .A2(n3077), .ZN(n3184) );
  NAND2_X4 U3540 ( .A1(net254857), .A2(net254858), .ZN(net254696) );
  NAND2_X4 U3541 ( .A1(n2376), .A2(n2375), .ZN(n2443) );
  OAI22_X4 U3542 ( .A1(n2032), .A2(n2033), .B1(net256018), .B2(n2031), .ZN(
        n2092) );
  NAND2_X4 U3543 ( .A1(n2271), .A2(n2270), .ZN(n2313) );
  NAND2_X4 U3544 ( .A1(n1766), .A2(n3105), .ZN(n3020) );
  NAND2_X4 U3545 ( .A1(n2088), .A2(n2089), .ZN(n2164) );
  NAND2_X1 U3546 ( .A1(n1922), .A2(n3915), .ZN(n3916) );
  NAND2_X1 U3547 ( .A1(net256183), .A2(n3915), .ZN(n3259) );
  NAND2_X4 U3548 ( .A1(n4096), .A2(n2118), .ZN(n2191) );
  NAND3_X1 U3549 ( .A1(n2588), .A2(n2688), .A3(n2455), .ZN(n2456) );
  NAND2_X4 U3550 ( .A1(n2853), .A2(n2852), .ZN(n2856) );
  OAI21_X1 U3551 ( .B1(n2731), .B2(n2853), .A(n2852), .ZN(n2802) );
  XNOR2_X1 U3552 ( .A(n2730), .B(n2853), .ZN(product_out[14]) );
  NAND2_X4 U3553 ( .A1(n2729), .A2(n2852), .ZN(n2853) );
  NAND2_X1 U3554 ( .A1(n3343), .A2(n1779), .ZN(n3256) );
  NAND3_X4 U3555 ( .A1(a[16]), .A2(n2972), .A3(net256117), .ZN(n3116) );
  NAND2_X2 U3556 ( .A1(n2825), .A2(n2826), .ZN(n3041) );
  NAND3_X4 U3557 ( .A1(n1802), .A2(n2104), .A3(n1954), .ZN(net255910) );
  NAND2_X1 U3558 ( .A1(n1780), .A2(n2016), .ZN(n2018) );
  INV_X2 U3559 ( .A(net255225), .ZN(net255383) );
  NAND2_X4 U3560 ( .A1(n2983), .A2(n2982), .ZN(net254467) );
  NAND2_X4 U3561 ( .A1(n1997), .A2(n2108), .ZN(net255874) );
  NAND2_X2 U3562 ( .A1(n2316), .A2(n1324), .ZN(n2263) );
  NAND2_X4 U3563 ( .A1(n3438), .A2(n3290), .ZN(n3240) );
  NAND2_X4 U3564 ( .A1(net256032), .A2(net256033), .ZN(net256420) );
  NAND2_X4 U3565 ( .A1(n1999), .A2(n2067), .ZN(n2104) );
  OAI22_X2 U3566 ( .A1(n3564), .A2(n1915), .B1(n3564), .B2(n1963), .ZN(n3565)
         );
  NAND2_X4 U3567 ( .A1(n2419), .A2(n2421), .ZN(n2404) );
  NAND2_X4 U3568 ( .A1(n2305), .A2(n2304), .ZN(n2419) );
  NAND2_X4 U3569 ( .A1(n2020), .A2(a[1]), .ZN(n2071) );
  NAND4_X4 U3570 ( .A1(n2015), .A2(n2014), .A3(n2013), .A4(net256050), .ZN(
        n2020) );
  NOR2_X2 U3571 ( .A1(net256362), .A2(net253819), .ZN(n3610) );
  OAI211_X4 U3572 ( .C1(n2594), .C2(n2593), .A(n2592), .B(n2687), .ZN(n2690)
         );
  NAND2_X4 U3573 ( .A1(net254682), .A2(net254683), .ZN(net254688) );
  NAND3_X2 U3574 ( .A1(n3711), .A2(n3712), .A3(n3713), .ZN(n3808) );
  NAND3_X2 U3575 ( .A1(n3711), .A2(n3712), .A3(n3713), .ZN(n3683) );
  NAND2_X4 U3576 ( .A1(n3713), .A2(n3680), .ZN(n3597) );
  NAND2_X4 U3577 ( .A1(n3591), .A2(n3590), .ZN(n3713) );
  AOI21_X2 U3578 ( .B1(n1903), .B2(n3636), .A(n3634), .ZN(n3644) );
  OAI22_X4 U3579 ( .A1(n2430), .A2(n2429), .B1(n2427), .B2(n4103), .ZN(
        net255328) );
  NAND2_X4 U3580 ( .A1(n2978), .A2(n2979), .ZN(n3141) );
  NAND2_X4 U3581 ( .A1(n2057), .A2(n2058), .ZN(n2190) );
  INV_X4 U3582 ( .A(n1951), .ZN(n2281) );
  OAI21_X2 U3583 ( .B1(n2956), .B2(n2955), .A(net257979), .ZN(n2957) );
  OAI21_X1 U3584 ( .B1(n2732), .B2(n2658), .A(n2734), .ZN(n2724) );
  NAND3_X1 U3585 ( .A1(n1857), .A2(n1873), .A3(n2613), .ZN(n2508) );
  NAND2_X4 U3586 ( .A1(n2387), .A2(n2388), .ZN(n2609) );
  OAI22_X4 U3587 ( .A1(n2038), .A2(n2039), .B1(n2037), .B2(n2036), .ZN(n2094)
         );
  NAND3_X1 U3588 ( .A1(n2308), .A2(n2307), .A3(n2306), .ZN(n2282) );
  NAND2_X1 U3589 ( .A1(n2445), .A2(net256909), .ZN(n2329) );
  NAND2_X1 U3590 ( .A1(n2445), .A2(net256909), .ZN(n2327) );
  INV_X8 U3591 ( .A(n2445), .ZN(n2377) );
  NAND3_X4 U3592 ( .A1(n1792), .A2(net257586), .A3(n2249), .ZN(n2445) );
  NAND2_X4 U3593 ( .A1(net256032), .A2(net256033), .ZN(n1999) );
  INV_X16 U3594 ( .A(net256157), .ZN(net256153) );
  INV_X8 U3595 ( .A(n3640), .ZN(n3564) );
  XNOR2_X1 U3596 ( .A(n2933), .B(n3098), .ZN(product_out[17]) );
  NOR2_X4 U3597 ( .A1(n2989), .A2(n2990), .ZN(n2002) );
  NAND2_X1 U3598 ( .A1(a[11]), .A2(net256165), .ZN(n3107) );
  NOR3_X2 U3600 ( .A1(n3778), .A2(n3779), .A3(n3777), .ZN(product_out[27]) );
  NOR2_X2 U3601 ( .A1(n3773), .A2(n3772), .ZN(n3778) );
  NAND2_X4 U3602 ( .A1(n1182), .A2(n3315), .ZN(n3442) );
  NAND2_X4 U3603 ( .A1(n1817), .A2(n1937), .ZN(n3678) );
  NAND2_X4 U3604 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  NAND2_X4 U3605 ( .A1(n2877), .A2(n2876), .ZN(n2922) );
  NAND2_X4 U3606 ( .A1(n3019), .A2(n1766), .ZN(n3109) );
  NAND2_X4 U3607 ( .A1(net254004), .A2(n3453), .ZN(n3454) );
  NAND2_X4 U3608 ( .A1(n4095), .A2(n3327), .ZN(n3536) );
  NAND2_X4 U3609 ( .A1(n2732), .A2(n2734), .ZN(n3011) );
  NOR2_X4 U3610 ( .A1(n3386), .A2(n1410), .ZN(net256362) );
  NAND2_X4 U3611 ( .A1(n2525), .A2(n2682), .ZN(n2683) );
  NAND2_X4 U3612 ( .A1(n2523), .A2(n2524), .ZN(n2682) );
  NAND3_X2 U3613 ( .A1(n2535), .A2(n2536), .A3(n2629), .ZN(n2423) );
  NAND2_X4 U3614 ( .A1(n2795), .A2(n2796), .ZN(n3015) );
  NOR2_X4 U3615 ( .A1(n1886), .A2(n2796), .ZN(n2005) );
  NAND2_X4 U3616 ( .A1(n3805), .A2(n3806), .ZN(net253270) );
  NAND2_X4 U3617 ( .A1(n3935), .A2(net253270), .ZN(net253462) );
  AOI21_X4 U3618 ( .B1(n1195), .B2(n3856), .A(n1125), .ZN(n3858) );
  NAND2_X2 U3619 ( .A1(n3280), .A2(n1438), .ZN(n3187) );
  NAND2_X4 U3620 ( .A1(n2338), .A2(n2339), .ZN(n2535) );
  NAND2_X4 U3621 ( .A1(n2344), .A2(n2345), .ZN(n2420) );
  AOI22_X2 U3622 ( .A1(n2488), .A2(n1945), .B1(n2488), .B2(net256095), .ZN(
        n2479) );
  NAND2_X4 U3623 ( .A1(n3472), .A2(n3471), .ZN(n3856) );
  NAND2_X4 U3624 ( .A1(n3490), .A2(n3491), .ZN(net253182) );
  INV_X8 U3626 ( .A(n2878), .ZN(n2952) );
  NAND2_X4 U3627 ( .A1(n3710), .A2(net253643), .ZN(net253458) );
  INV_X8 U3629 ( .A(n3025), .ZN(n3177) );
  AOI22_X4 U3630 ( .A1(net254670), .A2(net257880), .B1(net254671), .B2(
        net254465), .ZN(net254635) );
  NAND3_X2 U3631 ( .A1(n1936), .A2(n3430), .A3(n3353), .ZN(n3312) );
  NAND2_X4 U3632 ( .A1(n3135), .A2(n3352), .ZN(n3204) );
  INV_X2 U3633 ( .A(n2590), .ZN(n2591) );
  INV_X4 U3634 ( .A(n2005), .ZN(n3012) );
  NOR2_X4 U3635 ( .A1(n3250), .A2(n1404), .ZN(n2006) );
  INV_X4 U3636 ( .A(n2006), .ZN(n3548) );
  NAND3_X2 U3637 ( .A1(net256306), .A2(net254562), .A3(net254761), .ZN(n2816)
         );
  NAND2_X4 U3638 ( .A1(n3113), .A2(net254467), .ZN(n3247) );
  NAND2_X4 U3639 ( .A1(n3031), .A2(n2960), .ZN(n3139) );
  NAND3_X2 U3640 ( .A1(n3437), .A2(n1844), .A3(n3442), .ZN(n3636) );
  INV_X8 U3642 ( .A(n2571), .ZN(n2737) );
  NAND2_X4 U3643 ( .A1(n2213), .A2(n2214), .ZN(n2314) );
  NAND2_X2 U3644 ( .A1(n2008), .A2(n2888), .ZN(n2685) );
  INV_X4 U3645 ( .A(n2007), .ZN(n2008) );
  INV_X8 U3646 ( .A(n2746), .ZN(n2949) );
  NOR2_X2 U3647 ( .A1(net253824), .A2(net253815), .ZN(n3414) );
  INV_X8 U3648 ( .A(net254052), .ZN(net253824) );
  INV_X4 U3649 ( .A(net256305), .ZN(net256306) );
  NAND2_X4 U3650 ( .A1(net255504), .A2(net255505), .ZN(net255092) );
  INV_X8 U3651 ( .A(n2193), .ZN(n2196) );
  NAND2_X4 U3652 ( .A1(n1168), .A2(n3412), .ZN(net253765) );
  NAND2_X4 U3653 ( .A1(n3439), .A2(n3440), .ZN(n3450) );
  OAI211_X4 U3654 ( .C1(n3444), .C2(n3451), .A(n3450), .B(n3449), .ZN(n3551)
         );
  NAND3_X2 U3655 ( .A1(n2247), .A2(n2246), .A3(net255724), .ZN(n2257) );
  NAND2_X4 U3656 ( .A1(n1864), .A2(n2224), .ZN(n2270) );
  NAND2_X4 U3657 ( .A1(n2633), .A2(n2634), .ZN(n2738) );
  XNOR2_X2 U3658 ( .A(n3456), .B(n3153), .ZN(net254414) );
  NAND2_X4 U3660 ( .A1(n2156), .A2(n1412), .ZN(n2185) );
  OAI22_X4 U3661 ( .A1(n1279), .A2(n2433), .B1(n2502), .B2(n2610), .ZN(n2465)
         );
  NAND2_X4 U3662 ( .A1(n2736), .A2(n3013), .ZN(n2846) );
  NAND2_X4 U3663 ( .A1(n3117), .A2(n3122), .ZN(n3206) );
  NAND2_X4 U3664 ( .A1(n3376), .A2(n3375), .ZN(n3637) );
  NAND2_X4 U3665 ( .A1(n1964), .A2(n3373), .ZN(n3563) );
  INV_X8 U3666 ( .A(n3709), .ZN(n3630) );
  NAND2_X4 U3667 ( .A1(n1935), .A2(n3395), .ZN(n3538) );
  NAND2_X4 U3668 ( .A1(n3698), .A2(net257630), .ZN(n3767) );
  OAI21_X2 U3669 ( .B1(n2672), .B2(n2671), .A(n1894), .ZN(n2716) );
  NAND2_X4 U3670 ( .A1(net253179), .A2(n3784), .ZN(n3698) );
  NAND2_X4 U3671 ( .A1(n1902), .A2(n2532), .ZN(n2944) );
  NAND2_X4 U3672 ( .A1(n2317), .A2(n2316), .ZN(n2427) );
  NAND3_X1 U3673 ( .A1(n3477), .A2(n1849), .A3(n1436), .ZN(n3478) );
  OAI211_X4 U3674 ( .C1(n3531), .C2(n1892), .A(n1436), .B(n3529), .ZN(n3542)
         );
  NAND2_X4 U3675 ( .A1(net256032), .A2(net256033), .ZN(n3955) );
  AOI21_X1 U3676 ( .B1(n3799), .B2(n1870), .A(n3806), .ZN(n3750) );
  NAND2_X4 U3677 ( .A1(n3799), .A2(n1870), .ZN(n3900) );
  NAND2_X4 U3678 ( .A1(n3041), .A2(n2829), .ZN(n3037) );
  NAND2_X4 U3679 ( .A1(n3188), .A2(n3189), .ZN(n3344) );
  NAND2_X4 U3680 ( .A1(n3091), .A2(n3092), .ZN(n3093) );
  NAND2_X4 U3681 ( .A1(n2938), .A2(n2806), .ZN(n2867) );
  AOI21_X4 U3682 ( .B1(n1134), .B2(n1914), .A(n3162), .ZN(n3163) );
  NAND3_X4 U3683 ( .A1(n2141), .A2(n1818), .A3(n1952), .ZN(n2193) );
  INV_X8 U3684 ( .A(n3613), .ZN(n3758) );
  NAND2_X4 U3686 ( .A1(n2512), .A2(n2592), .ZN(n2593) );
  OAI21_X4 U3687 ( .B1(n1479), .B2(n1753), .A(n3033), .ZN(n3197) );
  NAND2_X4 U3688 ( .A1(n2830), .A2(n1121), .ZN(n2889) );
  OAI211_X4 U3689 ( .C1(n2203), .C2(n2370), .A(n2371), .B(n2202), .ZN(n2323)
         );
  NAND2_X4 U3690 ( .A1(n2205), .A2(n2379), .ZN(net255726) );
  NAND2_X4 U3691 ( .A1(n2446), .A2(n2250), .ZN(n2379) );
  NAND2_X4 U3692 ( .A1(n2790), .A2(n2791), .ZN(n3179) );
  NAND2_X4 U3693 ( .A1(n2808), .A2(n2952), .ZN(n2789) );
  NAND2_X4 U3694 ( .A1(n3496), .A2(n3495), .ZN(n3499) );
  NAND2_X4 U3695 ( .A1(n2280), .A2(n1519), .ZN(n2307) );
  NAND2_X4 U3696 ( .A1(n2211), .A2(n2212), .ZN(n2426) );
  NAND2_X4 U3697 ( .A1(n2813), .A2(n2812), .ZN(n2950) );
  NAND2_X4 U3698 ( .A1(n3049), .A2(n3050), .ZN(n3217) );
  NAND3_X2 U3699 ( .A1(n3462), .A2(n3461), .A3(n3460), .ZN(n3603) );
  NAND2_X4 U3700 ( .A1(n3060), .A2(n3205), .ZN(n3208) );
  NAND2_X4 U3701 ( .A1(n3055), .A2(n3054), .ZN(n3056) );
  NAND2_X4 U3702 ( .A1(n3236), .A2(n3237), .ZN(n3438) );
  NAND2_X4 U3703 ( .A1(n3183), .A2(n3182), .ZN(n3280) );
  NAND3_X2 U3704 ( .A1(n1760), .A2(n1790), .A3(n3550), .ZN(n3463) );
  NAND2_X4 U3705 ( .A1(n3192), .A2(n3063), .ZN(n3198) );
  NOR2_X1 U3706 ( .A1(n1929), .A2(n2830), .ZN(n2761) );
  NAND2_X4 U3707 ( .A1(n1410), .A2(n3386), .ZN(net254052) );
  NAND2_X4 U3709 ( .A1(n2389), .A2(n2609), .ZN(n2506) );
  OAI211_X4 U3711 ( .C1(n2616), .C2(n1918), .A(n2615), .B(n2614), .ZN(n2617)
         );
  NAND3_X4 U3712 ( .A1(n2757), .A2(net255045), .A3(n1786), .ZN(net254761) );
  NAND3_X2 U3713 ( .A1(n1109), .A2(n3457), .A3(n3455), .ZN(n3462) );
  AOI21_X4 U3714 ( .B1(n2501), .B2(net255318), .A(net255319), .ZN(n2529) );
  NAND2_X4 U3715 ( .A1(net253657), .A2(net253656), .ZN(net253411) );
  NAND2_X4 U3716 ( .A1(n3909), .A2(n3913), .ZN(n3992) );
  NAND3_X2 U3717 ( .A1(n2334), .A2(n2333), .A3(n1414), .ZN(net255426) );
  NAND2_X4 U3718 ( .A1(n3243), .A2(n1978), .ZN(n3453) );
  NAND3_X1 U3719 ( .A1(n2612), .A2(n2613), .A3(n2682), .ZN(n2614) );
  NAND3_X2 U3720 ( .A1(n1873), .A2(n1392), .A3(n2682), .ZN(n2678) );
  NAND2_X4 U3721 ( .A1(n3926), .A2(n3793), .ZN(n3919) );
  NAND2_X4 U3722 ( .A1(n2551), .A2(n2552), .ZN(n2652) );
  NAND2_X4 U3723 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
  NAND2_X4 U3724 ( .A1(n3197), .A2(n3196), .ZN(n3199) );
  NAND2_X4 U3726 ( .A1(n1809), .A2(n3380), .ZN(n3604) );
  NAND3_X2 U3727 ( .A1(net256909), .A2(n2443), .A3(n2441), .ZN(n2378) );
  INV_X8 U3728 ( .A(net253820), .ZN(net253816) );
  NAND2_X4 U3729 ( .A1(n3172), .A2(n1583), .ZN(n3271) );
  NAND3_X2 U3730 ( .A1(n3525), .A2(n1842), .A3(n3520), .ZN(n3172) );
  OAI21_X4 U3731 ( .B1(n2815), .B2(n2879), .A(n2814), .ZN(n2840) );
  INV_X8 U3732 ( .A(n2808), .ZN(n2879) );
  NAND2_X4 U3733 ( .A1(n2810), .A2(n2811), .ZN(n2881) );
  NAND2_X4 U3734 ( .A1(net255383), .A2(n2466), .ZN(n2579) );
  NAND2_X4 U3735 ( .A1(net253547), .A2(net253177), .ZN(n3774) );
  NAND2_X4 U3736 ( .A1(net254094), .A2(net254085), .ZN(n3709) );
  NAND2_X4 U3737 ( .A1(n2206), .A2(net255434), .ZN(net255433) );
  NAND3_X1 U3739 ( .A1(n2506), .A2(n1873), .A3(n2613), .ZN(n2507) );
  NAND2_X4 U3740 ( .A1(net254283), .A2(n3251), .ZN(net253764) );
  NAND2_X4 U3741 ( .A1(n2492), .A2(n2491), .ZN(n2570) );
  NAND2_X4 U3742 ( .A1(n2638), .A2(n2637), .ZN(n2656) );
  NAND2_X4 U3743 ( .A1(n2739), .A2(n2737), .ZN(n2636) );
  NAND3_X2 U3744 ( .A1(net255916), .A2(net257401), .A3(net255915), .ZN(
        net255856) );
  NAND2_X4 U3745 ( .A1(n1890), .A2(n2394), .ZN(n2536) );
  NAND3_X4 U3746 ( .A1(n1803), .A2(n3506), .A3(n3787), .ZN(net253179) );
  NAND2_X4 U3747 ( .A1(n1785), .A2(n1143), .ZN(n3780) );
  NAND2_X4 U3748 ( .A1(n2464), .A2(n1796), .ZN(n2612) );
  NAND2_X4 U3749 ( .A1(n2959), .A2(net254675), .ZN(net254459) );
  NAND2_X4 U3750 ( .A1(n2750), .A2(n2751), .ZN(n2755) );
  NAND2_X4 U3751 ( .A1(n3381), .A2(n3382), .ZN(n3550) );
  NAND2_X4 U3752 ( .A1(net254761), .A2(net256306), .ZN(n3031) );
  NAND2_X4 U3753 ( .A1(n2920), .A2(n1416), .ZN(n3025) );
  NAND3_X1 U3754 ( .A1(net257590), .A2(n1258), .A3(n2182), .ZN(n2145) );
  NAND3_X1 U3755 ( .A1(n1258), .A2(net255626), .A3(net255434), .ZN(n2246) );
  NAND2_X4 U3756 ( .A1(net256033), .A2(net256032), .ZN(net255611) );
  NAND2_X4 U3757 ( .A1(control[1]), .A2(net256087), .ZN(net253064) );
  INV_X32 U3758 ( .A(net256167), .ZN(net256165) );
  INV_X16 U3759 ( .A(net253271), .ZN(net256167) );
  INV_X32 U3760 ( .A(net256139), .ZN(net256135) );
  INV_X32 U3761 ( .A(control[0]), .ZN(net256089) );
  NAND2_X2 U3762 ( .A1(a[0]), .A2(net256151), .ZN(n3410) );
  INV_X4 U3763 ( .A(n3410), .ZN(n2803) );
  MUX2_X2 U3764 ( .A(product_in[0]), .B(n2803), .S(net256097), .Z(
        product_out[0]) );
  NAND2_X2 U3765 ( .A1(a[1]), .A2(net256147), .ZN(n2009) );
  XOR2_X2 U3766 ( .A(n2010), .B(n2009), .Z(n3510) );
  MUX2_X2 U3767 ( .A(product_in[1]), .B(n3510), .S(net256099), .Z(
        product_out[1]) );
  NAND2_X2 U3768 ( .A1(a[0]), .A2(net256117), .ZN(n2016) );
  INV_X4 U3769 ( .A(n2016), .ZN(n2118) );
  INV_X4 U3770 ( .A(n2019), .ZN(n3692) );
  MUX2_X2 U3771 ( .A(product_in[2]), .B(n3692), .S(net256097), .Z(
        product_out[2]) );
  NAND3_X2 U3772 ( .A1(a[1]), .A2(n4098), .A3(net257127), .ZN(n2027) );
  NAND2_X2 U3773 ( .A1(n2062), .A2(n2063), .ZN(n2026) );
  NAND4_X2 U3774 ( .A1(b[24]), .A2(n1466), .A3(a[1]), .A4(net257677), .ZN(
        n2024) );
  NAND4_X2 U3775 ( .A1(b[16]), .A2(control[0]), .A3(a[1]), .A4(net257782), 
        .ZN(n2023) );
  NAND4_X2 U3776 ( .A1(n2024), .A2(n2023), .A3(n2022), .A4(n2021), .ZN(n2025)
         );
  NOR2_X4 U3777 ( .A1(n2093), .A2(n2092), .ZN(n2041) );
  NOR2_X4 U3778 ( .A1(n2095), .A2(n2094), .ZN(n2040) );
  NAND2_X2 U3779 ( .A1(n2043), .A2(n2042), .ZN(n2045) );
  NAND2_X2 U3780 ( .A1(a[1]), .A2(net256119), .ZN(n2046) );
  INV_X4 U3781 ( .A(n2046), .ZN(n2058) );
  NAND2_X2 U3782 ( .A1(n2045), .A2(n2044), .ZN(n2056) );
  NAND2_X2 U3783 ( .A1(n2056), .A2(n2046), .ZN(n2192) );
  XNOR2_X2 U3784 ( .A(n2048), .B(n2059), .ZN(n2052) );
  NAND2_X2 U3785 ( .A1(net257721), .A2(net256371), .ZN(net253308) );
  AOI22_X2 U3786 ( .A1(b[27]), .A2(net253067), .B1(b[19]), .B2(n1922), .ZN(
        n2050) );
  AOI22_X2 U3787 ( .A1(b[3]), .A2(net256099), .B1(b[11]), .B2(net256183), .ZN(
        n2049) );
  NAND2_X2 U3788 ( .A1(n2050), .A2(n2049), .ZN(net253237) );
  NAND2_X2 U3789 ( .A1(a[0]), .A2(net256135), .ZN(n2051) );
  NAND2_X2 U3790 ( .A1(n2052), .A2(n2051), .ZN(n2055) );
  INV_X4 U3791 ( .A(n2051), .ZN(n2054) );
  INV_X4 U3792 ( .A(n2052), .ZN(n2053) );
  NAND2_X2 U3793 ( .A1(n2055), .A2(n2183), .ZN(n3762) );
  INV_X4 U3794 ( .A(n3762), .ZN(n2418) );
  MUX2_X2 U3795 ( .A(product_in[3]), .B(n2418), .S(net256099), .Z(
        product_out[3]) );
  INV_X4 U3796 ( .A(n2192), .ZN(n2060) );
  NAND2_X2 U3797 ( .A1(n2118), .A2(n4096), .ZN(n2059) );
  OAI21_X4 U3798 ( .B1(n2065), .B2(n2064), .A(a[3]), .ZN(n2066) );
  INV_X4 U3799 ( .A(net255936), .ZN(net255790) );
  XNOR2_X2 U3800 ( .A(n2069), .B(n2068), .ZN(n2076) );
  XNOR2_X2 U3801 ( .A(n2075), .B(net257565), .ZN(n2120) );
  XNOR2_X2 U3802 ( .A(n2078), .B(n2077), .ZN(n2080) );
  NAND2_X2 U3803 ( .A1(a[1]), .A2(net256137), .ZN(n2079) );
  INV_X4 U3804 ( .A(n2079), .ZN(n2081) );
  NAND2_X2 U3805 ( .A1(n2081), .A2(n2080), .ZN(n2186) );
  NAND2_X2 U3806 ( .A1(b[12]), .A2(net256183), .ZN(n2085) );
  NAND2_X2 U3807 ( .A1(b[4]), .A2(net256099), .ZN(n2084) );
  AOI22_X2 U3808 ( .A1(b[28]), .A2(net253067), .B1(b[20]), .B2(n1922), .ZN(
        n2083) );
  NAND2_X2 U3809 ( .A1(a[0]), .A2(net253231), .ZN(n2086) );
  NAND2_X2 U3810 ( .A1(n1923), .A2(n2086), .ZN(n2090) );
  INV_X4 U3811 ( .A(n2086), .ZN(n2089) );
  INV_X4 U3812 ( .A(n2125), .ZN(n2124) );
  NAND2_X2 U3813 ( .A1(a[3]), .A2(net256119), .ZN(n2146) );
  INV_X4 U3814 ( .A(n2146), .ZN(n2116) );
  NAND4_X2 U3815 ( .A1(n2099), .A2(n2098), .A3(n2097), .A4(n2096), .ZN(n2198)
         );
  NAND2_X2 U3816 ( .A1(n2198), .A2(net255936), .ZN(n2111) );
  NAND3_X2 U3817 ( .A1(n2104), .A2(n2105), .A3(n1954), .ZN(n2106) );
  INV_X4 U3818 ( .A(n2106), .ZN(n2197) );
  NAND3_X2 U3819 ( .A1(n2107), .A2(net255540), .A3(n1802), .ZN(n2108) );
  NAND2_X2 U3820 ( .A1(n2116), .A2(n2110), .ZN(n2113) );
  INV_X4 U3821 ( .A(n2111), .ZN(n2370) );
  NAND2_X2 U3822 ( .A1(n2113), .A2(n2112), .ZN(n2114) );
  NAND2_X2 U3823 ( .A1(n2114), .A2(n1835), .ZN(n2139) );
  OAI21_X4 U3824 ( .B1(n2115), .B2(n2116), .A(n2139), .ZN(n2154) );
  NAND3_X2 U3825 ( .A1(n1952), .A2(n2141), .A3(n2140), .ZN(n2153) );
  INV_X4 U3826 ( .A(n1979), .ZN(n2157) );
  NAND2_X2 U3827 ( .A1(a[1]), .A2(net256127), .ZN(n2128) );
  OAI21_X4 U3828 ( .B1(n2127), .B2(n2126), .A(n2128), .ZN(n2217) );
  INV_X4 U3829 ( .A(n2128), .ZN(n2264) );
  NAND2_X2 U3830 ( .A1(n2217), .A2(n2268), .ZN(n2130) );
  XNOR2_X2 U3831 ( .A(n2130), .B(n2164), .ZN(n2135) );
  NAND2_X2 U3832 ( .A1(b[13]), .A2(net256183), .ZN(n2133) );
  NAND2_X2 U3833 ( .A1(b[5]), .A2(net256099), .ZN(n2132) );
  AOI22_X2 U3834 ( .A1(b[29]), .A2(net253067), .B1(b[21]), .B2(n1922), .ZN(
        n2131) );
  NAND3_X4 U3835 ( .A1(n2133), .A2(n2132), .A3(n2131), .ZN(net253103) );
  NAND2_X2 U3836 ( .A1(a[0]), .A2(net256105), .ZN(n2134) );
  INV_X4 U3837 ( .A(n2134), .ZN(n2137) );
  INV_X4 U3838 ( .A(n2135), .ZN(n2136) );
  INV_X4 U3839 ( .A(n3918), .ZN(n2566) );
  MUX2_X2 U3840 ( .A(product_in[5]), .B(n2566), .S(net256099), .Z(
        product_out[5]) );
  NAND2_X2 U3841 ( .A1(a[1]), .A2(net253103), .ZN(n2220) );
  INV_X4 U3842 ( .A(a[6]), .ZN(net255718) );
  NAND2_X2 U3843 ( .A1(a[3]), .A2(net256137), .ZN(n2150) );
  INV_X4 U3844 ( .A(n2150), .ZN(n2182) );
  NAND2_X2 U3845 ( .A1(n2143), .A2(n2142), .ZN(n2148) );
  XNOR2_X2 U3846 ( .A(n2145), .B(n2144), .ZN(n2151) );
  XNOR2_X2 U3847 ( .A(net255725), .B(n2149), .ZN(n2180) );
  OAI21_X4 U3848 ( .B1(n2160), .B2(n2159), .A(n2158), .ZN(n2223) );
  XNOR2_X2 U3849 ( .A(n2223), .B(n2226), .ZN(n2161) );
  INV_X4 U3850 ( .A(n2224), .ZN(n2163) );
  NAND2_X2 U3851 ( .A1(n2266), .A2(n2217), .ZN(n2230) );
  NAND2_X2 U3852 ( .A1(n2220), .A2(n2167), .ZN(n2169) );
  XNOR2_X2 U3853 ( .A(n2170), .B(n2221), .ZN(n2175) );
  NAND2_X2 U3854 ( .A1(b[14]), .A2(net256183), .ZN(n2173) );
  NAND2_X2 U3855 ( .A1(b[6]), .A2(net256099), .ZN(n2172) );
  AOI22_X2 U3856 ( .A1(b[30]), .A2(net253067), .B1(b[22]), .B2(n1922), .ZN(
        n2171) );
  NAND2_X2 U3857 ( .A1(a[0]), .A2(net256173), .ZN(n2174) );
  INV_X4 U3859 ( .A(n2174), .ZN(n2177) );
  INV_X4 U3860 ( .A(n2175), .ZN(n2176) );
  INV_X4 U3861 ( .A(n2179), .ZN(n3983) );
  MUX2_X2 U3862 ( .A(product_in[6]), .B(n3983), .S(net256097), .Z(
        product_out[6]) );
  NAND2_X2 U3863 ( .A1(n2182), .A2(n2181), .ZN(n2319) );
  NOR2_X4 U3864 ( .A1(n2184), .A2(n2183), .ZN(n2188) );
  OAI21_X4 U3865 ( .B1(n2195), .B2(n2196), .A(n2194), .ZN(net255626) );
  INV_X4 U3866 ( .A(n2198), .ZN(n2199) );
  OAI21_X4 U3867 ( .B1(net255785), .B2(n1858), .A(n2200), .ZN(net255727) );
  INV_X4 U3868 ( .A(net255727), .ZN(net255776) );
  NAND2_X2 U3869 ( .A1(n1840), .A2(net255533), .ZN(n2202) );
  INV_X4 U3870 ( .A(n2204), .ZN(n2250) );
  INV_X4 U3871 ( .A(net255726), .ZN(net255777) );
  NAND2_X2 U3872 ( .A1(a[5]), .A2(net256119), .ZN(net255775) );
  NAND2_X2 U3873 ( .A1(a[4]), .A2(net256137), .ZN(n2207) );
  NAND2_X2 U3875 ( .A1(n2322), .A2(n2320), .ZN(n2209) );
  INV_X4 U3877 ( .A(n2212), .ZN(n2214) );
  INV_X4 U3878 ( .A(n2268), .ZN(n2216) );
  XNOR2_X2 U3879 ( .A(n1912), .B(n1824), .ZN(n2311) );
  INV_X4 U3880 ( .A(n2220), .ZN(n2229) );
  AOI21_X2 U3881 ( .B1(n1805), .B2(n2315), .A(n2229), .ZN(n2222) );
  XNOR2_X2 U3882 ( .A(n2225), .B(n2224), .ZN(n2227) );
  XNOR2_X2 U3883 ( .A(n2227), .B(n2226), .ZN(n2228) );
  NAND2_X2 U3884 ( .A1(n2229), .A2(n2228), .ZN(n2231) );
  XNOR2_X2 U3885 ( .A(n2231), .B(n2230), .ZN(n2232) );
  NAND2_X2 U3886 ( .A1(n2308), .A2(n2306), .ZN(n2234) );
  NAND2_X2 U3887 ( .A1(a[1]), .A2(net256175), .ZN(n2236) );
  INV_X4 U3888 ( .A(n2236), .ZN(n2239) );
  INV_X4 U3889 ( .A(n2237), .ZN(n2238) );
  XNOR2_X2 U3890 ( .A(n2240), .B(n2292), .ZN(n2241) );
  INV_X4 U3891 ( .A(n2241), .ZN(n2299) );
  NAND2_X2 U3892 ( .A1(b[15]), .A2(net256183), .ZN(n2244) );
  NAND2_X2 U3893 ( .A1(b[7]), .A2(net256099), .ZN(n2243) );
  AOI22_X2 U3894 ( .A1(b[31]), .A2(net253067), .B1(b[23]), .B2(n1922), .ZN(
        n2242) );
  XNOR2_X2 U3895 ( .A(n2299), .B(n1424), .ZN(n3397) );
  INV_X4 U3896 ( .A(n3397), .ZN(n4068) );
  MUX2_X2 U3897 ( .A(product_in[7]), .B(n4068), .S(net256097), .Z(
        product_out[7]) );
  NAND2_X2 U3898 ( .A1(product_in[8]), .A2(net256095), .ZN(n2301) );
  NAND2_X2 U3899 ( .A1(n1390), .A2(net256175), .ZN(n2288) );
  INV_X4 U3900 ( .A(n2288), .ZN(n2287) );
  NAND2_X2 U3901 ( .A1(a[6]), .A2(net256119), .ZN(net255624) );
  INV_X4 U3902 ( .A(a[7]), .ZN(n2248) );
  INV_X4 U3903 ( .A(a[8]), .ZN(n2434) );
  NOR2_X4 U3904 ( .A1(n2434), .A2(n2248), .ZN(net255720) );
  NOR2_X4 U3905 ( .A1(net255718), .A2(n2248), .ZN(n2249) );
  NAND2_X2 U3906 ( .A1(n2250), .A2(n2445), .ZN(n2255) );
  NOR2_X4 U3907 ( .A1(n1411), .A2(n2377), .ZN(n2252) );
  NAND2_X2 U3908 ( .A1(a[5]), .A2(net256137), .ZN(net255703) );
  XNOR2_X2 U3909 ( .A(n2258), .B(net255699), .ZN(n2260) );
  NAND2_X2 U3910 ( .A1(a[4]), .A2(net256125), .ZN(n2259) );
  INV_X4 U3911 ( .A(n2259), .ZN(n2262) );
  INV_X4 U3912 ( .A(n2260), .ZN(n2261) );
  INV_X4 U3913 ( .A(n2263), .ZN(n2275) );
  NAND3_X2 U3914 ( .A1(n2269), .A2(n2268), .A3(n2267), .ZN(n2271) );
  NAND2_X2 U3915 ( .A1(n2313), .A2(n2315), .ZN(n2273) );
  NAND2_X2 U3916 ( .A1(a[3]), .A2(net256105), .ZN(n2276) );
  INV_X4 U3917 ( .A(n2276), .ZN(n2277) );
  NAND2_X2 U3918 ( .A1(n2309), .A2(n2360), .ZN(n2285) );
  XNOR2_X2 U3919 ( .A(n2215), .B(n2279), .ZN(n2280) );
  NAND2_X2 U3920 ( .A1(n2281), .A2(n2307), .ZN(n2283) );
  XNOR2_X2 U3921 ( .A(n2285), .B(n2284), .ZN(n2289) );
  INV_X4 U3922 ( .A(n1831), .ZN(n2286) );
  OAI21_X4 U3923 ( .B1(n2293), .B2(n2292), .A(n2291), .ZN(n2304) );
  XNOR2_X2 U3924 ( .A(n2294), .B(n2304), .ZN(n2297) );
  INV_X4 U3925 ( .A(n2297), .ZN(n2295) );
  NAND2_X2 U3926 ( .A1(a[1]), .A2(net256165), .ZN(n2296) );
  INV_X4 U3927 ( .A(n2296), .ZN(n2298) );
  NAND2_X2 U3928 ( .A1(n2298), .A2(n2297), .ZN(n2348) );
  NAND2_X2 U3929 ( .A1(n1424), .A2(n2299), .ZN(n2349) );
  XNOR2_X2 U3930 ( .A(n2300), .B(n2349), .ZN(n3406) );
  INV_X4 U3931 ( .A(n2301), .ZN(n2303) );
  INV_X4 U3932 ( .A(n2416), .ZN(n2357) );
  NAND2_X2 U3933 ( .A1(product_in[9]), .A2(net256095), .ZN(n2354) );
  INV_X4 U3934 ( .A(n2354), .ZN(n2352) );
  INV_X4 U3935 ( .A(n3510), .ZN(n2351) );
  NAND3_X2 U3936 ( .A1(n2308), .A2(n2307), .A3(n2306), .ZN(n2310) );
  NAND2_X2 U3937 ( .A1(n2360), .A2(n2361), .ZN(n2341) );
  NAND2_X2 U3938 ( .A1(a[4]), .A2(net256105), .ZN(n2337) );
  NAND3_X2 U3939 ( .A1(n2315), .A2(n2314), .A3(n2313), .ZN(n2317) );
  INV_X4 U3940 ( .A(n2427), .ZN(n2318) );
  NAND3_X2 U3941 ( .A1(n1829), .A2(n2320), .A3(n2319), .ZN(net255322) );
  INV_X4 U3942 ( .A(n2379), .ZN(n2324) );
  INV_X4 U3943 ( .A(n2435), .ZN(n2375) );
  INV_X4 U3944 ( .A(net255606), .ZN(net255605) );
  AOI21_X4 U3945 ( .B1(n1858), .B2(n1840), .A(net255605), .ZN(n2330) );
  NAND3_X2 U3946 ( .A1(n1875), .A2(n2371), .A3(n2330), .ZN(n2331) );
  NAND2_X2 U3947 ( .A1(a[5]), .A2(net256125), .ZN(net255582) );
  INV_X4 U3948 ( .A(net255582), .ZN(net255453) );
  INV_X4 U3949 ( .A(n2337), .ZN(n2339) );
  NAND2_X2 U3950 ( .A1(n2362), .A2(n2535), .ZN(n2340) );
  XNOR2_X2 U3951 ( .A(n2341), .B(n2340), .ZN(n2344) );
  NAND2_X2 U3952 ( .A1(a[3]), .A2(net256175), .ZN(n2343) );
  INV_X4 U3953 ( .A(n2343), .ZN(n2345) );
  NAND2_X2 U3954 ( .A1(n2496), .A2(n2420), .ZN(n2405) );
  XNOR2_X2 U3955 ( .A(n2346), .B(n2405), .ZN(n2402) );
  OAI21_X4 U3956 ( .B1(n2350), .B2(n2349), .A(n2348), .ZN(n2401) );
  XNOR2_X2 U3957 ( .A(n2402), .B(n2401), .ZN(n3513) );
  NAND2_X2 U3958 ( .A1(n2352), .A2(n2353), .ZN(n2415) );
  INV_X4 U3959 ( .A(n2353), .ZN(n2355) );
  XNOR2_X2 U3960 ( .A(n2357), .B(n2356), .ZN(product_out[9]) );
  INV_X4 U3961 ( .A(a[3]), .ZN(net255484) );
  INV_X4 U3962 ( .A(n2496), .ZN(n2359) );
  OAI21_X4 U3963 ( .B1(n2359), .B2(n2358), .A(n2420), .ZN(n2398) );
  INV_X4 U3964 ( .A(n2360), .ZN(n2364) );
  OAI21_X4 U3965 ( .B1(n2363), .B2(n2364), .A(n2362), .ZN(n2629) );
  NAND2_X2 U3966 ( .A1(a[7]), .A2(net256137), .ZN(net255505) );
  INV_X4 U3967 ( .A(net255505), .ZN(net255506) );
  AND2_X2 U3968 ( .A1(net255426), .A2(net255434), .ZN(n2367) );
  NAND3_X2 U3969 ( .A1(net255542), .A2(n2368), .A3(n2505), .ZN(n2390) );
  NOR2_X4 U3970 ( .A1(n2374), .A2(n2373), .ZN(n2380) );
  AOI21_X4 U3971 ( .B1(n2380), .B2(n2379), .A(n2378), .ZN(n2385) );
  INV_X4 U3972 ( .A(n2382), .ZN(n2381) );
  NAND3_X4 U3973 ( .A1(n2381), .A2(a[9]), .A3(net257586), .ZN(n2688) );
  NAND2_X2 U3974 ( .A1(a[9]), .A2(net257586), .ZN(n2383) );
  NAND2_X2 U3975 ( .A1(a[8]), .A2(net256119), .ZN(n2386) );
  INV_X4 U3976 ( .A(n2386), .ZN(n2388) );
  NAND2_X2 U3977 ( .A1(a[5]), .A2(net256105), .ZN(n2392) );
  INV_X4 U3978 ( .A(n2392), .ZN(n2394) );
  XNOR2_X2 U3979 ( .A(n2396), .B(n2395), .ZN(net255490) );
  NAND3_X2 U3980 ( .A1(n4113), .A2(a[4]), .A3(net256173), .ZN(n2497) );
  INV_X4 U3981 ( .A(net255490), .ZN(net255489) );
  XNOR2_X2 U3982 ( .A(n2397), .B(n2398), .ZN(n2400) );
  OAI21_X4 U3983 ( .B1(net256167), .B2(net255484), .A(n2399), .ZN(n2558) );
  NAND2_X2 U3984 ( .A1(n2558), .A2(n2555), .ZN(n2408) );
  INV_X4 U3985 ( .A(n2403), .ZN(n2407) );
  XNOR2_X2 U3986 ( .A(n2405), .B(n2404), .ZN(n2406) );
  NAND2_X2 U3987 ( .A1(n2407), .A2(n2406), .ZN(n2554) );
  XNOR2_X2 U3988 ( .A(n2408), .B(n2476), .ZN(n3691) );
  INV_X4 U3989 ( .A(n3691), .ZN(n2995) );
  NAND2_X2 U3990 ( .A1(n3692), .A2(net256183), .ZN(n2409) );
  NAND2_X2 U3991 ( .A1(product_in[10]), .A2(net256095), .ZN(n2410) );
  INV_X4 U3992 ( .A(n2409), .ZN(n2412) );
  INV_X4 U3993 ( .A(n2410), .ZN(n2411) );
  NAND2_X2 U3994 ( .A1(n2412), .A2(n2411), .ZN(n2481) );
  OAI21_X4 U3996 ( .B1(n2417), .B2(n2416), .A(n2415), .ZN(n2480) );
  NAND2_X2 U3997 ( .A1(n2418), .A2(net256183), .ZN(n2488) );
  NAND2_X2 U3998 ( .A1(n2423), .A2(n1144), .ZN(n2472) );
  INV_X4 U3999 ( .A(net255458), .ZN(net255457) );
  NOR2_X4 U4000 ( .A1(n2425), .A2(net255453), .ZN(n2429) );
  NAND2_X2 U4001 ( .A1(a[7]), .A2(net256125), .ZN(net255376) );
  INV_X4 U4002 ( .A(net255376), .ZN(net255379) );
  OAI21_X4 U4003 ( .B1(net255429), .B2(net255428), .A(net255430), .ZN(n2504)
         );
  NAND2_X2 U4004 ( .A1(n2435), .A2(n2434), .ZN(n2438) );
  NAND3_X2 U4005 ( .A1(n2437), .A2(n2438), .A3(n2439), .ZN(n2583) );
  NAND2_X2 U4006 ( .A1(n2583), .A2(n2443), .ZN(n2517) );
  NAND2_X2 U4007 ( .A1(n2584), .A2(n2517), .ZN(n2455) );
  INV_X4 U4008 ( .A(n2455), .ZN(n2449) );
  NAND3_X2 U4009 ( .A1(n2440), .A2(n2201), .A3(n2441), .ZN(n2699) );
  XNOR2_X2 U4010 ( .A(n2513), .B(n2514), .ZN(n2588) );
  INV_X4 U4011 ( .A(n2588), .ZN(n2452) );
  INV_X4 U4012 ( .A(n2688), .ZN(n2515) );
  XNOR2_X2 U4013 ( .A(n2450), .B(n2515), .ZN(n2453) );
  OAI21_X4 U4014 ( .B1(n2452), .B2(n2451), .A(n2453), .ZN(n2458) );
  NAND2_X2 U4015 ( .A1(n2454), .A2(n2453), .ZN(n2457) );
  NAND2_X2 U4016 ( .A1(a[9]), .A2(net256119), .ZN(n2460) );
  INV_X4 U4017 ( .A(n2460), .ZN(n2463) );
  XNOR2_X2 U4019 ( .A(net255374), .B(n1110), .ZN(n2469) );
  NAND2_X2 U4020 ( .A1(a[6]), .A2(net256105), .ZN(n2468) );
  INV_X4 U4021 ( .A(n2468), .ZN(n2470) );
  NAND2_X2 U4022 ( .A1(a[5]), .A2(net256175), .ZN(n2493) );
  XNOR2_X2 U4023 ( .A(n2573), .B(n2473), .ZN(n2559) );
  INV_X4 U4024 ( .A(n1891), .ZN(n2475) );
  NAND2_X2 U4025 ( .A1(a[4]), .A2(net256165), .ZN(n2474) );
  INV_X4 U4026 ( .A(n2474), .ZN(n2560) );
  NAND2_X2 U4027 ( .A1(product_in[11]), .A2(net256095), .ZN(n2487) );
  INV_X4 U4028 ( .A(n2487), .ZN(n2478) );
  XNOR2_X2 U4029 ( .A(n2479), .B(n2478), .ZN(n2486) );
  INV_X4 U4030 ( .A(n2480), .ZN(n2483) );
  OAI21_X4 U4031 ( .B1(n2483), .B2(n2482), .A(n2481), .ZN(n2484) );
  INV_X4 U4032 ( .A(n2484), .ZN(n2485) );
  NOR2_X4 U4033 ( .A1(n2486), .A2(n2485), .ZN(n2490) );
  NOR2_X4 U4034 ( .A1(n2490), .A2(n2489), .ZN(n2646) );
  INV_X4 U4035 ( .A(n2493), .ZN(n2492) );
  INV_X4 U4036 ( .A(n2570), .ZN(n2664) );
  INV_X4 U4037 ( .A(n2499), .ZN(n2663) );
  NAND2_X2 U4038 ( .A1(a[7]), .A2(net256105), .ZN(n2532) );
  INV_X4 U4039 ( .A(n2532), .ZN(n2530) );
  NOR2_X4 U4040 ( .A1(n2753), .A2(n2749), .ZN(n2501) );
  NAND3_X2 U4041 ( .A1(n1953), .A2(n1392), .A3(n2503), .ZN(n2509) );
  NAND4_X2 U4042 ( .A1(n2509), .A2(n2681), .A3(n2508), .A4(n2507), .ZN(n2526)
         );
  INV_X4 U4043 ( .A(a[11]), .ZN(n2511) );
  NOR2_X4 U4044 ( .A1(n2511), .A2(net254628), .ZN(n2510) );
  OAI21_X4 U4045 ( .B1(net257585), .B2(n2511), .A(n2590), .ZN(n2512) );
  NAND2_X2 U4046 ( .A1(n2514), .A2(n2513), .ZN(n2687) );
  INV_X4 U4047 ( .A(n2687), .ZN(n2596) );
  NOR2_X4 U4048 ( .A1(n2596), .A2(n2515), .ZN(n2520) );
  NAND4_X2 U4049 ( .A1(n2699), .A2(n2517), .A3(n2518), .A4(n2700), .ZN(n2519)
         );
  NAND2_X2 U4050 ( .A1(a[10]), .A2(net256119), .ZN(n2522) );
  INV_X4 U4051 ( .A(n2522), .ZN(n2524) );
  XNOR2_X2 U4052 ( .A(n2526), .B(n2683), .ZN(n2528) );
  NAND2_X2 U4053 ( .A1(a[9]), .A2(net256135), .ZN(n2527) );
  INV_X4 U4054 ( .A(n2527), .ZN(n2577) );
  INV_X4 U4055 ( .A(n2528), .ZN(n2576) );
  XNOR2_X2 U4056 ( .A(n2529), .B(n1420), .ZN(net255231) );
  NAND2_X2 U4057 ( .A1(a[8]), .A2(net256125), .ZN(net255232) );
  XNOR2_X2 U4058 ( .A(net255284), .B(net256860), .ZN(n2531) );
  NOR2_X4 U4059 ( .A1(n1260), .A2(n2668), .ZN(n2542) );
  INV_X4 U4060 ( .A(n2534), .ZN(n2626) );
  XNOR2_X2 U4061 ( .A(n2542), .B(n1867), .ZN(n2543) );
  NAND2_X2 U4062 ( .A1(n2662), .A2(n2659), .ZN(n2547) );
  XNOR2_X2 U4063 ( .A(n2544), .B(n2547), .ZN(n2545) );
  NAND2_X2 U4064 ( .A1(a[5]), .A2(net256165), .ZN(n2546) );
  INV_X4 U4065 ( .A(n2546), .ZN(n2552) );
  INV_X4 U4066 ( .A(n2547), .ZN(n2550) );
  XNOR2_X2 U4067 ( .A(n2550), .B(n2549), .ZN(n2551) );
  AOI21_X4 U4068 ( .B1(n2558), .B2(n2557), .A(n2556), .ZN(n2655) );
  OAI21_X4 U4069 ( .B1(n2655), .B2(n2654), .A(n2653), .ZN(n2567) );
  XNOR2_X2 U4070 ( .A(n2561), .B(n1813), .ZN(n3794) );
  INV_X4 U4071 ( .A(n3794), .ZN(n3169) );
  NAND2_X2 U4072 ( .A1(product_in[12]), .A2(net256095), .ZN(n2562) );
  INV_X4 U4073 ( .A(net255247), .ZN(net255244) );
  INV_X4 U4074 ( .A(n2562), .ZN(n2563) );
  NAND2_X2 U4075 ( .A1(net255244), .A2(n2563), .ZN(n2644) );
  INV_X4 U4076 ( .A(n2645), .ZN(n2565) );
  NAND2_X2 U4077 ( .A1(n2566), .A2(net256183), .ZN(n2647) );
  INV_X4 U4078 ( .A(n2657), .ZN(n2569) );
  NAND2_X2 U4080 ( .A1(a[6]), .A2(net256165), .ZN(n2638) );
  OAI21_X4 U4081 ( .B1(n1811), .B2(n2570), .A(n2659), .ZN(n2571) );
  NAND3_X2 U4082 ( .A1(n2662), .A2(n2573), .A3(n2572), .ZN(n2739) );
  INV_X4 U4083 ( .A(net255232), .ZN(net255106) );
  NOR3_X4 U4084 ( .A1(n2575), .A2(net255218), .A3(net255217), .ZN(n2582) );
  OAI21_X4 U4085 ( .B1(n2581), .B2(n2582), .A(n2674), .ZN(n2621) );
  NAND2_X2 U4086 ( .A1(a[11]), .A2(net256119), .ZN(n2605) );
  INV_X4 U4087 ( .A(n2583), .ZN(n2585) );
  OAI21_X4 U4088 ( .B1(n2586), .B2(n2585), .A(n2584), .ZN(n2697) );
  NAND3_X2 U4089 ( .A1(n2700), .A2(n2699), .A3(n2587), .ZN(n2598) );
  NAND2_X2 U4090 ( .A1(a[12]), .A2(net257586), .ZN(n2589) );
  INV_X4 U4091 ( .A(n2686), .ZN(n2595) );
  NOR2_X4 U4092 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  NAND3_X2 U4093 ( .A1(n2598), .A2(n2688), .A3(n2597), .ZN(n2599) );
  NAND2_X2 U4094 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  OAI21_X4 U4095 ( .B1(n2603), .B2(n2602), .A(n2601), .ZN(n2604) );
  NAND2_X2 U4096 ( .A1(n2605), .A2(n2604), .ZN(n2608) );
  INV_X4 U4097 ( .A(n2605), .ZN(n2606) );
  INV_X4 U4098 ( .A(n2679), .ZN(n2616) );
  XNOR2_X2 U4099 ( .A(n2617), .B(n2759), .ZN(n2619) );
  INV_X4 U4100 ( .A(n2618), .ZN(n2751) );
  NAND2_X2 U4101 ( .A1(n2673), .A2(n2755), .ZN(n2620) );
  NAND2_X2 U4102 ( .A1(a[9]), .A2(net256125), .ZN(net255167) );
  NAND2_X2 U4103 ( .A1(a[8]), .A2(net256105), .ZN(n2622) );
  INV_X4 U4104 ( .A(n2622), .ZN(n2625) );
  OAI21_X4 U4105 ( .B1(n2627), .B2(n2626), .A(n2630), .ZN(n2669) );
  NAND3_X4 U4106 ( .A1(n2630), .A2(n2628), .A3(n1897), .ZN(n2945) );
  NAND2_X2 U4107 ( .A1(a[7]), .A2(net256175), .ZN(n2632) );
  INV_X4 U4108 ( .A(n2632), .ZN(n2634) );
  XNOR2_X2 U4109 ( .A(n2636), .B(n2635), .ZN(n2639) );
  INV_X4 U4110 ( .A(n1934), .ZN(n2637) );
  INV_X4 U4111 ( .A(n1944), .ZN(n2642) );
  XNOR2_X2 U4112 ( .A(n2643), .B(n1408), .ZN(n2649) );
  OAI21_X4 U4113 ( .B1(n2646), .B2(n2645), .A(n2644), .ZN(n2650) );
  INV_X4 U4114 ( .A(n2647), .ZN(n2648) );
  NAND2_X2 U4115 ( .A1(n1408), .A2(n2648), .ZN(n2851) );
  INV_X4 U4116 ( .A(n2649), .ZN(n2651) );
  NAND2_X2 U4117 ( .A1(a[8]), .A2(net256175), .ZN(n2718) );
  INV_X4 U4118 ( .A(n2674), .ZN(n2756) );
  INV_X4 U4119 ( .A(n2675), .ZN(n2752) );
  NOR2_X4 U4120 ( .A1(n2753), .A2(n2752), .ZN(n2677) );
  INV_X4 U4121 ( .A(n2678), .ZN(n2680) );
  NAND2_X2 U4122 ( .A1(n2680), .A2(n2679), .ZN(n2888) );
  INV_X4 U4123 ( .A(n2681), .ZN(n2684) );
  OAI21_X4 U4124 ( .B1(n2684), .B2(n2683), .A(n2682), .ZN(n2890) );
  INV_X4 U4125 ( .A(n2759), .ZN(n2886) );
  NAND3_X2 U4126 ( .A1(n1970), .A2(n2690), .A3(n2689), .ZN(n2693) );
  NAND2_X2 U4127 ( .A1(n2691), .A2(n1423), .ZN(n2692) );
  NAND2_X2 U4128 ( .A1(n2693), .A2(n2692), .ZN(n2694) );
  INV_X4 U4129 ( .A(n2694), .ZN(n2769) );
  NAND2_X2 U4130 ( .A1(a[14]), .A2(net256151), .ZN(n2702) );
  INV_X4 U4131 ( .A(n2702), .ZN(n2701) );
  NAND2_X2 U4132 ( .A1(n2771), .A2(n2703), .ZN(n2772) );
  XNOR2_X2 U4133 ( .A(n2765), .B(n2772), .ZN(n2706) );
  NAND2_X2 U4134 ( .A1(a[12]), .A2(net256119), .ZN(n2705) );
  NAND2_X2 U4135 ( .A1(n2704), .A2(n2705), .ZN(n2708) );
  INV_X4 U4136 ( .A(n2705), .ZN(n2707) );
  INV_X4 U4137 ( .A(n2710), .ZN(n2711) );
  NAND2_X2 U4138 ( .A1(a[9]), .A2(net256105), .ZN(n2712) );
  NAND3_X2 U4140 ( .A1(a[7]), .A2(n2722), .A3(net256165), .ZN(n3013) );
  NAND2_X2 U4141 ( .A1(a[7]), .A2(net256165), .ZN(n3008) );
  NAND2_X2 U4144 ( .A1(product_in[14]), .A2(net256095), .ZN(n2726) );
  NAND2_X2 U4145 ( .A1(n3983), .A2(net256183), .ZN(n2725) );
  INV_X4 U4146 ( .A(n2725), .ZN(n2728) );
  INV_X4 U4147 ( .A(n2726), .ZN(n2727) );
  INV_X4 U4148 ( .A(n2730), .ZN(n2731) );
  NAND3_X2 U4149 ( .A1(n3011), .A2(n3010), .A3(n2735), .ZN(n2736) );
  NAND3_X4 U4150 ( .A1(n2739), .A2(n2738), .A3(n2737), .ZN(n2740) );
  NAND3_X4 U4151 ( .A1(n2741), .A2(n2740), .A3(n1273), .ZN(n2938) );
  NAND2_X2 U4152 ( .A1(n2938), .A2(n2004), .ZN(n2793) );
  OAI21_X4 U4153 ( .B1(n2743), .B2(n1894), .A(n1278), .ZN(n2878) );
  NAND3_X4 U4154 ( .A1(n1916), .A2(n2949), .A3(n2948), .ZN(n2808) );
  NAND3_X2 U4155 ( .A1(net254992), .A2(n2677), .A3(n2754), .ZN(n2757) );
  NAND2_X2 U4156 ( .A1(a[12]), .A2(net256135), .ZN(n2784) );
  INV_X4 U4157 ( .A(n2784), .ZN(n2782) );
  NAND2_X2 U4158 ( .A1(n2886), .A2(n2888), .ZN(n2763) );
  OAI21_X4 U4159 ( .B1(n2764), .B2(n2763), .A(n2762), .ZN(n2781) );
  NAND2_X2 U4160 ( .A1(a[15]), .A2(net256147), .ZN(n2766) );
  INV_X4 U4161 ( .A(n2766), .ZN(n2822) );
  XNOR2_X2 U4162 ( .A(n1425), .B(n2822), .ZN(n2770) );
  INV_X4 U4163 ( .A(n2768), .ZN(n2775) );
  AOI21_X4 U4164 ( .B1(n2772), .B2(n2771), .A(n2770), .ZN(n2773) );
  OAI21_X4 U4165 ( .B1(n2775), .B2(n2774), .A(n2773), .ZN(n2821) );
  NAND2_X2 U4166 ( .A1(a[13]), .A2(net256119), .ZN(n2779) );
  XNOR2_X2 U4167 ( .A(n2781), .B(n2780), .ZN(n2783) );
  INV_X4 U4168 ( .A(n2783), .ZN(n2785) );
  NAND2_X2 U4169 ( .A1(a[10]), .A2(net256105), .ZN(n2788) );
  INV_X4 U4170 ( .A(n2788), .ZN(n2811) );
  NAND2_X2 U4171 ( .A1(n1946), .A2(n2812), .ZN(n2880) );
  NAND2_X2 U4172 ( .A1(a[9]), .A2(net256175), .ZN(n2791) );
  INV_X4 U4173 ( .A(n2791), .ZN(n2805) );
  NAND2_X2 U4174 ( .A1(n2805), .A2(n1855), .ZN(n3175) );
  XNOR2_X2 U4175 ( .A(n2793), .B(n2792), .ZN(n2795) );
  INV_X4 U4176 ( .A(n2794), .ZN(n2796) );
  NAND2_X2 U4177 ( .A1(product_in[15]), .A2(net256095), .ZN(n2798) );
  NAND2_X2 U4178 ( .A1(net256183), .A2(n4068), .ZN(n2797) );
  INV_X4 U4179 ( .A(n2797), .ZN(n2800) );
  INV_X4 U4180 ( .A(n2798), .ZN(n2799) );
  NAND2_X2 U4181 ( .A1(n2800), .A2(n2799), .ZN(n2859) );
  XNOR2_X2 U4182 ( .A(n2802), .B(n1854), .ZN(product_out[15]) );
  NAND2_X2 U4183 ( .A1(product_in[16]), .A2(net256095), .ZN(n2863) );
  NAND2_X2 U4184 ( .A1(n2803), .A2(n1922), .ZN(n2804) );
  AOI21_X4 U4185 ( .B1(n2805), .B2(n1957), .A(n2940), .ZN(n2806) );
  NAND2_X2 U4186 ( .A1(n2950), .A2(n2881), .ZN(n2814) );
  NAND2_X2 U4187 ( .A1(a[11]), .A2(net256105), .ZN(net254858) );
  NAND2_X2 U4188 ( .A1(a[14]), .A2(net256117), .ZN(n2828) );
  INV_X4 U4189 ( .A(n2828), .ZN(n2825) );
  NAND2_X2 U4190 ( .A1(a[15]), .A2(n1460), .ZN(n2817) );
  NAND2_X2 U4191 ( .A1(a[16]), .A2(net256147), .ZN(n2818) );
  NAND2_X2 U4192 ( .A1(n2817), .A2(n2818), .ZN(n2820) );
  INV_X4 U4193 ( .A(n2818), .ZN(n2819) );
  NAND2_X2 U4194 ( .A1(n2820), .A2(n2900), .ZN(n2901) );
  INV_X4 U4195 ( .A(n2901), .ZN(n2824) );
  NOR2_X4 U4196 ( .A1(n2899), .A2(n1407), .ZN(n2823) );
  XNOR2_X2 U4197 ( .A(n2824), .B(n2823), .ZN(n2826) );
  INV_X4 U4198 ( .A(n2889), .ZN(n2831) );
  NAND3_X2 U4199 ( .A1(n2888), .A2(n2832), .A3(n2890), .ZN(n2836) );
  NAND3_X4 U4200 ( .A1(n2836), .A2(n1814), .A3(n2892), .ZN(n3038) );
  XNOR2_X2 U4201 ( .A(n3038), .B(n3037), .ZN(n2837) );
  NAND2_X2 U4202 ( .A1(a[12]), .A2(net256125), .ZN(net254871) );
  NAND2_X2 U4203 ( .A1(a[10]), .A2(net256175), .ZN(n2841) );
  INV_X4 U4204 ( .A(n2841), .ZN(n2844) );
  OAI21_X4 U4205 ( .B1(n2847), .B2(n1269), .A(n3015), .ZN(n2848) );
  NAND3_X4 U4206 ( .A1(n2857), .A2(n2856), .A3(n2855), .ZN(n2860) );
  INV_X4 U4207 ( .A(n2859), .ZN(n2862) );
  OAI21_X4 U4208 ( .B1(n2861), .B2(n2862), .A(n1839), .ZN(n3091) );
  INV_X4 U4209 ( .A(n2863), .ZN(n2865) );
  NAND2_X2 U4210 ( .A1(n2865), .A2(n2864), .ZN(n3092) );
  INV_X4 U4211 ( .A(n2866), .ZN(n2869) );
  NAND2_X2 U4212 ( .A1(a[10]), .A2(net256165), .ZN(n2925) );
  INV_X4 U4213 ( .A(n2925), .ZN(n2924) );
  OAI21_X4 U4214 ( .B1(n2874), .B2(n2873), .A(n3024), .ZN(n2877) );
  NAND2_X2 U4215 ( .A1(n2875), .A2(n1848), .ZN(n2876) );
  NOR2_X4 U4216 ( .A1(n2879), .A2(n1904), .ZN(n2884) );
  OAI21_X4 U4217 ( .B1(n2883), .B2(n2884), .A(n2882), .ZN(n2919) );
  INV_X4 U4218 ( .A(a[14]), .ZN(n2913) );
  NOR2_X4 U4219 ( .A1(n3037), .A2(n2887), .ZN(n2891) );
  NAND4_X2 U4220 ( .A1(n2891), .A2(n2888), .A3(n2889), .A4(n2890), .ZN(n2898)
         );
  INV_X4 U4221 ( .A(n2892), .ZN(n2896) );
  INV_X4 U4222 ( .A(n3037), .ZN(n2894) );
  OAI21_X4 U4223 ( .B1(n2896), .B2(n2895), .A(n2894), .ZN(n2897) );
  NAND3_X4 U4224 ( .A1(n2898), .A2(n2897), .A3(n1928), .ZN(n2964) );
  NOR2_X4 U4225 ( .A1(n2899), .A2(n1407), .ZN(n2902) );
  OAI21_X4 U4226 ( .B1(n2902), .B2(n2901), .A(n2900), .ZN(n3049) );
  NAND2_X2 U4227 ( .A1(a[17]), .A2(net256151), .ZN(n2903) );
  INV_X4 U4228 ( .A(n2903), .ZN(n2966) );
  XNOR2_X2 U4229 ( .A(n1426), .B(n2966), .ZN(n3048) );
  INV_X4 U4230 ( .A(n3048), .ZN(n2905) );
  NAND2_X2 U4231 ( .A1(n2905), .A2(n3049), .ZN(n2967) );
  NAND2_X2 U4232 ( .A1(a[15]), .A2(net256117), .ZN(n2908) );
  INV_X4 U4233 ( .A(n2908), .ZN(n2906) );
  NAND3_X2 U4234 ( .A1(n2907), .A2(n2967), .A3(n2906), .ZN(n3040) );
  INV_X4 U4235 ( .A(n2907), .ZN(n2909) );
  OAI21_X4 U4236 ( .B1(n2910), .B2(n2909), .A(n2908), .ZN(n2911) );
  XNOR2_X2 U4237 ( .A(n2964), .B(n1955), .ZN(n2914) );
  INV_X4 U4238 ( .A(n2914), .ZN(n2912) );
  OAI21_X4 U4239 ( .B1(net256139), .B2(n2913), .A(n2912), .ZN(n3196) );
  INV_X4 U4240 ( .A(n3196), .ZN(n3143) );
  NAND2_X2 U4241 ( .A1(n1866), .A2(n1111), .ZN(n2916) );
  NOR2_X4 U4242 ( .A1(n1139), .A2(net256095), .ZN(n2932) );
  NAND2_X2 U4243 ( .A1(product_in[17]), .A2(net256095), .ZN(n2928) );
  NAND2_X2 U4244 ( .A1(n2927), .A2(n2928), .ZN(n2931) );
  INV_X4 U4245 ( .A(n2928), .ZN(n2930) );
  NAND2_X2 U4246 ( .A1(n2930), .A2(n2929), .ZN(n3094) );
  OAI21_X4 U4247 ( .B1(n2932), .B2(n2931), .A(n3094), .ZN(n3098) );
  INV_X4 U4248 ( .A(n2935), .ZN(n3005) );
  NAND2_X2 U4249 ( .A1(n2937), .A2(n2936), .ZN(n3688) );
  INV_X4 U4250 ( .A(n3688), .ZN(n2992) );
  NAND3_X2 U4251 ( .A1(n2949), .A2(n2948), .A3(n2747), .ZN(n2951) );
  AOI21_X4 U4252 ( .B1(n2951), .B2(n2952), .A(n2950), .ZN(n2953) );
  NAND2_X2 U4253 ( .A1(a[13]), .A2(net253103), .ZN(net254634) );
  NAND2_X2 U4254 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  NAND2_X2 U4255 ( .A1(a[14]), .A2(net256125), .ZN(n2982) );
  INV_X4 U4256 ( .A(n2982), .ZN(n2981) );
  OAI21_X4 U4257 ( .B1(n2965), .B2(n1955), .A(n3040), .ZN(n2975) );
  NAND2_X2 U4258 ( .A1(n1426), .A2(n2966), .ZN(n3046) );
  NAND2_X2 U4259 ( .A1(a[18]), .A2(net256147), .ZN(n2968) );
  INV_X4 U4260 ( .A(n2968), .ZN(n2970) );
  INV_X4 U4261 ( .A(a[17]), .ZN(net254656) );
  XNOR2_X2 U4262 ( .A(n2971), .B(n3047), .ZN(n2972) );
  NAND2_X2 U4263 ( .A1(a[16]), .A2(net256117), .ZN(n2973) );
  NAND2_X2 U4264 ( .A1(n2973), .A2(n1837), .ZN(n2974) );
  XNOR2_X2 U4265 ( .A(n2975), .B(n3207), .ZN(n2978) );
  NAND2_X2 U4266 ( .A1(a[15]), .A2(net256135), .ZN(n2977) );
  INV_X4 U4267 ( .A(n2977), .ZN(n2979) );
  INV_X4 U4268 ( .A(n2985), .ZN(n2986) );
  XNOR2_X2 U4269 ( .A(n2988), .B(n2987), .ZN(n3108) );
  NAND2_X2 U4270 ( .A1(n2994), .A2(n3688), .ZN(n3001) );
  NAND2_X2 U4271 ( .A1(n3692), .A2(n1922), .ZN(n2999) );
  NAND2_X2 U4272 ( .A1(product_in[19]), .A2(net256095), .ZN(n3006) );
  NAND3_X2 U4273 ( .A1(n3011), .A2(n3010), .A3(n3009), .ZN(n3014) );
  NAND3_X2 U4274 ( .A1(n1267), .A2(n1778), .A3(n3021), .ZN(n3022) );
  OAI21_X4 U4275 ( .B1(n3028), .B2(n1996), .A(n4104), .ZN(n3161) );
  NAND2_X2 U4276 ( .A1(net254671), .A2(net257880), .ZN(n3029) );
  OAI21_X4 U4277 ( .B1(n3032), .B2(net254562), .A(n1449), .ZN(n3146) );
  NOR2_X4 U4278 ( .A1(n3042), .A2(n3037), .ZN(n3039) );
  NOR2_X4 U4279 ( .A1(n3043), .A2(n3119), .ZN(n3044) );
  NAND2_X2 U4280 ( .A1(n3046), .A2(n3045), .ZN(n3216) );
  INV_X4 U4281 ( .A(n3216), .ZN(n3051) );
  NAND2_X2 U4282 ( .A1(a[19]), .A2(net256147), .ZN(n3052) );
  INV_X4 U4283 ( .A(n3052), .ZN(n3125) );
  XNOR2_X2 U4284 ( .A(n1427), .B(n3125), .ZN(n3054) );
  INV_X4 U4285 ( .A(n3054), .ZN(n3221) );
  INV_X4 U4286 ( .A(n3126), .ZN(n3059) );
  INV_X4 U4287 ( .A(n3056), .ZN(n3058) );
  NAND2_X2 U4288 ( .A1(a[17]), .A2(net256117), .ZN(n3057) );
  OAI21_X4 U4289 ( .B1(n3059), .B2(n3058), .A(n3057), .ZN(n3060) );
  XNOR2_X2 U4290 ( .A(n3061), .B(n1614), .ZN(n3192) );
  NAND2_X2 U4291 ( .A1(a[16]), .A2(net256135), .ZN(n3191) );
  INV_X4 U4292 ( .A(n3191), .ZN(n3063) );
  NAND2_X2 U4293 ( .A1(n3138), .A2(n3198), .ZN(n3064) );
  XNOR2_X2 U4294 ( .A(n3065), .B(n3064), .ZN(n3068) );
  NAND2_X2 U4295 ( .A1(a[15]), .A2(net256125), .ZN(n3067) );
  INV_X4 U4296 ( .A(n3067), .ZN(n3069) );
  NAND2_X2 U4297 ( .A1(a[13]), .A2(net256175), .ZN(n3074) );
  INV_X4 U4298 ( .A(n3074), .ZN(n3077) );
  XNOR2_X2 U4300 ( .A(n1134), .B(n3078), .ZN(n3082) );
  INV_X4 U4301 ( .A(n1433), .ZN(n3080) );
  NAND2_X2 U4302 ( .A1(a[12]), .A2(net256165), .ZN(n3081) );
  INV_X4 U4303 ( .A(n3081), .ZN(n3083) );
  XNOR2_X2 U4305 ( .A(n3085), .B(n3084), .ZN(n3086) );
  AOI21_X2 U4306 ( .B1(net256183), .B2(n3759), .A(n3087), .ZN(n3088) );
  OAI21_X4 U4307 ( .B1(n3761), .B2(net256095), .A(n3088), .ZN(n3089) );
  INV_X4 U4308 ( .A(n3094), .ZN(n3096) );
  NOR2_X4 U4309 ( .A1(n3096), .A2(n3095), .ZN(n3097) );
  OAI21_X4 U4310 ( .B1(n3099), .B2(n3098), .A(n3097), .ZN(n3496) );
  NAND2_X2 U4311 ( .A1(n3103), .A2(n3102), .ZN(n3335) );
  INV_X4 U4312 ( .A(n3105), .ZN(n3106) );
  OAI21_X4 U4313 ( .B1(n3111), .B2(n1852), .A(n1799), .ZN(n3525) );
  INV_X4 U4314 ( .A(n3248), .ZN(n3244) );
  NAND2_X2 U4315 ( .A1(n3114), .A2(n3115), .ZN(n3153) );
  NAND2_X2 U4316 ( .A1(a[16]), .A2(net256125), .ZN(n3152) );
  INV_X4 U4317 ( .A(n3152), .ZN(n3243) );
  INV_X4 U4318 ( .A(n3208), .ZN(n3122) );
  NAND2_X2 U4319 ( .A1(n3206), .A2(n3205), .ZN(n3118) );
  INV_X4 U4320 ( .A(n3118), .ZN(n3210) );
  INV_X4 U4321 ( .A(n3119), .ZN(n3121) );
  NAND3_X2 U4322 ( .A1(n3209), .A2(n3123), .A3(n3122), .ZN(n3124) );
  NAND2_X2 U4323 ( .A1(a[18]), .A2(net256117), .ZN(n3133) );
  NAND2_X2 U4324 ( .A1(n1427), .A2(n3125), .ZN(n3215) );
  NAND2_X2 U4325 ( .A1(n3126), .A2(n3215), .ZN(n3131) );
  NAND2_X2 U4326 ( .A1(a[19]), .A2(n1460), .ZN(n3127) );
  NAND2_X2 U4327 ( .A1(a[20]), .A2(net256147), .ZN(n3128) );
  NAND2_X2 U4328 ( .A1(n3127), .A2(n3128), .ZN(n3130) );
  INV_X4 U4329 ( .A(n3128), .ZN(n3129) );
  NAND2_X2 U4330 ( .A1(n3130), .A2(n3297), .ZN(n3219) );
  XNOR2_X2 U4331 ( .A(n3131), .B(n3219), .ZN(n3134) );
  INV_X4 U4332 ( .A(n3134), .ZN(n3132) );
  NAND2_X2 U4333 ( .A1(n3133), .A2(n3132), .ZN(n3135) );
  NAND3_X2 U4334 ( .A1(a[18]), .A2(n3134), .A3(net256117), .ZN(n3352) );
  NAND3_X4 U4335 ( .A1(n3136), .A2(a[17]), .A3(net256135), .ZN(n3291) );
  NAND2_X2 U4336 ( .A1(a[17]), .A2(net256135), .ZN(n3137) );
  OAI21_X4 U4337 ( .B1(n3145), .B2(n1949), .A(n3144), .ZN(n3147) );
  OAI21_X4 U4338 ( .B1(n3148), .B2(n3147), .A(n1437), .ZN(n3149) );
  XNOR2_X2 U4339 ( .A(n3149), .B(n3150), .ZN(n3242) );
  INV_X4 U4340 ( .A(n3242), .ZN(n3151) );
  NAND2_X2 U4341 ( .A1(n3249), .A2(net254291), .ZN(n3456) );
  NAND2_X2 U4342 ( .A1(a[15]), .A2(net253103), .ZN(net254415) );
  NAND2_X2 U4343 ( .A1(net254415), .A2(net254414), .ZN(net254235) );
  NAND2_X2 U4344 ( .A1(a[14]), .A2(net256175), .ZN(n3156) );
  INV_X4 U4345 ( .A(n3156), .ZN(n3159) );
  NAND2_X2 U4346 ( .A1(a[13]), .A2(net256165), .ZN(n3165) );
  INV_X4 U4347 ( .A(n3165), .ZN(n3167) );
  OAI22_X2 U4348 ( .A1(n3512), .A2(net254390), .B1(n3169), .B2(net256184), 
        .ZN(n3266) );
  INV_X4 U4349 ( .A(n3266), .ZN(n3170) );
  OAI21_X4 U4350 ( .B1(n1846), .B2(net256095), .A(n3170), .ZN(n3171) );
  NAND2_X2 U4351 ( .A1(product_in[20]), .A2(net256095), .ZN(n3265) );
  NAND2_X2 U4352 ( .A1(product_in[21]), .A2(net256095), .ZN(n3262) );
  INV_X4 U4353 ( .A(n3262), .ZN(n3260) );
  AOI21_X4 U4354 ( .B1(n3178), .B2(n3180), .A(n3177), .ZN(n3183) );
  NAND3_X2 U4355 ( .A1(n3180), .A2(n3181), .A3(n1301), .ZN(n3182) );
  NAND3_X2 U4356 ( .A1(n3187), .A2(n1825), .A3(n3186), .ZN(n3188) );
  INV_X4 U4357 ( .A(n3193), .ZN(n3194) );
  NAND3_X4 U4358 ( .A1(n3199), .A2(n3200), .A3(n3198), .ZN(n3201) );
  NAND3_X4 U4359 ( .A1(n3201), .A2(n3202), .A3(n3203), .ZN(n3289) );
  INV_X4 U4360 ( .A(n3204), .ZN(n3214) );
  OAI211_X2 U4361 ( .C1(n1614), .C2(n3207), .A(n3206), .B(n3205), .ZN(n3213)
         );
  INV_X4 U4362 ( .A(n3209), .ZN(n3211) );
  NAND3_X4 U4363 ( .A1(n3214), .A2(n3212), .A3(n3213), .ZN(n3353) );
  INV_X4 U4364 ( .A(n3215), .ZN(n3222) );
  NOR2_X4 U4365 ( .A1(n3222), .A2(n3216), .ZN(n3218) );
  INV_X4 U4366 ( .A(n3304), .ZN(n3223) );
  INV_X4 U4367 ( .A(n3219), .ZN(n3220) );
  OAI21_X4 U4368 ( .B1(n3222), .B2(n3221), .A(n3220), .ZN(n3302) );
  OAI21_X4 U4369 ( .B1(n3223), .B2(n3302), .A(n3297), .ZN(n3226) );
  NAND2_X2 U4370 ( .A1(a[20]), .A2(n1460), .ZN(n3298) );
  INV_X4 U4371 ( .A(n3298), .ZN(n3225) );
  NAND2_X2 U4372 ( .A1(a[21]), .A2(net256147), .ZN(n3299) );
  INV_X4 U4373 ( .A(n3299), .ZN(n3224) );
  XNOR2_X2 U4374 ( .A(n3225), .B(n3224), .ZN(n3227) );
  INV_X4 U4375 ( .A(n3227), .ZN(n3305) );
  NAND2_X2 U4376 ( .A1(n3226), .A2(n3305), .ZN(n3233) );
  INV_X4 U4377 ( .A(n3233), .ZN(n3231) );
  INV_X4 U4378 ( .A(n3226), .ZN(n3228) );
  NAND2_X2 U4379 ( .A1(n3228), .A2(n3227), .ZN(n3232) );
  INV_X4 U4380 ( .A(n3232), .ZN(n3230) );
  NAND2_X2 U4381 ( .A1(a[19]), .A2(net256117), .ZN(n3229) );
  OAI21_X4 U4382 ( .B1(n3231), .B2(n3230), .A(n3229), .ZN(n3234) );
  NAND4_X2 U4383 ( .A1(a[19]), .A2(n3233), .A3(n3232), .A4(net256117), .ZN(
        n3430) );
  XNOR2_X2 U4384 ( .A(n1293), .B(n3427), .ZN(n3238) );
  NAND2_X2 U4385 ( .A1(a[18]), .A2(net256135), .ZN(n3237) );
  INV_X4 U4386 ( .A(n3237), .ZN(n3239) );
  NAND2_X2 U4387 ( .A1(n3239), .A2(n3238), .ZN(n3290) );
  XNOR2_X2 U4388 ( .A(n3241), .B(n3240), .ZN(n3250) );
  NAND2_X2 U4389 ( .A1(a[16]), .A2(net256105), .ZN(net254285) );
  INV_X4 U4390 ( .A(n3455), .ZN(n3246) );
  NAND3_X4 U4391 ( .A1(n1317), .A2(n1668), .A3(n3453), .ZN(net254298) );
  OAI21_X4 U4392 ( .B1(net254293), .B2(n3248), .A(n3324), .ZN(net254001) );
  NAND2_X2 U4393 ( .A1(n1404), .A2(n4086), .ZN(n3348) );
  XNOR2_X2 U4394 ( .A(net258069), .B(net254192), .ZN(net254242) );
  NAND2_X2 U4395 ( .A1(a[15]), .A2(net256173), .ZN(n3251) );
  INV_X4 U4396 ( .A(n3251), .ZN(n3277) );
  XNOR2_X2 U4397 ( .A(n3344), .B(n3388), .ZN(n3253) );
  NAND2_X2 U4398 ( .A1(a[14]), .A2(net256165), .ZN(n3343) );
  INV_X4 U4399 ( .A(n3343), .ZN(n3255) );
  NAND2_X2 U4400 ( .A1(n3256), .A2(n1769), .ZN(n3274) );
  INV_X4 U4401 ( .A(n3265), .ZN(n3267) );
  NAND2_X2 U4402 ( .A1(n3267), .A2(n3266), .ZN(n3337) );
  NOR2_X4 U4403 ( .A1(n3272), .A2(n1892), .ZN(n3276) );
  NAND2_X2 U4404 ( .A1(n3274), .A2(n1769), .ZN(n3275) );
  OAI21_X4 U4405 ( .B1(n3276), .B2(n1971), .A(n3275), .ZN(n3329) );
  NAND3_X4 U4406 ( .A1(n3280), .A2(n1340), .A3(n3282), .ZN(n3283) );
  NAND2_X2 U4408 ( .A1(a[18]), .A2(net256125), .ZN(n3458) );
  INV_X4 U4409 ( .A(n3458), .ZN(n3320) );
  NAND3_X4 U4410 ( .A1(n3289), .A2(n3290), .A3(n3291), .ZN(n3437) );
  NAND2_X2 U4411 ( .A1(n3437), .A2(n1844), .ZN(n3292) );
  NAND2_X2 U4412 ( .A1(a[20]), .A2(net256117), .ZN(n3309) );
  NAND2_X2 U4413 ( .A1(a[21]), .A2(n1460), .ZN(n3293) );
  NAND2_X2 U4414 ( .A1(a[22]), .A2(net256147), .ZN(n3294) );
  NAND2_X2 U4415 ( .A1(n3293), .A2(n3294), .ZN(n3296) );
  INV_X4 U4416 ( .A(n3294), .ZN(n3295) );
  NAND2_X2 U4417 ( .A1(n3296), .A2(n3359), .ZN(n3360) );
  INV_X4 U4418 ( .A(n3297), .ZN(n3301) );
  NOR2_X4 U4419 ( .A1(n3299), .A2(n3298), .ZN(n3300) );
  NOR2_X4 U4420 ( .A1(n3301), .A2(n3300), .ZN(n3307) );
  INV_X4 U4421 ( .A(n3302), .ZN(n3303) );
  NAND3_X2 U4422 ( .A1(n3305), .A2(n3304), .A3(n3303), .ZN(n3306) );
  XNOR2_X2 U4423 ( .A(n3360), .B(n3358), .ZN(n3310) );
  INV_X4 U4424 ( .A(n3310), .ZN(n3308) );
  NAND2_X2 U4425 ( .A1(n3309), .A2(n3308), .ZN(n3311) );
  NAND3_X2 U4426 ( .A1(a[20]), .A2(n3310), .A3(net256117), .ZN(n3429) );
  NAND2_X2 U4427 ( .A1(n3427), .A2(n3430), .ZN(n3313) );
  XNOR2_X2 U4428 ( .A(n3431), .B(n3314), .ZN(n3316) );
  NAND2_X2 U4429 ( .A1(a[19]), .A2(net256135), .ZN(n3315) );
  INV_X4 U4430 ( .A(n3315), .ZN(n3318) );
  XNOR2_X2 U4431 ( .A(n3441), .B(n3321), .ZN(n3319) );
  XNOR2_X2 U4432 ( .A(n3322), .B(n3321), .ZN(n3459) );
  INV_X4 U4433 ( .A(n3549), .ZN(n3347) );
  NAND2_X2 U4434 ( .A1(n3323), .A2(n1292), .ZN(n3325) );
  XNOR2_X2 U4435 ( .A(net254179), .B(n3629), .ZN(n3533) );
  NAND2_X2 U4436 ( .A1(a[15]), .A2(net256165), .ZN(n3532) );
  INV_X4 U4437 ( .A(n3532), .ZN(n3327) );
  NAND2_X2 U4438 ( .A1(n3536), .A2(n3535), .ZN(n3328) );
  XNOR2_X2 U4439 ( .A(n3329), .B(n3328), .ZN(n3986) );
  NAND2_X2 U4440 ( .A1(n3983), .A2(n1922), .ZN(n3330) );
  OAI21_X4 U4441 ( .B1(n4111), .B2(net256184), .A(n3330), .ZN(n3341) );
  INV_X4 U4442 ( .A(n3341), .ZN(n3332) );
  INV_X4 U4443 ( .A(n3340), .ZN(n3333) );
  NAND2_X2 U4444 ( .A1(n3333), .A2(n3341), .ZN(n3493) );
  XNOR2_X2 U4445 ( .A(n3388), .B(n3343), .ZN(n3345) );
  OAI221_X2 U4446 ( .B1(n3474), .B2(n1436), .C1(n3474), .C2(n1849), .A(n1992), 
        .ZN(n3396) );
  INV_X4 U4447 ( .A(net257068), .ZN(net254058) );
  INV_X4 U4448 ( .A(n3395), .ZN(n3472) );
  NAND2_X2 U4449 ( .A1(a[17]), .A2(net256175), .ZN(net254085) );
  INV_X4 U4450 ( .A(n3547), .ZN(n3349) );
  NOR2_X4 U4451 ( .A1(n3428), .A2(n3427), .ZN(n3356) );
  OAI21_X4 U4452 ( .B1(n3356), .B2(n3355), .A(n3354), .ZN(n3372) );
  NAND2_X2 U4453 ( .A1(a[23]), .A2(net256151), .ZN(n3357) );
  INV_X4 U4454 ( .A(n3357), .ZN(n3415) );
  XNOR2_X2 U4455 ( .A(n1428), .B(n3415), .ZN(n3364) );
  INV_X4 U4456 ( .A(n3364), .ZN(n3362) );
  INV_X4 U4457 ( .A(n3358), .ZN(n3361) );
  OAI21_X4 U4458 ( .B1(n3361), .B2(n3360), .A(n3359), .ZN(n3363) );
  NAND2_X2 U4460 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  NAND2_X2 U4461 ( .A1(n3416), .A2(n3366), .ZN(n3369) );
  INV_X4 U4462 ( .A(n3369), .ZN(n3368) );
  NAND2_X2 U4463 ( .A1(a[21]), .A2(net256117), .ZN(n3370) );
  INV_X4 U4464 ( .A(n3370), .ZN(n3367) );
  NAND2_X2 U4465 ( .A1(n3368), .A2(n3367), .ZN(n3568) );
  NAND2_X2 U4466 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  NAND2_X2 U4467 ( .A1(n3568), .A2(n3371), .ZN(n3432) );
  XNOR2_X2 U4468 ( .A(n3372), .B(n3432), .ZN(n3374) );
  NAND2_X2 U4469 ( .A1(a[20]), .A2(net256135), .ZN(n3373) );
  INV_X4 U4470 ( .A(n3373), .ZN(n3376) );
  INV_X4 U4471 ( .A(n3374), .ZN(n3375) );
  NAND3_X4 U4472 ( .A1(n3437), .A2(n3442), .A3(n1844), .ZN(n3377) );
  XNOR2_X2 U4473 ( .A(n3379), .B(n3378), .ZN(n3381) );
  NAND2_X2 U4474 ( .A1(a[19]), .A2(net256125), .ZN(n3380) );
  INV_X4 U4475 ( .A(n3380), .ZN(n3382) );
  XNOR2_X2 U4476 ( .A(net254082), .B(net254083), .ZN(n3391) );
  NOR2_X4 U4477 ( .A1(n3630), .A2(n3391), .ZN(n3392) );
  INV_X4 U4478 ( .A(n3392), .ZN(n3393) );
  NOR2_X4 U4479 ( .A1(n1189), .A2(net256095), .ZN(n3403) );
  OAI22_X2 U4480 ( .A1(n3397), .A2(n3512), .B1(n1129), .B2(net256184), .ZN(
        n3400) );
  INV_X4 U4481 ( .A(n3400), .ZN(n3398) );
  NAND2_X2 U4482 ( .A1(product_in[23]), .A2(net256095), .ZN(n3399) );
  NAND2_X2 U4483 ( .A1(n3398), .A2(n3399), .ZN(n3402) );
  INV_X4 U4484 ( .A(n3399), .ZN(n3401) );
  NAND2_X2 U4485 ( .A1(n3401), .A2(n3400), .ZN(n3784) );
  OAI21_X4 U4486 ( .B1(n3403), .B2(n3402), .A(n3784), .ZN(n3505) );
  NAND2_X2 U4487 ( .A1(n1922), .A2(n3407), .ZN(n3408) );
  NAND2_X2 U4488 ( .A1(n3786), .A2(net256095), .ZN(n3481) );
  NAND2_X2 U4489 ( .A1(product_in[24]), .A2(net256095), .ZN(n3785) );
  NAND2_X2 U4490 ( .A1(n3481), .A2(n3785), .ZN(n3486) );
  NAND2_X2 U4491 ( .A1(a[17]), .A2(net256165), .ZN(n3469) );
  INV_X4 U4492 ( .A(n3469), .ZN(n3468) );
  NAND2_X2 U4493 ( .A1(a[19]), .A2(net256105), .ZN(n3608) );
  NAND2_X2 U4494 ( .A1(a[22]), .A2(net256117), .ZN(n3424) );
  NAND2_X2 U4495 ( .A1(n1428), .A2(n3415), .ZN(n3417) );
  NAND2_X2 U4496 ( .A1(a[23]), .A2(net256143), .ZN(n3419) );
  NAND2_X2 U4497 ( .A1(a[24]), .A2(net256147), .ZN(n3420) );
  NAND2_X2 U4498 ( .A1(n3419), .A2(n3420), .ZN(n3422) );
  INV_X4 U4499 ( .A(n3420), .ZN(n3421) );
  NAND2_X2 U4500 ( .A1(n3422), .A2(n3574), .ZN(n3575) );
  XNOR2_X2 U4501 ( .A(n3576), .B(n3423), .ZN(n3425) );
  NAND2_X2 U4502 ( .A1(n3424), .A2(n1913), .ZN(n3426) );
  NAND3_X2 U4503 ( .A1(a[22]), .A2(n3425), .A3(net256117), .ZN(n3569) );
  NAND2_X2 U4504 ( .A1(a[21]), .A2(net256135), .ZN(n3557) );
  XNOR2_X2 U4505 ( .A(n3570), .B(n3557), .ZN(n3436) );
  INV_X4 U4506 ( .A(n3432), .ZN(n3433) );
  OAI21_X4 U4507 ( .B1(n3435), .B2(n3434), .A(n3433), .ZN(n3567) );
  XNOR2_X2 U4508 ( .A(n3436), .B(n3558), .ZN(n3638) );
  INV_X4 U4509 ( .A(n3638), .ZN(n3443) );
  NOR2_X4 U4510 ( .A1(n3634), .A2(n3443), .ZN(n3440) );
  NAND3_X2 U4511 ( .A1(n3636), .A2(n1903), .A3(n3637), .ZN(n3439) );
  NAND3_X4 U4512 ( .A1(n1908), .A2(n1915), .A3(n3441), .ZN(n3447) );
  NOR2_X4 U4513 ( .A1(n3451), .A2(n3444), .ZN(n3445) );
  NAND2_X2 U4514 ( .A1(a[20]), .A2(net256125), .ZN(n3448) );
  INV_X4 U4515 ( .A(n3448), .ZN(n3449) );
  INV_X4 U4516 ( .A(n3454), .ZN(n3457) );
  INV_X4 U4517 ( .A(n3473), .ZN(n3477) );
  NAND2_X2 U4518 ( .A1(n3785), .A2(n3507), .ZN(n3482) );
  INV_X4 U4519 ( .A(n3481), .ZN(n3480) );
  AOI22_X2 U4520 ( .A1(n3482), .A2(n3481), .B1(n3480), .B2(n3785), .ZN(n3483)
         );
  INV_X4 U4521 ( .A(n3485), .ZN(n3489) );
  INV_X4 U4522 ( .A(n3543), .ZN(n3487) );
  NOR2_X4 U4523 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  INV_X4 U4524 ( .A(n3493), .ZN(n3781) );
  NAND3_X2 U4525 ( .A1(n1440), .A2(n3503), .A3(n3501), .ZN(n3504) );
  NAND2_X2 U4526 ( .A1(net253179), .A2(n3784), .ZN(n3509) );
  XNOR2_X2 U4527 ( .A(net253936), .B(n3509), .ZN(product_out[24]) );
  INV_X4 U4528 ( .A(n3785), .ZN(n3508) );
  INV_X4 U4529 ( .A(net253187), .ZN(net253535) );
  NAND2_X2 U4530 ( .A1(net253067), .A2(n3510), .ZN(n3511) );
  NAND2_X2 U4531 ( .A1(product_in[25]), .A2(net256095), .ZN(n3515) );
  NAND2_X2 U4532 ( .A1(n3514), .A2(n3515), .ZN(net253183) );
  INV_X4 U4533 ( .A(n3515), .ZN(n3517) );
  NAND2_X2 U4534 ( .A1(net253183), .A2(n3790), .ZN(n3763) );
  XNOR2_X2 U4535 ( .A(n3518), .B(n3763), .ZN(n3620) );
  INV_X4 U4536 ( .A(n1842), .ZN(n3522) );
  XNOR2_X2 U4537 ( .A(n3528), .B(n3527), .ZN(n3529) );
  NOR2_X4 U4538 ( .A1(n1879), .A2(n3539), .ZN(n3540) );
  NAND3_X4 U4539 ( .A1(n3542), .A2(n3540), .A3(n3541), .ZN(n3855) );
  INV_X4 U4540 ( .A(n3616), .ZN(n3618) );
  NAND2_X2 U4541 ( .A1(a[20]), .A2(net256105), .ZN(n3598) );
  INV_X4 U4542 ( .A(n3598), .ZN(n3686) );
  AOI211_X4 U4543 ( .C1(n3604), .C2(n3552), .A(n3682), .B(n3677), .ZN(n3553)
         );
  OAI21_X4 U4544 ( .B1(n3555), .B2(n3554), .A(n3553), .ZN(n3596) );
  NAND2_X2 U4545 ( .A1(a[21]), .A2(net256125), .ZN(n3592) );
  INV_X4 U4546 ( .A(n3592), .ZN(n3591) );
  NAND2_X2 U4547 ( .A1(n3636), .A2(n1903), .ZN(n3562) );
  INV_X4 U4548 ( .A(n3557), .ZN(n3560) );
  XNOR2_X2 U4549 ( .A(n3558), .B(n3570), .ZN(n3559) );
  INV_X4 U4550 ( .A(n3637), .ZN(n3561) );
  NOR3_X4 U4551 ( .A1(n3562), .A2(n3564), .A3(n3561), .ZN(n3566) );
  NAND2_X2 U4552 ( .A1(n1830), .A2(n3568), .ZN(n3649) );
  NAND2_X2 U4553 ( .A1(n3570), .A2(n1830), .ZN(n3647) );
  OAI21_X4 U4554 ( .B1(n3650), .B2(n3649), .A(n3647), .ZN(n3584) );
  NAND2_X2 U4555 ( .A1(a[23]), .A2(net256117), .ZN(n3580) );
  INV_X4 U4556 ( .A(n3571), .ZN(n3659) );
  NAND2_X2 U4557 ( .A1(a[25]), .A2(net256147), .ZN(n3572) );
  INV_X4 U4558 ( .A(n3572), .ZN(n3658) );
  XNOR2_X2 U4559 ( .A(n3659), .B(n3658), .ZN(n3573) );
  INV_X4 U4560 ( .A(n3573), .ZN(n3578) );
  OAI21_X4 U4561 ( .B1(n3576), .B2(n3575), .A(n3574), .ZN(n3577) );
  NAND2_X2 U4563 ( .A1(n3580), .A2(n3579), .ZN(n3583) );
  INV_X4 U4564 ( .A(n3579), .ZN(n3582) );
  INV_X4 U4565 ( .A(n3580), .ZN(n3581) );
  NAND2_X2 U4566 ( .A1(n3582), .A2(n3581), .ZN(n3651) );
  XNOR2_X2 U4567 ( .A(n3584), .B(n3646), .ZN(n3586) );
  NAND3_X4 U4568 ( .A1(a[22]), .A2(n1901), .A3(net256135), .ZN(n3645) );
  INV_X4 U4569 ( .A(n3645), .ZN(n3717) );
  NAND2_X2 U4570 ( .A1(a[22]), .A2(net256135), .ZN(n3585) );
  NOR2_X4 U4571 ( .A1(n3717), .A2(n3639), .ZN(n3588) );
  XNOR2_X2 U4572 ( .A(n3589), .B(n3588), .ZN(n3593) );
  INV_X4 U4573 ( .A(n1797), .ZN(n3590) );
  NOR2_X4 U4574 ( .A1(n1337), .A2(n3598), .ZN(n3599) );
  XNOR2_X2 U4575 ( .A(n3600), .B(n3599), .ZN(n3601) );
  NAND2_X2 U4576 ( .A1(a[19]), .A2(net256173), .ZN(net253780) );
  XNOR2_X2 U4577 ( .A(n3607), .B(n3678), .ZN(n3609) );
  OAI21_X4 U4578 ( .B1(net253816), .B2(net253815), .A(n3610), .ZN(n3613) );
  NOR2_X4 U4579 ( .A1(net257838), .A2(net253780), .ZN(n3611) );
  NAND3_X2 U4580 ( .A1(net253448), .A2(net253647), .A3(n3614), .ZN(n3621) );
  NAND2_X2 U4582 ( .A1(n3620), .A2(n3619), .ZN(product_out[25]) );
  INV_X4 U4583 ( .A(net253780), .ZN(net253762) );
  XNOR2_X2 U4584 ( .A(net253770), .B(n3631), .ZN(n3632) );
  OAI21_X4 U4585 ( .B1(n1977), .B2(n3702), .A(n3701), .ZN(n3857) );
  NOR2_X4 U4586 ( .A1(n3708), .A2(n3857), .ZN(n3687) );
  NAND2_X2 U4587 ( .A1(a[20]), .A2(net256173), .ZN(net253643) );
  NAND2_X2 U4588 ( .A1(a[21]), .A2(net256105), .ZN(n3756) );
  INV_X4 U4589 ( .A(n3756), .ZN(n3796) );
  NAND2_X2 U4590 ( .A1(n3640), .A2(n3637), .ZN(n3643) );
  AOI21_X4 U4591 ( .B1(n3641), .B2(n3640), .A(n3639), .ZN(n3642) );
  OAI21_X4 U4592 ( .B1(n3644), .B2(n3643), .A(n3642), .ZN(n3714) );
  NAND2_X2 U4593 ( .A1(n3714), .A2(n3645), .ZN(n3672) );
  NAND2_X2 U4594 ( .A1(a[23]), .A2(net256135), .ZN(n3668) );
  OAI211_X2 U4595 ( .C1(n3650), .C2(n3649), .A(n3648), .B(n3647), .ZN(n3652)
         );
  NAND2_X2 U4596 ( .A1(n3652), .A2(n3651), .ZN(n3653) );
  INV_X4 U4597 ( .A(n3653), .ZN(n3720) );
  NAND2_X2 U4598 ( .A1(a[24]), .A2(net256117), .ZN(n3663) );
  NAND2_X2 U4599 ( .A1(a[25]), .A2(net256143), .ZN(n3654) );
  NAND2_X2 U4600 ( .A1(a[26]), .A2(net256147), .ZN(n3655) );
  NAND2_X2 U4601 ( .A1(n3654), .A2(n3655), .ZN(n3657) );
  INV_X4 U4602 ( .A(n3655), .ZN(n3656) );
  NAND2_X2 U4603 ( .A1(n3657), .A2(n3723), .ZN(n3724) );
  NAND2_X2 U4604 ( .A1(n3659), .A2(n3658), .ZN(n3661) );
  XNOR2_X2 U4605 ( .A(n3724), .B(n3722), .ZN(n3664) );
  INV_X4 U4606 ( .A(n3664), .ZN(n3662) );
  NAND2_X2 U4607 ( .A1(n3663), .A2(n3662), .ZN(n3665) );
  NAND3_X2 U4608 ( .A1(a[24]), .A2(n3664), .A3(net256117), .ZN(n3718) );
  INV_X4 U4609 ( .A(n3719), .ZN(n3666) );
  XNOR2_X2 U4610 ( .A(n3720), .B(n3666), .ZN(n3669) );
  NAND2_X2 U4612 ( .A1(n3668), .A2(n3667), .ZN(n3715) );
  INV_X4 U4613 ( .A(n3668), .ZN(n3670) );
  NAND2_X2 U4615 ( .A1(n3715), .A2(n3836), .ZN(n3671) );
  XNOR2_X2 U4616 ( .A(n3672), .B(n3671), .ZN(n3675) );
  NAND2_X2 U4617 ( .A1(a[22]), .A2(net256125), .ZN(n3674) );
  NAND2_X2 U4618 ( .A1(n3673), .A2(n3674), .ZN(n3807) );
  INV_X4 U4619 ( .A(n3674), .ZN(n3676) );
  NAND2_X2 U4620 ( .A1(n3807), .A2(n3809), .ZN(n3684) );
  XNOR2_X2 U4621 ( .A(net253693), .B(net253694), .ZN(n3710) );
  XNOR2_X2 U4622 ( .A(n3687), .B(net253415), .ZN(n3697) );
  NAND2_X2 U4623 ( .A1(n1922), .A2(n1841), .ZN(n3694) );
  NAND2_X2 U4624 ( .A1(n3692), .A2(net253067), .ZN(n3693) );
  NAND2_X2 U4625 ( .A1(product_in[26]), .A2(net256095), .ZN(n3764) );
  XNOR2_X2 U4626 ( .A(n3765), .B(n3764), .ZN(n3696) );
  NOR2_X4 U4627 ( .A1(n3776), .A2(net253535), .ZN(n3699) );
  OAI21_X4 U4628 ( .B1(n3699), .B2(n3763), .A(n3790), .ZN(n3700) );
  NAND2_X2 U4630 ( .A1(a[22]), .A2(net256105), .ZN(n3801) );
  INV_X4 U4631 ( .A(n3801), .ZN(n3806) );
  INV_X4 U4632 ( .A(a[23]), .ZN(n3746) );
  OAI21_X4 U4633 ( .B1(n3717), .B2(n3716), .A(n3715), .ZN(n3835) );
  NAND2_X2 U4634 ( .A1(a[24]), .A2(net256135), .ZN(n3740) );
  OAI21_X4 U4635 ( .B1(n3720), .B2(n3719), .A(n3718), .ZN(n3721) );
  INV_X4 U4636 ( .A(n3721), .ZN(n3814) );
  NAND2_X2 U4637 ( .A1(a[25]), .A2(net256117), .ZN(n3734) );
  INV_X4 U4638 ( .A(n3722), .ZN(n3725) );
  OAI21_X4 U4639 ( .B1(n3725), .B2(n3724), .A(n3723), .ZN(n3730) );
  INV_X4 U4640 ( .A(n3730), .ZN(n3728) );
  INV_X4 U4641 ( .A(n3726), .ZN(n3817) );
  NAND2_X2 U4642 ( .A1(a[27]), .A2(net256151), .ZN(n3727) );
  INV_X4 U4643 ( .A(n3727), .ZN(n3816) );
  XNOR2_X2 U4644 ( .A(n3817), .B(n3816), .ZN(n3729) );
  NAND2_X2 U4645 ( .A1(n3728), .A2(n3729), .ZN(n3732) );
  INV_X4 U4646 ( .A(n3729), .ZN(n3731) );
  NAND2_X2 U4647 ( .A1(n3731), .A2(n3730), .ZN(n3818) );
  NAND2_X2 U4648 ( .A1(n3732), .A2(n3818), .ZN(n3733) );
  NAND2_X2 U4649 ( .A1(n3734), .A2(n3733), .ZN(n3737) );
  INV_X4 U4650 ( .A(n3733), .ZN(n3736) );
  INV_X4 U4651 ( .A(n3734), .ZN(n3735) );
  NAND2_X2 U4652 ( .A1(n3736), .A2(n3735), .ZN(n3812) );
  NAND2_X2 U4653 ( .A1(n3737), .A2(n3812), .ZN(n3813) );
  INV_X4 U4654 ( .A(n3813), .ZN(n3738) );
  XNOR2_X2 U4655 ( .A(n3814), .B(n3738), .ZN(n3741) );
  INV_X4 U4656 ( .A(n3741), .ZN(n3739) );
  NAND2_X2 U4657 ( .A1(n3740), .A2(n3739), .ZN(n3838) );
  INV_X4 U4658 ( .A(n3740), .ZN(n3742) );
  NAND2_X2 U4659 ( .A1(n3742), .A2(n3741), .ZN(n3839) );
  XNOR2_X2 U4660 ( .A(n3744), .B(n3743), .ZN(n3747) );
  OAI21_X4 U4661 ( .B1(n1648), .B2(n3746), .A(n3745), .ZN(n3899) );
  NAND2_X2 U4662 ( .A1(n3800), .A2(n3801), .ZN(n3748) );
  INV_X4 U4663 ( .A(n3748), .ZN(n3749) );
  XNOR2_X2 U4664 ( .A(n3750), .B(n3749), .ZN(n3754) );
  XNOR2_X2 U4665 ( .A(n3752), .B(n3751), .ZN(n3753) );
  NAND2_X2 U4666 ( .A1(a[21]), .A2(net256173), .ZN(net253450) );
  NAND2_X2 U4667 ( .A1(n1922), .A2(n3759), .ZN(n3760) );
  NAND2_X2 U4668 ( .A1(product_in[27]), .A2(net256095), .ZN(net253571) );
  INV_X4 U4669 ( .A(net253571), .ZN(net253569) );
  NAND2_X2 U4670 ( .A1(net253569), .A2(net253570), .ZN(net253177) );
  INV_X4 U4671 ( .A(n3763), .ZN(n3789) );
  INV_X4 U4672 ( .A(n3764), .ZN(n3766) );
  NAND2_X2 U4673 ( .A1(n3766), .A2(n3765), .ZN(net253533) );
  NAND2_X2 U4674 ( .A1(n3789), .A2(net253535), .ZN(n3770) );
  NOR2_X2 U4675 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  INV_X4 U4676 ( .A(n3780), .ZN(n3783) );
  NOR2_X4 U4677 ( .A1(n1828), .A2(n3781), .ZN(n3782) );
  NOR2_X4 U4678 ( .A1(n3783), .A2(n3782), .ZN(n3788) );
  OAI21_X4 U4679 ( .B1(n3786), .B2(n3785), .A(n3784), .ZN(net253188) );
  AOI21_X4 U4680 ( .B1(n3788), .B2(n3787), .A(net253188), .ZN(n3792) );
  NAND2_X2 U4681 ( .A1(net253533), .A2(n3790), .ZN(net253185) );
  OAI21_X4 U4682 ( .B1(n3792), .B2(n3791), .A(net257159), .ZN(n3926) );
  OAI21_X4 U4684 ( .B1(n3804), .B2(n3803), .A(n3862), .ZN(n3935) );
  NAND2_X2 U4685 ( .A1(n1870), .A2(n3939), .ZN(n3810) );
  OAI21_X4 U4686 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3815) );
  INV_X4 U4687 ( .A(n3815), .ZN(n3873) );
  NAND2_X2 U4688 ( .A1(n3817), .A2(n3816), .ZN(n3819) );
  NAND2_X2 U4689 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  INV_X4 U4690 ( .A(n3820), .ZN(n3876) );
  NAND2_X2 U4691 ( .A1(a[28]), .A2(net256147), .ZN(n3822) );
  NAND2_X2 U4692 ( .A1(n3821), .A2(n3822), .ZN(n3824) );
  INV_X4 U4693 ( .A(n3822), .ZN(n3823) );
  NAND2_X2 U4694 ( .A1(n3824), .A2(n3874), .ZN(n3875) );
  INV_X4 U4695 ( .A(n3875), .ZN(n3825) );
  XNOR2_X2 U4696 ( .A(n3876), .B(n3825), .ZN(n3827) );
  NAND2_X2 U4697 ( .A1(a[26]), .A2(net256117), .ZN(n3826) );
  NAND2_X2 U4698 ( .A1(n1826), .A2(n3826), .ZN(n3829) );
  INV_X4 U4699 ( .A(n3826), .ZN(n3828) );
  NAND2_X2 U4700 ( .A1(n3828), .A2(n3827), .ZN(n3871) );
  NAND2_X2 U4701 ( .A1(n3829), .A2(n3871), .ZN(n3872) );
  INV_X4 U4702 ( .A(n3872), .ZN(n3830) );
  XNOR2_X2 U4703 ( .A(n3873), .B(n3830), .ZN(n3833) );
  INV_X4 U4704 ( .A(n3833), .ZN(n3831) );
  NAND2_X2 U4705 ( .A1(a[25]), .A2(net256135), .ZN(n3832) );
  NAND2_X2 U4706 ( .A1(n3831), .A2(n3832), .ZN(n3867) );
  INV_X4 U4707 ( .A(n3832), .ZN(n3834) );
  NAND2_X2 U4708 ( .A1(n3834), .A2(n3833), .ZN(n3868) );
  INV_X4 U4709 ( .A(n3837), .ZN(n3841) );
  INV_X4 U4710 ( .A(n3838), .ZN(n3840) );
  OAI21_X4 U4711 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3866) );
  NAND2_X2 U4712 ( .A1(a[24]), .A2(net256125), .ZN(n3843) );
  INV_X4 U4713 ( .A(n3843), .ZN(n3845) );
  XNOR2_X2 U4714 ( .A(n3847), .B(n3846), .ZN(n3849) );
  NAND2_X2 U4715 ( .A1(a[23]), .A2(net256105), .ZN(n3848) );
  INV_X4 U4716 ( .A(n3848), .ZN(n3864) );
  XNOR2_X2 U4717 ( .A(net253462), .B(net253463), .ZN(n3850) );
  NAND2_X2 U4718 ( .A1(a[22]), .A2(net256173), .ZN(net253401) );
  INV_X4 U4719 ( .A(net253401), .ZN(net253460) );
  OAI21_X4 U4720 ( .B1(n1451), .B2(net253453), .A(net253323), .ZN(net253431)
         );
  XNOR2_X2 U4721 ( .A(net253451), .B(net253452), .ZN(net253442) );
  XNOR2_X2 U4722 ( .A(n1783), .B(n3853), .ZN(net253204) );
  NAND2_X2 U4723 ( .A1(net253421), .A2(net253205), .ZN(n3859) );
  OAI21_X4 U4724 ( .B1(net253393), .B2(net253392), .A(net257650), .ZN(n3912)
         );
  INV_X4 U4725 ( .A(n3867), .ZN(n3869) );
  OAI21_X4 U4726 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(n3948) );
  NAND2_X2 U4727 ( .A1(a[26]), .A2(net256135), .ZN(n3888) );
  OAI21_X4 U4728 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3889) );
  INV_X4 U4729 ( .A(n3889), .ZN(n3963) );
  OAI21_X4 U4730 ( .B1(n3876), .B2(n3875), .A(n3874), .ZN(n3880) );
  INV_X4 U4731 ( .A(n3880), .ZN(n3878) );
  NAND2_X2 U4732 ( .A1(a[29]), .A2(net256147), .ZN(n3877) );
  INV_X4 U4733 ( .A(n3877), .ZN(n3952) );
  XNOR2_X2 U4734 ( .A(n1429), .B(n3952), .ZN(n3879) );
  NAND2_X2 U4735 ( .A1(n3878), .A2(n3879), .ZN(n3882) );
  INV_X4 U4736 ( .A(n3879), .ZN(n3881) );
  NAND2_X2 U4737 ( .A1(n3881), .A2(n3880), .ZN(n3953) );
  NAND4_X2 U4738 ( .A1(a[27]), .A2(n3882), .A3(n3953), .A4(net256117), .ZN(
        n3961) );
  INV_X4 U4739 ( .A(n3882), .ZN(n3885) );
  INV_X4 U4740 ( .A(n3953), .ZN(n3884) );
  NAND2_X2 U4741 ( .A1(a[27]), .A2(net256117), .ZN(n3883) );
  OAI21_X4 U4742 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(n3886) );
  NAND2_X2 U4743 ( .A1(n3961), .A2(n3886), .ZN(n3962) );
  XNOR2_X2 U4744 ( .A(n3963), .B(n3962), .ZN(n3887) );
  NAND2_X2 U4745 ( .A1(n3888), .A2(n3887), .ZN(n3947) );
  XNOR2_X2 U4746 ( .A(n3889), .B(n3962), .ZN(n3890) );
  NAND3_X2 U4747 ( .A1(n3890), .A2(net256135), .A3(a[26]), .ZN(n3949) );
  NAND2_X2 U4748 ( .A1(n3947), .A2(n3949), .ZN(n3891) );
  XNOR2_X2 U4749 ( .A(n3948), .B(n3891), .ZN(n3894) );
  NAND2_X2 U4750 ( .A1(a[25]), .A2(net256125), .ZN(n3893) );
  NAND2_X2 U4751 ( .A1(n3892), .A2(n3893), .ZN(n3896) );
  INV_X4 U4752 ( .A(n3893), .ZN(n3895) );
  NAND2_X2 U4753 ( .A1(n3895), .A2(n3894), .ZN(n3944) );
  INV_X4 U4754 ( .A(n3945), .ZN(n3904) );
  INV_X4 U4755 ( .A(n3942), .ZN(n3901) );
  NAND2_X2 U4756 ( .A1(a[24]), .A2(net256105), .ZN(n3905) );
  NAND2_X2 U4757 ( .A1(n3905), .A2(n1871), .ZN(n3937) );
  INV_X4 U4758 ( .A(n3905), .ZN(n3906) );
  XNOR2_X2 U4759 ( .A(n3908), .B(n3907), .ZN(n3914) );
  INV_X4 U4760 ( .A(n1938), .ZN(n3909) );
  NAND2_X2 U4761 ( .A1(a[23]), .A2(net256173), .ZN(n3913) );
  INV_X4 U4762 ( .A(n3913), .ZN(n3910) );
  XNOR2_X2 U4763 ( .A(n3912), .B(n3911), .ZN(net253279) );
  NAND2_X2 U4764 ( .A1(product_in[29]), .A2(net253304), .ZN(net253194) );
  INV_X4 U4765 ( .A(net253173), .ZN(net253301) );
  NAND2_X2 U4766 ( .A1(n1958), .A2(net253287), .ZN(n3920) );
  OAI21_X4 U4767 ( .B1(n3922), .B2(n3921), .A(n3920), .ZN(n3923) );
  INV_X4 U4768 ( .A(net253177), .ZN(net253294) );
  INV_X4 U4769 ( .A(net253287), .ZN(net253295) );
  NOR2_X4 U4770 ( .A1(net253294), .A2(net253295), .ZN(n3924) );
  NAND2_X2 U4771 ( .A1(n3924), .A2(net253194), .ZN(n3925) );
  NOR2_X4 U4772 ( .A1(n3927), .A2(net253289), .ZN(n3930) );
  NAND2_X2 U4773 ( .A1(net253287), .A2(net253194), .ZN(n3929) );
  OAI21_X4 U4774 ( .B1(n3930), .B2(n3929), .A(n3928), .ZN(n3931) );
  NOR2_X4 U4775 ( .A1(n3931), .A2(n3932), .ZN(n3991) );
  NAND2_X2 U4776 ( .A1(a[24]), .A2(net256175), .ZN(n4003) );
  NAND2_X2 U4777 ( .A1(a[23]), .A2(net256165), .ZN(n4073) );
  INV_X4 U4778 ( .A(n3975), .ZN(n3972) );
  NAND3_X2 U4779 ( .A1(n3936), .A2(n3937), .A3(n1115), .ZN(n3976) );
  INV_X4 U4780 ( .A(n3976), .ZN(n3971) );
  INV_X4 U4781 ( .A(n3947), .ZN(n3951) );
  INV_X4 U4782 ( .A(n3948), .ZN(n3950) );
  OAI21_X4 U4783 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3967) );
  INV_X4 U4784 ( .A(n3967), .ZN(n3965) );
  NAND2_X2 U4785 ( .A1(n1429), .A2(n3952), .ZN(n3954) );
  NAND2_X2 U4786 ( .A1(n3954), .A2(n3953), .ZN(n4025) );
  NAND2_X2 U4787 ( .A1(a[30]), .A2(net256151), .ZN(n3958) );
  INV_X4 U4788 ( .A(n3958), .ZN(n3957) );
  NAND2_X2 U4789 ( .A1(a[29]), .A2(net256143), .ZN(n3959) );
  INV_X4 U4790 ( .A(n3959), .ZN(n3956) );
  NAND2_X2 U4791 ( .A1(n3957), .A2(n3956), .ZN(n4033) );
  NAND2_X2 U4792 ( .A1(n3959), .A2(n3958), .ZN(n3960) );
  NAND2_X2 U4793 ( .A1(n4033), .A2(n3960), .ZN(n4024) );
  XNOR2_X2 U4794 ( .A(n4025), .B(n4024), .ZN(n4022) );
  NAND2_X2 U4795 ( .A1(a[28]), .A2(net256117), .ZN(n4021) );
  XNOR2_X2 U4796 ( .A(n4022), .B(n4021), .ZN(n4020) );
  OAI21_X4 U4797 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(n4019) );
  NAND2_X2 U4798 ( .A1(a[27]), .A2(net256135), .ZN(n4015) );
  XNOR2_X2 U4799 ( .A(n4019), .B(n4015), .ZN(n3964) );
  XNOR2_X2 U4800 ( .A(n4020), .B(n3964), .ZN(n3966) );
  NAND2_X2 U4801 ( .A1(n3965), .A2(n3966), .ZN(n4012) );
  NAND2_X2 U4802 ( .A1(n3968), .A2(n3967), .ZN(n4011) );
  NAND2_X2 U4803 ( .A1(a[26]), .A2(net256125), .ZN(n4014) );
  XNOR2_X2 U4804 ( .A(n3969), .B(n4014), .ZN(n4004) );
  NAND2_X2 U4805 ( .A1(a[25]), .A2(net253103), .ZN(n4005) );
  XNOR2_X2 U4806 ( .A(n4004), .B(n4005), .ZN(n3970) );
  XNOR2_X2 U4807 ( .A(n3970), .B(n4010), .ZN(n3973) );
  OAI21_X4 U4808 ( .B1(n3972), .B2(n3971), .A(n1116), .ZN(n4001) );
  INV_X4 U4809 ( .A(n3992), .ZN(n3977) );
  NOR2_X4 U4810 ( .A1(n3977), .A2(net253220), .ZN(n3979) );
  NAND2_X2 U4811 ( .A1(n3983), .A2(net253067), .ZN(n3984) );
  NAND2_X2 U4812 ( .A1(n3987), .A2(net256095), .ZN(net253192) );
  NAND2_X2 U4813 ( .A1(product_in[30]), .A2(net256095), .ZN(net253193) );
  INV_X4 U4814 ( .A(net253193), .ZN(net253191) );
  NAND2_X2 U4815 ( .A1(net253191), .A2(net253192), .ZN(net253163) );
  INV_X4 U4816 ( .A(n3999), .ZN(n4072) );
  NAND2_X2 U4817 ( .A1(n4071), .A2(n4072), .ZN(n4066) );
  INV_X4 U4818 ( .A(n1112), .ZN(n4009) );
  XNOR2_X2 U4819 ( .A(n4009), .B(n4010), .ZN(n4006) );
  NOR2_X4 U4820 ( .A1(n4008), .A2(n4007), .ZN(n4062) );
  NAND2_X2 U4821 ( .A1(n4010), .A2(n4009), .ZN(n4060) );
  XNOR2_X2 U4822 ( .A(n4020), .B(n4019), .ZN(n4016) );
  NOR2_X2 U4823 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  NOR2_X4 U4824 ( .A1(n4018), .A2(n4017), .ZN(n4056) );
  NAND2_X2 U4825 ( .A1(n4020), .A2(n4019), .ZN(n4054) );
  INV_X4 U4826 ( .A(n4021), .ZN(n4023) );
  NAND2_X2 U4827 ( .A1(n4023), .A2(n4022), .ZN(n4052) );
  INV_X4 U4828 ( .A(n4024), .ZN(n4026) );
  NAND2_X2 U4829 ( .A1(n4026), .A2(n4025), .ZN(n4050) );
  INV_X4 U4830 ( .A(a[31]), .ZN(n4027) );
  INV_X4 U4831 ( .A(a[30]), .ZN(n4028) );
  INV_X4 U4832 ( .A(a[24]), .ZN(n4029) );
  NOR2_X4 U4833 ( .A1(net256167), .A2(n4029), .ZN(n4030) );
  FA_X1 U4834 ( .A(n4032), .B(n4031), .CI(n4030), .S(n4036) );
  INV_X4 U4835 ( .A(n4033), .ZN(n4034) );
  INV_X4 U4836 ( .A(a[29]), .ZN(net253111) );
  XNOR2_X2 U4837 ( .A(n4034), .B(net253109), .ZN(n4035) );
  XNOR2_X2 U4838 ( .A(n4036), .B(n4035), .ZN(n4048) );
  INV_X4 U4839 ( .A(a[25]), .ZN(n4037) );
  INV_X4 U4840 ( .A(a[26]), .ZN(n4038) );
  XOR2_X2 U4841 ( .A(n4040), .B(n4039), .Z(n4046) );
  INV_X4 U4842 ( .A(a[27]), .ZN(n4041) );
  NOR2_X4 U4843 ( .A1(n1648), .A2(n4041), .ZN(n4044) );
  INV_X4 U4844 ( .A(a[28]), .ZN(n4042) );
  NOR2_X4 U4845 ( .A1(net256139), .A2(n4042), .ZN(n4043) );
  XNOR2_X2 U4846 ( .A(n4044), .B(n4043), .ZN(n4045) );
  XNOR2_X2 U4847 ( .A(n4046), .B(n4045), .ZN(n4047) );
  XNOR2_X2 U4848 ( .A(n4048), .B(n4047), .ZN(n4049) );
  XNOR2_X2 U4849 ( .A(n4050), .B(n4049), .ZN(n4051) );
  XNOR2_X2 U4850 ( .A(n4052), .B(n4051), .ZN(n4053) );
  XNOR2_X2 U4851 ( .A(n4054), .B(n4053), .ZN(n4055) );
  XNOR2_X2 U4852 ( .A(n4056), .B(n4055), .ZN(n4057) );
  XNOR2_X2 U4853 ( .A(n4058), .B(n4057), .ZN(n4059) );
  XNOR2_X2 U4854 ( .A(n4060), .B(n4059), .ZN(n4061) );
  XNOR2_X2 U4855 ( .A(n4062), .B(n4061), .ZN(n4063) );
  XNOR2_X2 U4856 ( .A(n4064), .B(n4063), .ZN(n4065) );
  XNOR2_X2 U4857 ( .A(n4066), .B(n4065), .ZN(net253044) );
  NAND2_X2 U4858 ( .A1(net253067), .A2(n4068), .ZN(n4069) );
  NAND2_X2 U4859 ( .A1(product_in[31]), .A2(net256095), .ZN(net253050) );
  XNOR2_X2 U4860 ( .A(n4072), .B(n4071), .ZN(n4074) );
  INV_X1 U1145 ( .A(net254364), .ZN(n1106) );
  INV_X2 U1161 ( .A(net255581), .ZN(net255454) );
  XNOR2_X2 U1165 ( .A(n3241), .B(n3240), .ZN(n4086) );
  OAI21_X2 U1172 ( .B1(n3608), .B2(n3609), .A(net253823), .ZN(net253586) );
  INV_X2 U1180 ( .A(net254682), .ZN(net254952) );
  INV_X2 U1189 ( .A(n3669), .ZN(n3667) );
  NAND2_X4 U1201 ( .A1(n3670), .A2(n3669), .ZN(n3836) );
  OAI21_X2 U1206 ( .B1(n3578), .B2(n3577), .A(n3660), .ZN(n3579) );
  INV_X2 U1214 ( .A(n3363), .ZN(n3365) );
  INV_X4 U1225 ( .A(n2619), .ZN(n2750) );
  INV_X4 U1227 ( .A(n2680), .ZN(n1918) );
  NAND2_X4 U1241 ( .A1(n3166), .A2(n3167), .ZN(n4087) );
  NAND2_X2 U1244 ( .A1(n3166), .A2(n3167), .ZN(n3273) );
  XNOR2_X2 U1251 ( .A(n3104), .B(n1845), .ZN(product_out[20]) );
  INV_X4 U1257 ( .A(n3104), .ZN(n3268) );
  INV_X1 U1359 ( .A(n1933), .ZN(n3264) );
  INV_X2 U1361 ( .A(n3264), .ZN(n1845) );
  NAND2_X2 U1386 ( .A1(n1365), .A2(n1366), .ZN(n1368) );
  NAND2_X2 U1395 ( .A1(n2166), .A2(n2165), .ZN(n1367) );
  AND2_X2 U1405 ( .A1(n1821), .A2(n1583), .ZN(n4088) );
  NAND2_X4 U1422 ( .A1(n1272), .A2(n1300), .ZN(n1821) );
  AND2_X2 U1490 ( .A1(n1821), .A2(n1583), .ZN(n1847) );
  OAI21_X4 U1514 ( .B1(net254575), .B2(net254576), .A(net257864), .ZN(n3073)
         );
  INV_X8 U1515 ( .A(n1919), .ZN(n3076) );
  NAND2_X4 U1620 ( .A1(n1353), .A2(n1354), .ZN(n1919) );
  CLKBUF_X2 U1668 ( .A(n3474), .Z(n1850) );
  INV_X4 U1682 ( .A(n3701), .ZN(n4089) );
  INV_X2 U1704 ( .A(n3701), .ZN(n3705) );
  INV_X1 U1786 ( .A(n3768), .ZN(n4090) );
  INV_X8 U1787 ( .A(net253433), .ZN(net253415) );
  NAND2_X2 U1788 ( .A1(n3855), .A2(n3856), .ZN(n3625) );
  CLKBUF_X3 U1796 ( .A(n3281), .Z(n1340) );
  INV_X1 U1826 ( .A(n1943), .ZN(n4091) );
  INV_X2 U1865 ( .A(n4091), .ZN(n4092) );
  AND3_X2 U1867 ( .A1(net253776), .A2(n3472), .A3(net257109), .ZN(n1880) );
  OR2_X2 U1889 ( .A1(n3539), .A2(n1879), .ZN(n3475) );
  INV_X2 U1890 ( .A(n3523), .ZN(n3524) );
  INV_X1 U1905 ( .A(n3274), .ZN(n1164) );
  INV_X4 U1929 ( .A(n2641), .ZN(n1576) );
  OAI21_X2 U1934 ( .B1(n2569), .B2(n2568), .A(n1435), .ZN(n2641) );
  NAND2_X4 U1952 ( .A1(n3180), .A2(n1995), .ZN(n2921) );
  NAND2_X4 U1968 ( .A1(n3504), .A2(n4094), .ZN(n1803) );
  NAND2_X2 U1979 ( .A1(n2920), .A2(n1416), .ZN(n4093) );
  INV_X8 U1980 ( .A(n3633), .ZN(n3624) );
  NAND2_X4 U1996 ( .A1(n1395), .A2(n1396), .ZN(n3633) );
  NAND2_X2 U2091 ( .A1(n3624), .A2(n3623), .ZN(n3854) );
  NOR2_X2 U2099 ( .A1(n3494), .A2(n3781), .ZN(n4094) );
  INV_X8 U2103 ( .A(n3492), .ZN(n3494) );
  INV_X2 U2105 ( .A(net255040), .ZN(n1217) );
  AOI21_X2 U2136 ( .B1(n3926), .B2(net257211), .A(n3925), .ZN(n3932) );
  NOR2_X2 U2137 ( .A1(net256159), .A2(n2071), .ZN(n4097) );
  INV_X2 U2144 ( .A(n3533), .ZN(n4095) );
  XNOR2_X2 U2152 ( .A(n1967), .B(n4097), .ZN(n4096) );
  CLKBUF_X2 U2161 ( .A(n2020), .Z(n4098) );
  NAND2_X1 U2220 ( .A1(n1922), .A2(n3794), .ZN(net253525) );
  INV_X2 U2242 ( .A(n2119), .ZN(n4099) );
  INV_X4 U2243 ( .A(n4099), .ZN(n4100) );
  INV_X4 U2248 ( .A(n1128), .ZN(n4101) );
  NAND2_X4 U2254 ( .A1(n3339), .A2(n1183), .ZN(n1128) );
  NAND2_X4 U2289 ( .A1(n3534), .A2(n3535), .ZN(n3474) );
  NOR2_X2 U2447 ( .A1(n3285), .A2(n3284), .ZN(n3286) );
  INV_X4 U2451 ( .A(net254366), .ZN(net254575) );
  INV_X4 U2458 ( .A(net253776), .ZN(net254059) );
  XNOR2_X2 U2503 ( .A(n1394), .B(n3615), .ZN(n4102) );
  INV_X2 U2593 ( .A(n1545), .ZN(n1546) );
  XNOR2_X2 U2603 ( .A(n1912), .B(n1824), .ZN(n1827) );
  NAND2_X2 U2641 ( .A1(n2237), .A2(n2236), .ZN(n2290) );
  AND2_X2 U2645 ( .A1(n2211), .A2(n2212), .ZN(n4103) );
  NAND2_X4 U2650 ( .A1(a[3]), .A2(net256127), .ZN(n2212) );
  INV_X8 U2879 ( .A(n1925), .ZN(n1926) );
  INV_X4 U2908 ( .A(n3027), .ZN(n4104) );
  INV_X1 U2914 ( .A(n3027), .ZN(n1438) );
  INV_X1 U2916 ( .A(n3166), .ZN(n4105) );
  INV_X2 U2925 ( .A(n4105), .ZN(n4106) );
  NAND2_X1 U2942 ( .A1(n4106), .A2(n3167), .ZN(n4107) );
  CLKBUF_X2 U2973 ( .A(n3513), .Z(n4108) );
  OAI21_X1 U3029 ( .B1(n2417), .B2(n2416), .A(n2415), .ZN(n4109) );
  INV_X8 U3127 ( .A(n2414), .ZN(n2417) );
  INV_X4 U3131 ( .A(n2947), .ZN(n4110) );
  NAND2_X1 U3141 ( .A1(n2175), .A2(n2174), .ZN(n2178) );
  NAND2_X4 U3206 ( .A1(net255327), .A2(net255329), .ZN(net255498) );
  INV_X4 U3329 ( .A(n3919), .ZN(n3922) );
  NAND2_X2 U3365 ( .A1(n3080), .A2(n3081), .ZN(n1842) );
  NAND2_X4 U3527 ( .A1(n3082), .A2(n3083), .ZN(n3523) );
  AOI21_X2 U3599 ( .B1(n3526), .B2(n1300), .A(n3524), .ZN(n3531) );
  NAND2_X2 U3625 ( .A1(n1123), .A2(n3072), .ZN(n1353) );
  NAND2_X4 U3628 ( .A1(n3190), .A2(n1107), .ZN(n3072) );
  NOR2_X4 U3641 ( .A1(n1568), .A2(net257672), .ZN(n3793) );
  INV_X1 U3659 ( .A(n2662), .ZN(n1431) );
  INV_X8 U3685 ( .A(n1950), .ZN(n2923) );
  XNOR2_X2 U3708 ( .A(n3171), .B(n3267), .ZN(n1933) );
  INV_X2 U3710 ( .A(n3004), .ZN(n1174) );
  XNOR2_X2 U3725 ( .A(n2724), .B(n4112), .ZN(n4111) );
  INV_X4 U3738 ( .A(n4111), .ZN(n3982) );
  AND2_X2 U3858 ( .A1(n3013), .A2(n2735), .ZN(n4112) );
  NAND2_X2 U3874 ( .A1(n3622), .A2(n3621), .ZN(n1395) );
  XNOR2_X1 U3876 ( .A(n2396), .B(n2395), .ZN(n4113) );
  BUF_X4 U3995 ( .A(n2652), .Z(n1435) );
  NAND2_X2 U4018 ( .A1(n2657), .A2(n2652), .ZN(n2561) );
  INV_X2 U4079 ( .A(n1248), .ZN(n1218) );
  OAI21_X4 U4139 ( .B1(net253393), .B2(net253392), .A(net257650), .ZN(n1124)
         );
  OAI211_X4 U4142 ( .C1(n1185), .C2(n1184), .A(n2844), .B(n1187), .ZN(n3176)
         );
  INV_X2 U4143 ( .A(net254856), .ZN(n1185) );
  NAND2_X4 U4299 ( .A1(n3151), .A2(n3152), .ZN(net254291) );
  NOR2_X4 U4304 ( .A1(n1585), .A2(n2881), .ZN(n1586) );
  NAND2_X4 U4407 ( .A1(net255770), .A2(n2208), .ZN(n2320) );
  INV_X1 U4459 ( .A(n2207), .ZN(n2208) );
  NAND3_X2 U4562 ( .A1(n2715), .A2(n1219), .A3(n1220), .ZN(n2742) );
  INV_X2 U4581 ( .A(n2712), .ZN(n2715) );
  OAI211_X2 U4611 ( .C1(n1905), .C2(net253064), .A(n3985), .B(n3984), .ZN(
        n3988) );
  NAND2_X2 U4614 ( .A1(net253301), .A2(net253302), .ZN(net253287) );
  NAND2_X4 U4629 ( .A1(n3993), .A2(n3996), .ZN(n3978) );
  NAND2_X2 U4683 ( .A1(n1747), .A2(net253398), .ZN(n1746) );
  NAND2_X2 U4861 ( .A1(net253169), .A2(n4114), .ZN(n4115) );
  INV_X4 U4862 ( .A(n1636), .ZN(n4114) );
  INV_X4 U4863 ( .A(n4115), .ZN(net253166) );
  NAND2_X2 U4864 ( .A1(net255225), .A2(n2578), .ZN(net255091) );
  NAND2_X4 U4865 ( .A1(n1741), .A2(n1740), .ZN(n1434) );
  INV_X4 U4866 ( .A(net254857), .ZN(n1741) );
  AOI21_X4 U4867 ( .B1(n1658), .B2(n1657), .A(n1659), .ZN(n1653) );
  INV_X8 U4868 ( .A(net253043), .ZN(n1658) );
  OAI211_X4 U4869 ( .C1(n3681), .C2(n3682), .A(n3679), .B(n3680), .ZN(n3711)
         );
  INV_X4 U4870 ( .A(n3550), .ZN(n3682) );
  INV_X2 U4871 ( .A(n3678), .ZN(n3679) );
  AOI21_X4 U4872 ( .B1(n3856), .B2(n3855), .A(n3854), .ZN(n3708) );
  OAI21_X4 U4873 ( .B1(n2611), .B2(net255179), .A(n2610), .ZN(n2679) );
  INV_X4 U4874 ( .A(n2432), .ZN(n2610) );
endmodule

