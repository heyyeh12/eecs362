module wb(memRd, regWr, target, memWrData);
    
    input memRd;

endmodule // wb