
module dffa_N_BITS32 ( d, clk, rst, enable, q, aload, arst );
  input [31:0] d;
  output [31:0] q;
  input [31:0] aload;
  input clk, rst, enable, arst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262;

  DFFRS_X1 q_reg_31_ ( .D(n128), .CK(clk), .RN(n163), .SN(n126), .Q(q[31]), 
        .QN(n127) );
  DFFRS_X1 q_reg_30_ ( .D(n125), .CK(clk), .RN(n164), .SN(n123), .Q(q[30]), 
        .QN(n124) );
  DFFRS_X1 q_reg_29_ ( .D(n122), .CK(clk), .RN(n165), .SN(n120), .Q(q[29]), 
        .QN(n121) );
  DFFRS_X1 q_reg_28_ ( .D(n119), .CK(clk), .RN(n166), .SN(n117), .Q(q[28]), 
        .QN(n118) );
  DFFRS_X1 q_reg_27_ ( .D(n116), .CK(clk), .RN(n167), .SN(n114), .Q(q[27]), 
        .QN(n115) );
  DFFRS_X1 q_reg_26_ ( .D(n113), .CK(clk), .RN(n168), .SN(n111), .Q(q[26]), 
        .QN(n112) );
  DFFRS_X1 q_reg_25_ ( .D(n110), .CK(clk), .RN(n169), .SN(n108), .Q(q[25]), 
        .QN(n109) );
  DFFRS_X1 q_reg_24_ ( .D(n107), .CK(clk), .RN(n170), .SN(n105), .Q(q[24]), 
        .QN(n106) );
  DFFRS_X1 q_reg_23_ ( .D(n104), .CK(clk), .RN(n171), .SN(n102), .Q(q[23]), 
        .QN(n103) );
  DFFRS_X1 q_reg_22_ ( .D(n101), .CK(clk), .RN(n172), .SN(n99), .Q(q[22]), 
        .QN(n100) );
  DFFRS_X1 q_reg_21_ ( .D(n98), .CK(clk), .RN(n173), .SN(n96), .Q(q[21]), .QN(
        n97) );
  DFFRS_X1 q_reg_20_ ( .D(n95), .CK(clk), .RN(n174), .SN(n93), .Q(q[20]), .QN(
        n94) );
  DFFRS_X1 q_reg_19_ ( .D(n92), .CK(clk), .RN(n175), .SN(n90), .Q(q[19]), .QN(
        n91) );
  DFFRS_X1 q_reg_18_ ( .D(n89), .CK(clk), .RN(n176), .SN(n87), .Q(q[18]), .QN(
        n88) );
  DFFRS_X1 q_reg_17_ ( .D(n86), .CK(clk), .RN(n177), .SN(n84), .Q(q[17]), .QN(
        n85) );
  DFFRS_X1 q_reg_16_ ( .D(n83), .CK(clk), .RN(n178), .SN(n81), .Q(q[16]), .QN(
        n82) );
  DFFRS_X1 q_reg_15_ ( .D(n80), .CK(clk), .RN(n179), .SN(n78), .Q(q[15]), .QN(
        n79) );
  DFFRS_X1 q_reg_14_ ( .D(n77), .CK(clk), .RN(n180), .SN(n75), .Q(q[14]), .QN(
        n76) );
  DFFRS_X1 q_reg_13_ ( .D(n74), .CK(clk), .RN(n181), .SN(n72), .Q(q[13]), .QN(
        n73) );
  DFFRS_X1 q_reg_12_ ( .D(n71), .CK(clk), .RN(n182), .SN(n69), .Q(q[12]), .QN(
        n70) );
  DFFRS_X1 q_reg_11_ ( .D(n68), .CK(clk), .RN(n183), .SN(n66), .Q(q[11]), .QN(
        n67) );
  DFFRS_X1 q_reg_10_ ( .D(n65), .CK(clk), .RN(n184), .SN(n63), .Q(q[10]), .QN(
        n64) );
  DFFRS_X1 q_reg_9_ ( .D(n62), .CK(clk), .RN(n185), .SN(n60), .Q(q[9]), .QN(
        n61) );
  DFFRS_X1 q_reg_8_ ( .D(n59), .CK(clk), .RN(n186), .SN(n57), .Q(q[8]), .QN(
        n58) );
  DFFRS_X1 q_reg_7_ ( .D(n56), .CK(clk), .RN(n187), .SN(n54), .Q(q[7]), .QN(
        n55) );
  DFFRS_X1 q_reg_6_ ( .D(n53), .CK(clk), .RN(n188), .SN(n51), .Q(q[6]), .QN(
        n52) );
  DFFRS_X1 q_reg_5_ ( .D(n50), .CK(clk), .RN(n189), .SN(n48), .Q(q[5]), .QN(
        n49) );
  DFFRS_X1 q_reg_4_ ( .D(n47), .CK(clk), .RN(n190), .SN(n45), .Q(q[4]), .QN(
        n46) );
  DFFRS_X1 q_reg_3_ ( .D(n44), .CK(clk), .RN(n191), .SN(n42), .Q(q[3]), .QN(
        n43) );
  DFFRS_X1 q_reg_2_ ( .D(n41), .CK(clk), .RN(n192), .SN(n39), .Q(q[2]), .QN(
        n40) );
  DFFRS_X1 q_reg_1_ ( .D(n38), .CK(clk), .RN(n193), .SN(n36), .Q(q[1]), .QN(
        n37) );
  DFFRS_X1 q_reg_0_ ( .D(n35), .CK(clk), .RN(n194), .SN(n33), .Q(q[0]), .QN(
        n34) );
  OAI21_X1 U3 ( .B1(enable), .B2(n34), .A(n1), .ZN(n35) );
  NAND2_X1 U4 ( .A1(enable), .A2(d[0]), .ZN(n1) );
  OAI21_X1 U5 ( .B1(enable), .B2(n37), .A(n2), .ZN(n38) );
  NAND2_X1 U6 ( .A1(d[1]), .A2(enable), .ZN(n2) );
  OAI21_X1 U7 ( .B1(enable), .B2(n40), .A(n3), .ZN(n41) );
  NAND2_X1 U8 ( .A1(d[2]), .A2(enable), .ZN(n3) );
  OAI21_X1 U9 ( .B1(enable), .B2(n43), .A(n4), .ZN(n44) );
  NAND2_X1 U10 ( .A1(d[3]), .A2(enable), .ZN(n4) );
  OAI21_X1 U11 ( .B1(enable), .B2(n46), .A(n5), .ZN(n47) );
  NAND2_X1 U12 ( .A1(d[4]), .A2(enable), .ZN(n5) );
  OAI21_X1 U13 ( .B1(enable), .B2(n49), .A(n6), .ZN(n50) );
  NAND2_X1 U14 ( .A1(d[5]), .A2(enable), .ZN(n6) );
  OAI21_X1 U15 ( .B1(enable), .B2(n52), .A(n7), .ZN(n53) );
  NAND2_X1 U16 ( .A1(d[6]), .A2(enable), .ZN(n7) );
  OAI21_X1 U17 ( .B1(enable), .B2(n55), .A(n8), .ZN(n56) );
  NAND2_X1 U18 ( .A1(d[7]), .A2(enable), .ZN(n8) );
  OAI21_X1 U19 ( .B1(enable), .B2(n58), .A(n9), .ZN(n59) );
  NAND2_X1 U20 ( .A1(d[8]), .A2(enable), .ZN(n9) );
  OAI21_X1 U21 ( .B1(enable), .B2(n61), .A(n10), .ZN(n62) );
  NAND2_X1 U22 ( .A1(d[9]), .A2(enable), .ZN(n10) );
  OAI21_X1 U23 ( .B1(enable), .B2(n64), .A(n11), .ZN(n65) );
  NAND2_X1 U24 ( .A1(d[10]), .A2(enable), .ZN(n11) );
  OAI21_X1 U25 ( .B1(enable), .B2(n67), .A(n12), .ZN(n68) );
  NAND2_X1 U26 ( .A1(d[11]), .A2(enable), .ZN(n12) );
  OAI21_X1 U27 ( .B1(enable), .B2(n70), .A(n13), .ZN(n71) );
  NAND2_X1 U28 ( .A1(d[12]), .A2(enable), .ZN(n13) );
  OAI21_X1 U29 ( .B1(enable), .B2(n73), .A(n14), .ZN(n74) );
  NAND2_X1 U30 ( .A1(d[13]), .A2(enable), .ZN(n14) );
  OAI21_X1 U31 ( .B1(enable), .B2(n76), .A(n15), .ZN(n77) );
  NAND2_X1 U32 ( .A1(d[14]), .A2(enable), .ZN(n15) );
  OAI21_X1 U33 ( .B1(enable), .B2(n79), .A(n16), .ZN(n80) );
  NAND2_X1 U34 ( .A1(d[15]), .A2(enable), .ZN(n16) );
  OAI21_X1 U35 ( .B1(enable), .B2(n82), .A(n17), .ZN(n83) );
  NAND2_X1 U36 ( .A1(d[16]), .A2(enable), .ZN(n17) );
  OAI21_X1 U37 ( .B1(enable), .B2(n85), .A(n18), .ZN(n86) );
  NAND2_X1 U38 ( .A1(d[17]), .A2(enable), .ZN(n18) );
  OAI21_X1 U39 ( .B1(enable), .B2(n88), .A(n19), .ZN(n89) );
  NAND2_X1 U40 ( .A1(d[18]), .A2(enable), .ZN(n19) );
  OAI21_X1 U41 ( .B1(enable), .B2(n91), .A(n20), .ZN(n92) );
  NAND2_X1 U42 ( .A1(d[19]), .A2(enable), .ZN(n20) );
  OAI21_X1 U43 ( .B1(enable), .B2(n94), .A(n21), .ZN(n95) );
  NAND2_X1 U44 ( .A1(d[20]), .A2(enable), .ZN(n21) );
  OAI21_X1 U45 ( .B1(enable), .B2(n97), .A(n22), .ZN(n98) );
  NAND2_X1 U46 ( .A1(d[21]), .A2(enable), .ZN(n22) );
  OAI21_X1 U47 ( .B1(enable), .B2(n100), .A(n23), .ZN(n101) );
  NAND2_X1 U48 ( .A1(d[22]), .A2(enable), .ZN(n23) );
  OAI21_X1 U49 ( .B1(enable), .B2(n103), .A(n24), .ZN(n104) );
  NAND2_X1 U50 ( .A1(d[23]), .A2(enable), .ZN(n24) );
  OAI21_X1 U51 ( .B1(enable), .B2(n106), .A(n25), .ZN(n107) );
  NAND2_X1 U52 ( .A1(d[24]), .A2(enable), .ZN(n25) );
  OAI21_X1 U53 ( .B1(enable), .B2(n109), .A(n26), .ZN(n110) );
  NAND2_X1 U54 ( .A1(d[25]), .A2(enable), .ZN(n26) );
  OAI21_X1 U55 ( .B1(enable), .B2(n112), .A(n27), .ZN(n113) );
  NAND2_X1 U56 ( .A1(d[26]), .A2(enable), .ZN(n27) );
  OAI21_X1 U57 ( .B1(enable), .B2(n115), .A(n28), .ZN(n116) );
  NAND2_X1 U58 ( .A1(d[27]), .A2(enable), .ZN(n28) );
  OAI21_X1 U59 ( .B1(enable), .B2(n118), .A(n29), .ZN(n119) );
  NAND2_X1 U60 ( .A1(d[28]), .A2(enable), .ZN(n29) );
  OAI21_X1 U61 ( .B1(enable), .B2(n121), .A(n30), .ZN(n122) );
  NAND2_X1 U62 ( .A1(d[29]), .A2(enable), .ZN(n30) );
  OAI21_X1 U63 ( .B1(enable), .B2(n124), .A(n31), .ZN(n125) );
  NAND2_X1 U64 ( .A1(d[30]), .A2(enable), .ZN(n31) );
  OAI21_X1 U65 ( .B1(enable), .B2(n127), .A(n32), .ZN(n128) );
  NAND2_X1 U66 ( .A1(d[31]), .A2(enable), .ZN(n32) );
  INV_X4 U67 ( .A(n196), .ZN(n33) );
  INV_X4 U68 ( .A(n198), .ZN(n36) );
  INV_X4 U69 ( .A(n200), .ZN(n39) );
  INV_X4 U70 ( .A(n202), .ZN(n42) );
  INV_X4 U71 ( .A(n204), .ZN(n45) );
  INV_X4 U72 ( .A(n206), .ZN(n48) );
  INV_X4 U73 ( .A(n208), .ZN(n51) );
  INV_X4 U74 ( .A(n210), .ZN(n54) );
  INV_X4 U75 ( .A(n212), .ZN(n57) );
  INV_X4 U76 ( .A(n214), .ZN(n60) );
  INV_X4 U77 ( .A(n216), .ZN(n63) );
  INV_X4 U78 ( .A(n218), .ZN(n66) );
  INV_X4 U79 ( .A(n220), .ZN(n69) );
  INV_X4 U80 ( .A(n222), .ZN(n72) );
  INV_X4 U81 ( .A(n224), .ZN(n75) );
  INV_X4 U82 ( .A(n226), .ZN(n78) );
  INV_X4 U83 ( .A(n228), .ZN(n81) );
  INV_X4 U84 ( .A(n230), .ZN(n84) );
  INV_X4 U85 ( .A(n232), .ZN(n87) );
  INV_X4 U86 ( .A(n234), .ZN(n90) );
  INV_X4 U87 ( .A(n236), .ZN(n93) );
  INV_X4 U88 ( .A(n238), .ZN(n96) );
  INV_X4 U89 ( .A(n240), .ZN(n99) );
  INV_X4 U90 ( .A(n242), .ZN(n102) );
  INV_X4 U91 ( .A(n244), .ZN(n105) );
  INV_X4 U92 ( .A(n246), .ZN(n108) );
  INV_X4 U93 ( .A(n248), .ZN(n111) );
  INV_X4 U94 ( .A(n250), .ZN(n114) );
  INV_X4 U95 ( .A(n252), .ZN(n117) );
  INV_X4 U96 ( .A(n254), .ZN(n120) );
  INV_X4 U97 ( .A(n256), .ZN(n123) );
  INV_X4 U98 ( .A(n258), .ZN(n126) );
  NOR2_X1 U99 ( .A1(n261), .A2(n130), .ZN(n196) );
  INV_X1 U100 ( .A(aload[0]), .ZN(n130) );
  OAI21_X1 U101 ( .B1(arst), .B2(aload[0]), .A(rst), .ZN(n195) );
  NOR2_X1 U102 ( .A1(n260), .A2(n131), .ZN(n198) );
  INV_X1 U103 ( .A(aload[1]), .ZN(n131) );
  OAI21_X1 U104 ( .B1(arst), .B2(aload[1]), .A(rst), .ZN(n197) );
  NOR2_X1 U105 ( .A1(n262), .A2(n132), .ZN(n200) );
  INV_X1 U106 ( .A(aload[2]), .ZN(n132) );
  OAI21_X1 U107 ( .B1(arst), .B2(aload[2]), .A(rst), .ZN(n199) );
  NOR2_X1 U108 ( .A1(n261), .A2(n133), .ZN(n202) );
  INV_X1 U109 ( .A(aload[3]), .ZN(n133) );
  OAI21_X1 U110 ( .B1(arst), .B2(aload[3]), .A(rst), .ZN(n201) );
  NOR2_X1 U111 ( .A1(n260), .A2(n134), .ZN(n204) );
  INV_X1 U112 ( .A(aload[4]), .ZN(n134) );
  OAI21_X1 U113 ( .B1(arst), .B2(aload[4]), .A(rst), .ZN(n203) );
  NOR2_X1 U114 ( .A1(n262), .A2(n135), .ZN(n206) );
  INV_X1 U115 ( .A(aload[5]), .ZN(n135) );
  OAI21_X1 U116 ( .B1(arst), .B2(aload[5]), .A(rst), .ZN(n205) );
  NOR2_X1 U117 ( .A1(n261), .A2(n136), .ZN(n208) );
  INV_X1 U118 ( .A(aload[6]), .ZN(n136) );
  OAI21_X1 U119 ( .B1(arst), .B2(aload[6]), .A(rst), .ZN(n207) );
  NOR2_X1 U120 ( .A1(n260), .A2(n137), .ZN(n210) );
  INV_X1 U121 ( .A(aload[7]), .ZN(n137) );
  OAI21_X1 U122 ( .B1(arst), .B2(aload[7]), .A(rst), .ZN(n209) );
  NOR2_X1 U123 ( .A1(n262), .A2(n138), .ZN(n212) );
  INV_X1 U124 ( .A(aload[8]), .ZN(n138) );
  OAI21_X1 U125 ( .B1(arst), .B2(aload[8]), .A(rst), .ZN(n211) );
  NOR2_X1 U126 ( .A1(n261), .A2(n139), .ZN(n214) );
  INV_X1 U127 ( .A(aload[9]), .ZN(n139) );
  OAI21_X1 U128 ( .B1(arst), .B2(aload[9]), .A(rst), .ZN(n213) );
  NOR2_X1 U129 ( .A1(n260), .A2(n140), .ZN(n216) );
  INV_X1 U130 ( .A(aload[10]), .ZN(n140) );
  OAI21_X1 U131 ( .B1(arst), .B2(aload[10]), .A(rst), .ZN(n215) );
  NOR2_X1 U132 ( .A1(n262), .A2(n141), .ZN(n218) );
  INV_X1 U133 ( .A(aload[11]), .ZN(n141) );
  OAI21_X1 U134 ( .B1(arst), .B2(aload[11]), .A(rst), .ZN(n217) );
  NOR2_X1 U135 ( .A1(n261), .A2(n142), .ZN(n220) );
  INV_X1 U136 ( .A(aload[12]), .ZN(n142) );
  OAI21_X1 U137 ( .B1(arst), .B2(aload[12]), .A(rst), .ZN(n219) );
  NOR2_X1 U138 ( .A1(n260), .A2(n143), .ZN(n222) );
  INV_X1 U139 ( .A(aload[13]), .ZN(n143) );
  OAI21_X1 U140 ( .B1(arst), .B2(aload[13]), .A(rst), .ZN(n221) );
  NOR2_X1 U141 ( .A1(n262), .A2(n144), .ZN(n224) );
  INV_X1 U142 ( .A(aload[14]), .ZN(n144) );
  OAI21_X1 U143 ( .B1(arst), .B2(aload[14]), .A(rst), .ZN(n223) );
  NOR2_X1 U144 ( .A1(n261), .A2(n145), .ZN(n226) );
  INV_X1 U145 ( .A(aload[15]), .ZN(n145) );
  OAI21_X1 U146 ( .B1(arst), .B2(aload[15]), .A(rst), .ZN(n225) );
  NOR2_X1 U147 ( .A1(n260), .A2(n146), .ZN(n228) );
  INV_X1 U148 ( .A(aload[16]), .ZN(n146) );
  OAI21_X1 U149 ( .B1(arst), .B2(aload[16]), .A(rst), .ZN(n227) );
  NOR2_X1 U150 ( .A1(n262), .A2(n147), .ZN(n230) );
  INV_X1 U151 ( .A(aload[17]), .ZN(n147) );
  OAI21_X1 U152 ( .B1(arst), .B2(aload[17]), .A(rst), .ZN(n229) );
  NOR2_X1 U153 ( .A1(n261), .A2(n148), .ZN(n232) );
  INV_X1 U154 ( .A(aload[18]), .ZN(n148) );
  OAI21_X1 U155 ( .B1(arst), .B2(aload[18]), .A(rst), .ZN(n231) );
  NOR2_X1 U156 ( .A1(n260), .A2(n149), .ZN(n234) );
  INV_X1 U157 ( .A(aload[19]), .ZN(n149) );
  OAI21_X1 U158 ( .B1(arst), .B2(aload[19]), .A(rst), .ZN(n233) );
  NOR2_X1 U159 ( .A1(n262), .A2(n150), .ZN(n236) );
  INV_X1 U160 ( .A(aload[20]), .ZN(n150) );
  OAI21_X1 U161 ( .B1(arst), .B2(aload[20]), .A(rst), .ZN(n235) );
  NOR2_X1 U162 ( .A1(n261), .A2(n151), .ZN(n238) );
  INV_X1 U163 ( .A(aload[21]), .ZN(n151) );
  OAI21_X1 U164 ( .B1(arst), .B2(aload[21]), .A(rst), .ZN(n237) );
  NOR2_X1 U165 ( .A1(n260), .A2(n152), .ZN(n240) );
  INV_X1 U166 ( .A(aload[22]), .ZN(n152) );
  OAI21_X1 U167 ( .B1(arst), .B2(aload[22]), .A(rst), .ZN(n239) );
  NOR2_X1 U168 ( .A1(n262), .A2(n153), .ZN(n242) );
  INV_X1 U169 ( .A(aload[23]), .ZN(n153) );
  OAI21_X1 U170 ( .B1(arst), .B2(aload[23]), .A(rst), .ZN(n241) );
  NOR2_X1 U171 ( .A1(n261), .A2(n154), .ZN(n244) );
  INV_X1 U172 ( .A(aload[24]), .ZN(n154) );
  OAI21_X1 U173 ( .B1(arst), .B2(aload[24]), .A(rst), .ZN(n243) );
  NOR2_X1 U174 ( .A1(n260), .A2(n155), .ZN(n246) );
  INV_X1 U175 ( .A(aload[25]), .ZN(n155) );
  OAI21_X1 U176 ( .B1(arst), .B2(aload[25]), .A(rst), .ZN(n245) );
  NOR2_X1 U177 ( .A1(n262), .A2(n156), .ZN(n248) );
  INV_X1 U178 ( .A(aload[26]), .ZN(n156) );
  OAI21_X1 U179 ( .B1(arst), .B2(aload[26]), .A(rst), .ZN(n247) );
  NOR2_X1 U180 ( .A1(n261), .A2(n157), .ZN(n250) );
  INV_X1 U181 ( .A(aload[27]), .ZN(n157) );
  OAI21_X1 U182 ( .B1(arst), .B2(aload[27]), .A(rst), .ZN(n249) );
  NOR2_X1 U183 ( .A1(n260), .A2(n158), .ZN(n252) );
  INV_X1 U184 ( .A(aload[28]), .ZN(n158) );
  OAI21_X1 U185 ( .B1(arst), .B2(aload[28]), .A(rst), .ZN(n251) );
  NOR2_X1 U186 ( .A1(n262), .A2(n159), .ZN(n254) );
  INV_X1 U187 ( .A(aload[29]), .ZN(n159) );
  OAI21_X1 U188 ( .B1(arst), .B2(aload[29]), .A(rst), .ZN(n253) );
  NOR2_X1 U189 ( .A1(n261), .A2(n160), .ZN(n256) );
  INV_X1 U190 ( .A(aload[30]), .ZN(n160) );
  OAI21_X1 U191 ( .B1(arst), .B2(aload[30]), .A(rst), .ZN(n255) );
  NOR2_X1 U192 ( .A1(n260), .A2(n161), .ZN(n258) );
  INV_X1 U193 ( .A(aload[31]), .ZN(n161) );
  NAND2_X1 U194 ( .A1(rst), .A2(n162), .ZN(n129) );
  INV_X1 U195 ( .A(arst), .ZN(n162) );
  OAI21_X1 U196 ( .B1(arst), .B2(aload[31]), .A(rst), .ZN(n257) );
  INV_X4 U197 ( .A(n257), .ZN(n163) );
  INV_X4 U198 ( .A(n255), .ZN(n164) );
  INV_X4 U199 ( .A(n253), .ZN(n165) );
  INV_X4 U200 ( .A(n251), .ZN(n166) );
  INV_X4 U201 ( .A(n249), .ZN(n167) );
  INV_X4 U202 ( .A(n247), .ZN(n168) );
  INV_X4 U203 ( .A(n245), .ZN(n169) );
  INV_X4 U204 ( .A(n243), .ZN(n170) );
  INV_X4 U205 ( .A(n241), .ZN(n171) );
  INV_X4 U206 ( .A(n239), .ZN(n172) );
  INV_X4 U207 ( .A(n237), .ZN(n173) );
  INV_X4 U208 ( .A(n235), .ZN(n174) );
  INV_X4 U209 ( .A(n233), .ZN(n175) );
  INV_X4 U210 ( .A(n231), .ZN(n176) );
  INV_X4 U211 ( .A(n229), .ZN(n177) );
  INV_X4 U212 ( .A(n227), .ZN(n178) );
  INV_X4 U213 ( .A(n225), .ZN(n179) );
  INV_X4 U214 ( .A(n223), .ZN(n180) );
  INV_X4 U215 ( .A(n221), .ZN(n181) );
  INV_X4 U216 ( .A(n219), .ZN(n182) );
  INV_X4 U217 ( .A(n217), .ZN(n183) );
  INV_X4 U218 ( .A(n215), .ZN(n184) );
  INV_X4 U219 ( .A(n213), .ZN(n185) );
  INV_X4 U220 ( .A(n211), .ZN(n186) );
  INV_X4 U221 ( .A(n209), .ZN(n187) );
  INV_X4 U222 ( .A(n207), .ZN(n188) );
  INV_X4 U223 ( .A(n205), .ZN(n189) );
  INV_X4 U224 ( .A(n203), .ZN(n190) );
  INV_X4 U225 ( .A(n201), .ZN(n191) );
  INV_X4 U226 ( .A(n199), .ZN(n192) );
  INV_X4 U227 ( .A(n197), .ZN(n193) );
  INV_X4 U228 ( .A(n195), .ZN(n194) );
  INV_X1 U229 ( .A(n129), .ZN(n259) );
  INV_X1 U230 ( .A(n259), .ZN(n260) );
  INV_X1 U231 ( .A(n259), .ZN(n261) );
  INV_X1 U232 ( .A(n259), .ZN(n262) );
endmodule

