`define R0 32'b0
