
module pipeline ( clk, rst, initPC, instruction, iAddr, memInstr, memAddr, 
        memRdData, memWrData, dSize, memWr, busA, busB, busFP, rs1, rs2, rd, 
        regWrData, regWr, fp );
  input [31:0] initPC;
  input [31:0] instruction;
  output [31:0] iAddr;
  output [31:0] memInstr;
  output [31:0] memAddr;
  input [31:0] memRdData;
  output [31:0] memWrData;
  output [1:0] dSize;
  input [31:0] busA;
  input [31:0] busB;
  input [31:0] busFP;
  output [4:0] rs1;
  output [4:0] rs2;
  output [4:0] rd;
  output [31:0] regWrData;
  input clk, rst;
  output memWr, regWr, fp;
  wire   not_trap_3, op0_1, valid_2, valid_3, setInv_2, op0_2, zeroExt_2,
         not_trap_2, op0_3, hazard_detect_multiplier_fsm_N19,
         hazard_detect_multiplier_fsm_N18, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3577, n3578, n3579, n3580, n3581, n3583, n3584, n3586,
         n3587, n3589, n3590, n3591, n3592, n3593, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3607, n3608, n3609,
         n3610, n3611, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3712,
         n3714, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3724, n3726,
         n3728, n3729, n3730, n3731, n3732, n3734, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3963, n3965, n3966, n3970, n3971,
         n3972, n3975, n3976, n3978, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196;
  wire   [4:0] rd_2;
  wire   [4:0] rd_3;
  wire   [31:0] aluRes_2;
  wire   [1:0] reg31Val_3;
  wire   [31:0] reg31Val_0;
  wire   [31:0] wb_dsize_reg_z2;
  wire   [28:8] ex_multing_set_product_in_sig_z1;

  DFFR_X1 ex_mem_product_in_q_reg_0_ ( .D(aluRes_2[0]), .CK(clk), .RN(n4846), 
        .Q(n4590) );
  DFFR_X1 ex_mem_product_in_q_reg_24_ ( .D(aluRes_2[24]), .CK(clk), .RN(n4854), 
        .Q(ex_multing_set_product_in_sig_z1[24]) );
  DFFR_X1 ex_mem_product_in_q_reg_31_ ( .D(aluRes_2[31]), .CK(clk), .RN(n4849), 
        .Q(n4588) );
  DFFR_X1 ex_mem_product_in_q_reg_7_ ( .D(n4451), .CK(clk), .RN(n4852), .QN(
        n7574) );
  DFFR_X1 ex_mem_product_in_q_reg_23_ ( .D(aluRes_2[23]), .CK(clk), .RN(n4855), 
        .Q(n4571) );
  DFFR_X1 ex_mem_product_in_q_reg_26_ ( .D(aluRes_2[26]), .CK(clk), .RN(n4850), 
        .Q(ex_multing_set_product_in_sig_z1[26]) );
  DFFR_X1 ex_mem_product_in_q_reg_11_ ( .D(n9180), .CK(clk), .RN(n4858), .Q(
        n4460) );
  DFFR_X1 ex_mem_product_in_q_reg_28_ ( .D(aluRes_2[28]), .CK(clk), .RN(n4853), 
        .Q(ex_multing_set_product_in_sig_z1[28]) );
  DFFR_X1 ex_mem_product_in_q_reg_13_ ( .D(n9182), .CK(clk), .RN(n4859), .Q(
        n4461) );
  DFFR_X1 ex_mem_product_in_q_reg_30_ ( .D(aluRes_2[30]), .CK(clk), .RN(n4851), 
        .Q(n4573) );
  DFFR_X1 ex_mem_product_in_q_reg_15_ ( .D(aluRes_2[15]), .CK(clk), .RN(n4840), 
        .Q(n4580) );
  DFFR_X1 ex_mem_product_in_q_reg_16_ ( .D(aluRes_2[16]), .CK(clk), .RN(n4840), 
        .Q(n4561) );
  DFFR_X1 ex_mem_product_in_q_reg_10_ ( .D(n9185), .CK(clk), .RN(n4840), .Q(
        ex_multing_set_product_in_sig_z1[10]) );
  DFFR_X1 ex_mem_product_in_q_reg_1_ ( .D(n9186), .CK(clk), .RN(n4840), .Q(
        n4589) );
  DFFR_X1 ex_mem_product_in_q_reg_20_ ( .D(aluRes_2[20]), .CK(clk), .RN(n4840), 
        .Q(ex_multing_set_product_in_sig_z1[20]) );
  DFFR_X1 hazard_detect_multiplier_fsm_cur_state_reg_0_ ( .D(n9187), .CK(clk), 
        .RN(n4840), .Q(n4537), .QN(n7573) );
  DFFR_X1 hazard_detect_multiplier_fsm_cur_state_reg_1_ ( .D(
        hazard_detect_multiplier_fsm_N18), .CK(clk), .RN(n4840), .Q(n4135), 
        .QN(n7572) );
  DFFR_X1 ex_mem_product_in_q_reg_21_ ( .D(aluRes_2[21]), .CK(clk), .RN(n4840), 
        .Q(n4581) );
  DFFR_X1 ex_mem_product_in_q_reg_22_ ( .D(aluRes_2[22]), .CK(clk), .RN(n4840), 
        .Q(ex_multing_set_product_in_sig_z1[22]) );
  DFFR_X1 ex_mem_product_in_q_reg_9_ ( .D(n9188), .CK(clk), .RN(n4840), .Q(
        n4455), .QN(n7571) );
  DFFR_X1 ex_mem_product_in_q_reg_17_ ( .D(n9183), .CK(clk), .RN(n4840), .Q(
        n4570) );
  DFFR_X1 ex_mem_product_in_q_reg_12_ ( .D(n9181), .CK(clk), .RN(n4840), .Q(
        ex_multing_set_product_in_sig_z1[12]) );
  DFFR_X1 ex_mem_product_in_q_reg_29_ ( .D(aluRes_2[29]), .CK(clk), .RN(n4839), 
        .Q(n4584) );
  DFFR_X1 ex_mem_product_in_q_reg_8_ ( .D(n9189), .CK(clk), .RN(n4839), .Q(
        ex_multing_set_product_in_sig_z1[8]) );
  DFFR_X1 ex_mem_product_in_q_reg_25_ ( .D(aluRes_2[25]), .CK(clk), .RN(n4839), 
        .Q(n4572) );
  DFFR_X1 ex_mem_product_in_q_reg_18_ ( .D(aluRes_2[18]), .CK(clk), .RN(n4839), 
        .Q(ex_multing_set_product_in_sig_z1[18]) );
  DFFR_X1 ex_mem_product_in_q_reg_27_ ( .D(aluRes_2[27]), .CK(clk), .RN(n4839), 
        .Q(n4583) );
  DFFR_X1 ex_mem_product_in_q_reg_4_ ( .D(n9192), .CK(clk), .RN(n4839), .QN(
        n7570) );
  DFFR_X1 ex_mem_product_in_q_reg_19_ ( .D(aluRes_2[19]), .CK(clk), .RN(n4839), 
        .Q(n4582) );
  DFFR_X1 ex_mem_product_in_q_reg_2_ ( .D(n9194), .CK(clk), .RN(n4839), .QN(
        n7569) );
  DFFR_X1 ex_mem_product_in_q_reg_5_ ( .D(n9191), .CK(clk), .RN(n4839), .QN(
        n7568) );
  DFFR_X1 ex_mem_product_in_q_reg_6_ ( .D(n9190), .CK(clk), .RN(n4839), .QN(
        n7567) );
  DFFR_X1 ex_mem_product_in_q_reg_14_ ( .D(n9184), .CK(clk), .RN(n4839), .Q(
        n4493) );
  DFFR_X1 ex_mem_product_in_q_reg_3_ ( .D(n9193), .CK(clk), .RN(n4839), .QN(
        n7566) );
  DFFR_X1 ex_mem_aluRes_q_reg_0_ ( .D(n3978), .CK(clk), .RN(n4858), .Q(
        memAddr[0]), .QN(n9055) );
  DFFR_X1 ex_mem_aluRes_q_reg_24_ ( .D(n9163), .CK(clk), .RN(n4857), .Q(
        memAddr[24]), .QN(n9034) );
  DFFR_X1 ex_mem_aluRes_q_reg_31_ ( .D(n3976), .CK(clk), .RN(n4857), .Q(
        memAddr[31]), .QN(n8988) );
  DFFR_X1 ex_mem_aluRes_q_reg_7_ ( .D(n3975), .CK(clk), .RN(n4859), .Q(
        memAddr[7]), .QN(n9000) );
  DFFR_X1 ex_mem_aluRes_q_reg_23_ ( .D(n9162), .CK(clk), .RN(n4859), .Q(
        memAddr[23]), .QN(n9031) );
  DFFR_X1 ex_mem_aluRes_q_reg_26_ ( .D(n9165), .CK(clk), .RN(n4857), .Q(
        memAddr[26]), .QN(n9039) );
  DFFR_X1 ex_mem_aluRes_q_reg_11_ ( .D(n3972), .CK(clk), .RN(n4858), .Q(
        memAddr[11]), .QN(n9007) );
  DFFR_X1 ex_mem_aluRes_q_reg_28_ ( .D(n3971), .CK(clk), .RN(n4857), .Q(
        memAddr[28]), .QN(n9043) );
  DFFR_X1 ex_mem_aluRes_q_reg_13_ ( .D(n3970), .CK(clk), .RN(n4858), .Q(
        memAddr[13]), .QN(n9009) );
  DFFR_X1 ex_mem_aluRes_q_reg_30_ ( .D(n9168), .CK(clk), .RN(n4859), .Q(
        memAddr[30]), .QN(n9049) );
  DFFR_X1 ex_mem_aluRes_q_reg_15_ ( .D(n9155), .CK(clk), .RN(n4858), .Q(
        memAddr[15]), .QN(n9013) );
  DFFR_X1 ex_mem_aluRes_q_reg_16_ ( .D(n9156), .CK(clk), .RN(n4858), .Q(
        memAddr[16]), .QN(n9016) );
  DFFR_X1 ex_mem_aluRes_q_reg_10_ ( .D(n3966), .CK(clk), .RN(n4858), .Q(
        memAddr[10]), .QN(n9006) );
  DFFR_X1 ex_mem_aluRes_q_reg_1_ ( .D(n3965), .CK(clk), .RN(n4858), .Q(
        memAddr[1]), .QN(n8989) );
  DFFR_X1 ex_mem_aluRes_q_reg_20_ ( .D(n9159), .CK(clk), .RN(n4857), .Q(
        memAddr[20]), .QN(n9024) );
  DFFR_X1 ex_mem_isZero_q_reg ( .D(n3963), .CK(clk), .RN(n4850), .Q(n4388), 
        .QN(n8846) );
  DFFR_X1 id_ex_busA_q_reg_0_ ( .D(n9122), .CK(clk), .RN(n4866), .Q(n4372) );
  DFFR_X1 id_ex_busA_q_reg_1_ ( .D(n9121), .CK(clk), .RN(n4849), .Q(n4371) );
  DFFR_X1 id_ex_busA_q_reg_2_ ( .D(n9120), .CK(clk), .RN(n4867), .Q(n4336), 
        .QN(n8982) );
  DFFR_X1 id_ex_busA_q_reg_3_ ( .D(n9119), .CK(clk), .RN(n4848), .Q(n4340), 
        .QN(n8981) );
  DFFR_X1 id_ex_busA_q_reg_4_ ( .D(n9118), .CK(clk), .RN(n4867), .Q(n4335), 
        .QN(n8980) );
  DFFR_X1 id_ex_busA_q_reg_5_ ( .D(n9117), .CK(clk), .RN(n4848), .Q(n4337), 
        .QN(n8979) );
  DFFR_X1 id_ex_busA_q_reg_6_ ( .D(n9116), .CK(clk), .RN(n4867), .Q(n4338), 
        .QN(n8978) );
  DFFR_X1 id_ex_busA_q_reg_7_ ( .D(n9115), .CK(clk), .RN(n4848), .Q(n4206) );
  DFFR_X1 id_ex_busA_q_reg_8_ ( .D(n9114), .CK(clk), .RN(n4867), .Q(n4560), 
        .QN(n8977) );
  DFFR_X1 id_ex_busA_q_reg_9_ ( .D(n9113), .CK(clk), .RN(n4848), .Q(n4559), 
        .QN(n8976) );
  DFFR_X1 id_ex_busA_q_reg_10_ ( .D(n9112), .CK(clk), .RN(n4849), .Q(n4209) );
  DFFR_X1 id_ex_busA_q_reg_11_ ( .D(n9111), .CK(clk), .RN(n4866), .Q(n4207) );
  DFFR_X1 id_ex_busA_q_reg_12_ ( .D(n9110), .CK(clk), .RN(n4849), .Q(n4334), 
        .QN(n8984) );
  DFFR_X1 id_ex_busA_q_reg_13_ ( .D(n9109), .CK(clk), .RN(n4866), .Q(n4208) );
  DFFR_X1 id_ex_busA_q_reg_14_ ( .D(n9108), .CK(clk), .RN(n4849), .Q(n4339), 
        .QN(n8983) );
  DFFR_X1 id_ex_busA_q_reg_15_ ( .D(n9107), .CK(clk), .RN(n4866), .Q(n4418) );
  DFFR_X1 id_ex_busA_q_reg_16_ ( .D(n9106), .CK(clk), .RN(n4849), .Q(n4659), 
        .QN(n8952) );
  DFFR_X1 id_ex_busA_q_reg_17_ ( .D(n9105), .CK(clk), .RN(n4866), .Q(n4665), 
        .QN(n8951) );
  DFFR_X1 id_ex_busA_q_reg_18_ ( .D(n9104), .CK(clk), .RN(n4849), .Q(n4568), 
        .QN(n8950) );
  DFFR_X1 id_ex_busA_q_reg_19_ ( .D(n9103), .CK(clk), .RN(n4866), .Q(n4662), 
        .QN(n8949) );
  DFFR_X1 id_ex_busA_q_reg_20_ ( .D(n9102), .CK(clk), .RN(n4866), .Q(n4417) );
  DFFR_X1 id_ex_busA_q_reg_21_ ( .D(n9101), .CK(clk), .RN(n4849), .Q(n4667), 
        .QN(n8948) );
  DFFR_X1 id_ex_busA_q_reg_22_ ( .D(n9100), .CK(clk), .RN(n4867), .Q(n4666), 
        .QN(n8947) );
  DFFR_X1 id_ex_busA_q_reg_23_ ( .D(n9099), .CK(clk), .RN(n4849), .Q(n4656), 
        .QN(n9030) );
  DFFR_X1 id_ex_busA_q_reg_24_ ( .D(n9098), .CK(clk), .RN(n4867), .Q(n4657), 
        .QN(n9033) );
  DFFR_X1 id_ex_busA_q_reg_25_ ( .D(n9097), .CK(clk), .RN(n4848), .Q(n4664), 
        .QN(n9036) );
  DFFR_X1 id_ex_busA_q_reg_26_ ( .D(n9096), .CK(clk), .RN(n4867), .Q(n4475) );
  DFFR_X1 id_ex_busA_q_reg_27_ ( .D(n9095), .CK(clk), .RN(n4848), .Q(n4663), 
        .QN(n8946) );
  DFFR_X1 id_ex_busA_q_reg_28_ ( .D(n9094), .CK(clk), .RN(n4867), .Q(n4711) );
  DFFR_X1 id_ex_busA_q_reg_29_ ( .D(n9093), .CK(clk), .RN(n4848), .Q(n4714) );
  DFFR_X1 id_ex_busA_q_reg_30_ ( .D(n9092), .CK(clk), .RN(n4848), .Q(n4712) );
  DFFR_X1 id_ex_busA_q_reg_31_ ( .D(n9091), .CK(clk), .RN(n4867), .Q(n4474) );
  DFFR_X1 id_ex_busB_q_reg_0_ ( .D(n9154), .CK(clk), .RN(n4867), .Q(n4348), 
        .QN(n9056) );
  DFFR_X1 id_ex_busB_q_reg_1_ ( .D(n9153), .CK(clk), .RN(n4847), .Q(n4347), 
        .QN(n8990) );
  DFFR_X1 id_ex_busB_q_reg_2_ ( .D(n9152), .CK(clk), .RN(n4868), .Q(n4661), 
        .QN(n8992) );
  DFFR_X1 id_ex_busB_q_reg_3_ ( .D(n9151), .CK(clk), .RN(n4847), .Q(n4658), 
        .QN(n8994) );
  DFFR_X1 id_ex_busB_q_reg_4_ ( .D(n9150), .CK(clk), .RN(n4868), .Q(n4713) );
  DFFR_X1 id_ex_busB_q_reg_5_ ( .D(n9149), .CK(clk), .RN(n4847), .Q(n4660), 
        .QN(n8997) );
  DFFR_X1 id_ex_busB_q_reg_6_ ( .D(n9148), .CK(clk), .RN(n4869), .Q(n4655), 
        .QN(n8999) );
  DFFR_X1 id_ex_busB_q_reg_7_ ( .D(n9147), .CK(clk), .RN(n4847), .Q(n4668), 
        .QN(n9001) );
  DFFR_X1 id_ex_busB_q_reg_8_ ( .D(n9146), .CK(clk), .RN(n4869), .Q(n4346), 
        .QN(n9003) );
  DFFR_X1 id_ex_busB_q_reg_9_ ( .D(n9145), .CK(clk), .RN(n4846), .Q(n4345), 
        .QN(n9005) );
  DFFR_X1 id_ex_busB_q_reg_10_ ( .D(n9144), .CK(clk), .RN(n4848), .Q(n4704) );
  DFFR_X1 id_ex_busB_q_reg_11_ ( .D(n9143), .CK(clk), .RN(n4867), .Q(n4715) );
  DFFR_X1 id_ex_busB_q_reg_12_ ( .D(n9142), .CK(clk), .RN(n4848), .Q(n4707) );
  DFFR_X1 id_ex_busB_q_reg_13_ ( .D(n9141), .CK(clk), .RN(n4868), .Q(n4669), 
        .QN(n9010) );
  DFFR_X1 id_ex_busB_q_reg_14_ ( .D(n9140), .CK(clk), .RN(n4848), .Q(n4671), 
        .QN(n9012) );
  DFFR_X1 id_ex_busB_q_reg_15_ ( .D(n9139), .CK(clk), .RN(n4868), .Q(n4652), 
        .QN(n9014) );
  DFFR_X1 id_ex_busB_q_reg_16_ ( .D(n9138), .CK(clk), .RN(n4847), .Q(n4344), 
        .QN(n9015) );
  DFFR_X1 id_ex_busB_q_reg_17_ ( .D(n9137), .CK(clk), .RN(n4868), .Q(n4343), 
        .QN(n9017) );
  DFFR_X1 id_ex_busB_q_reg_18_ ( .D(n9136), .CK(clk), .RN(n4847), .Q(n4708), 
        .QN(n9019) );
  DFFR_X1 id_ex_busB_q_reg_19_ ( .D(n9135), .CK(clk), .RN(n4868), .Q(n4710), 
        .QN(n9021) );
  DFFR_X1 id_ex_busB_q_reg_20_ ( .D(n9134), .CK(clk), .RN(n4868), .Q(n4653), 
        .QN(n9023) );
  DFFR_X1 id_ex_busB_q_reg_21_ ( .D(n9133), .CK(clk), .RN(n4847), .Q(n4705), 
        .QN(n9025) );
  DFFR_X1 id_ex_busB_q_reg_22_ ( .D(n9132), .CK(clk), .RN(n4868), .Q(n4706), 
        .QN(n9027) );
  DFFR_X1 id_ex_busB_q_reg_23_ ( .D(n9131), .CK(clk), .RN(n4847), .Q(n4333), 
        .QN(n9029) );
  DFFR_X1 id_ex_busB_q_reg_24_ ( .D(n9130), .CK(clk), .RN(n4868), .Q(n4342), 
        .QN(n9032) );
  DFFR_X1 id_ex_busB_q_reg_25_ ( .D(n9129), .CK(clk), .RN(n4847), .Q(n4341), 
        .QN(n9035) );
  DFFR_X1 id_ex_busB_q_reg_26_ ( .D(n9128), .CK(clk), .RN(n4868), .Q(n4553), 
        .QN(n9038) );
  DFFR_X1 id_ex_busB_q_reg_27_ ( .D(n9127), .CK(clk), .RN(n4847), .Q(n4709), 
        .QN(n9040) );
  DFFR_X1 id_ex_busB_q_reg_28_ ( .D(n9126), .CK(clk), .RN(n4868), .Q(n4552), 
        .QN(n9042) );
  DFFR_X1 id_ex_busB_q_reg_29_ ( .D(n9125), .CK(clk), .RN(n4847), .Q(n4654), 
        .QN(n9044) );
  DFFR_X1 id_ex_busB_q_reg_30_ ( .D(n9124), .CK(clk), .RN(n4847), .Q(n4551), 
        .QN(n9046) );
  DFFR_X1 id_ex_busB_q_reg_31_ ( .D(n9123), .CK(clk), .RN(n4868), .Q(n4550), 
        .QN(n8987) );
  DFFR_X1 id_ex_aluCtrl_q_reg_2_ ( .D(n3898), .CK(clk), .RN(n4866), .Q(n4545), 
        .QN(n9050) );
  DFFR_X1 if_id_instr_q_reg_31_ ( .D(n3893), .CK(clk), .RN(n4841), .Q(n4275), 
        .QN(n8958) );
  DFFR_X1 if_id_instr_q_reg_29_ ( .D(n3891), .CK(clk), .RN(n4876), .Q(n4119), 
        .QN(n8953) );
  DFFR_X1 id_ex_memRd_q_reg ( .D(n3890), .CK(clk), .RN(n4873), .QN(n8845) );
  DFFR_X1 if_id_instr_q_reg_28_ ( .D(n3889), .CK(clk), .RN(n4841), .Q(n4538), 
        .QN(n8957) );
  DFFR_X1 if_id_instr_q_reg_27_ ( .D(n3888), .CK(clk), .RN(n4876), .Q(n4120), 
        .QN(n8954) );
  DFFR_X1 id_ex_branch_q_reg ( .D(n3887), .CK(clk), .RN(n4849), .Q(n4629), 
        .QN(n8844) );
  DFFR_X1 id_ex_jr_q_reg ( .D(n3886), .CK(clk), .RN(n4856), .Q(n4630), .QN(
        n8843) );
  DFFR_X1 id_ex_op0_q_reg ( .D(n9178), .CK(clk), .RN(n4876), .Q(op0_2) );
  DFFR_X1 id_ex_link_q_reg ( .D(n9179), .CK(clk), .RN(n4857), .Q(n4628), .QN(
        n8932) );
  DFFR_X1 id_ex_dSize_q_reg_1_ ( .D(n3882), .CK(clk), .RN(n4846), .Q(n4634), 
        .QN(n8842) );
  DFFR_X1 id_ex_dSize_q_reg_0_ ( .D(n3881), .CK(clk), .RN(n4869), .Q(n4633), 
        .QN(n8841) );
  DFFR_X1 id_ex_imm32_q_reg_4_ ( .D(n3880), .CK(clk), .RN(n4845), .Q(n4370), 
        .QN(n8964) );
  DFFR_X1 id_ex_imm32_q_reg_2_ ( .D(n3879), .CK(clk), .RN(n4845), .QN(n8840)
         );
  DFFR_X1 id_ex_imm32_q_reg_0_ ( .D(n3878), .CK(clk), .RN(n4846), .QN(n8839)
         );
  DFFR_X1 id_ex_jump_q_reg ( .D(n3877), .CK(clk), .RN(n4873), .QN(n8838) );
  DFFR_X1 id_ex_aluSrc_q_reg ( .D(n3876), .CK(clk), .RN(n4866), .Q(n4452), 
        .QN(n9054) );
  DFFR_X1 if_id_instr_q_reg_25_ ( .D(n3875), .CK(clk), .RN(n4876), .Q(rs1[4]), 
        .QN(n4528) );
  DFFR_X1 if_id_instr_q_reg_24_ ( .D(n3874), .CK(clk), .RN(n4841), .Q(rs1[3]), 
        .QN(n4529) );
  DFFR_X1 if_id_instr_q_reg_23_ ( .D(n3873), .CK(clk), .RN(n4876), .Q(rs1[2]), 
        .QN(n4527) );
  DFFR_X1 if_id_instr_q_reg_22_ ( .D(n3872), .CK(clk), .RN(n4841), .Q(rs1[1]), 
        .QN(n4531) );
  DFFR_X1 if_id_instr_q_reg_21_ ( .D(n3871), .CK(clk), .RN(n4875), .Q(rs1[0]), 
        .QN(n4530) );
  DFFR_X1 if_id_instr_q_reg_20_ ( .D(n3870), .CK(clk), .RN(n4841), .Q(n4332), 
        .QN(n8904) );
  DFFR_X1 if_id_instr_q_reg_19_ ( .D(n3869), .CK(clk), .RN(n4841), .Q(n4548), 
        .QN(n8905) );
  DFFR_X1 if_id_instr_q_reg_18_ ( .D(n3868), .CK(clk), .RN(n4875), .Q(n4547), 
        .QN(n8906) );
  DFFR_X1 if_id_instr_q_reg_17_ ( .D(n3867), .CK(clk), .RN(n4841), .Q(n4328), 
        .QN(n8907) );
  DFFR_X1 if_id_instr_q_reg_16_ ( .D(n3866), .CK(clk), .RN(n4875), .Q(n4329), 
        .QN(n8908) );
  DFFR_X1 if_id_instr_q_reg_15_ ( .D(n3865), .CK(clk), .RN(n4841), .Q(n4546), 
        .QN(n8945) );
  DFFR_X1 id_ex_imm32_q_reg_15_ ( .D(n3864), .CK(clk), .RN(n4846), .QN(n8837)
         );
  DFFR_X1 id_ex_imm32_q_reg_31_ ( .D(n3863), .CK(clk), .RN(n4845), .QN(n8836)
         );
  DFFR_X1 id_ex_imm32_q_reg_20_ ( .D(n3862), .CK(clk), .RN(n4846), .Q(n4557), 
        .QN(n8970) );
  DFFR_X1 id_ex_imm32_q_reg_18_ ( .D(n3861), .CK(clk), .RN(n4869), .Q(n4138), 
        .QN(n8972) );
  DFFR_X1 id_ex_imm32_q_reg_16_ ( .D(n3860), .CK(clk), .RN(n4869), .Q(n4564), 
        .QN(n8974) );
  DFFR_X1 if_id_instr_q_reg_14_ ( .D(n3859), .CK(clk), .RN(n4875), .QN(n8835)
         );
  DFFR_X1 id_ex_imm32_q_reg_30_ ( .D(n3858), .CK(clk), .RN(n4870), .QN(n8834)
         );
  DFFR_X1 id_ex_imm32_q_reg_14_ ( .D(n3857), .CK(clk), .RN(n4869), .QN(n8833)
         );
  DFFR_X1 if_id_instr_q_reg_13_ ( .D(n3856), .CK(clk), .RN(n4841), .QN(n8832)
         );
  DFFR_X1 id_ex_imm32_q_reg_29_ ( .D(n3855), .CK(clk), .RN(n4870), .QN(n8831)
         );
  DFFR_X1 id_ex_imm32_q_reg_13_ ( .D(n3854), .CK(clk), .RN(n4846), .QN(n8830)
         );
  DFFR_X1 if_id_instr_q_reg_12_ ( .D(n3853), .CK(clk), .RN(n4875), .QN(n8829)
         );
  DFFR_X1 id_ex_imm32_q_reg_28_ ( .D(n3852), .CK(clk), .RN(n4845), .QN(n8966)
         );
  DFFR_X1 id_ex_imm32_q_reg_12_ ( .D(n3851), .CK(clk), .RN(n4869), .Q(n4413), 
        .QN(n8828) );
  DFFR_X1 if_id_instr_q_reg_11_ ( .D(n3850), .CK(clk), .RN(n4841), .QN(n8827)
         );
  DFFR_X1 id_ex_imm32_q_reg_27_ ( .D(n3849), .CK(clk), .RN(n4870), .Q(n4177), 
        .QN(n8826) );
  DFFR_X1 id_ex_imm32_q_reg_11_ ( .D(n3848), .CK(clk), .RN(n4846), .Q(n4414), 
        .QN(n8825) );
  DFFR_X1 if_id_instr_q_reg_10_ ( .D(n3847), .CK(clk), .RN(n4875), .QN(n8824)
         );
  DFFR_X1 id_ex_imm32_q_reg_26_ ( .D(n3846), .CK(clk), .RN(n4845), .QN(n8968)
         );
  DFFR_X1 id_ex_imm32_q_reg_10_ ( .D(n3845), .CK(clk), .RN(n4869), .Q(n4415), 
        .QN(n8823) );
  DFFR_X1 if_id_instr_q_reg_9_ ( .D(n3844), .CK(clk), .RN(n4876), .QN(n8934)
         );
  DFFR_X1 id_ex_imm32_q_reg_9_ ( .D(n3843), .CK(clk), .RN(n4870), .QN(n8822)
         );
  DFFR_X1 id_ex_imm32_q_reg_25_ ( .D(n3842), .CK(clk), .RN(n4870), .Q(n4565), 
        .QN(n8933) );
  DFFR_X1 if_id_instr_q_reg_8_ ( .D(n3841), .CK(clk), .RN(n4847), .QN(n8936)
         );
  DFFR_X1 id_ex_imm32_q_reg_8_ ( .D(n3840), .CK(clk), .RN(n4845), .QN(n8960)
         );
  DFFR_X1 id_ex_imm32_q_reg_24_ ( .D(n3839), .CK(clk), .RN(n4846), .Q(n4566), 
        .QN(n8935) );
  DFFR_X1 if_id_instr_q_reg_7_ ( .D(n3838), .CK(clk), .RN(n4876), .QN(n8938)
         );
  DFFR_X1 id_ex_imm32_q_reg_7_ ( .D(n3837), .CK(clk), .RN(n4870), .QN(n8821)
         );
  DFFR_X1 id_ex_imm32_q_reg_23_ ( .D(n3836), .CK(clk), .RN(n4870), .Q(n4467), 
        .QN(n8937) );
  DFFR_X1 if_id_instr_q_reg_6_ ( .D(n3835), .CK(clk), .RN(n4848), .QN(n8940)
         );
  DFFR_X1 id_ex_imm32_q_reg_6_ ( .D(n3834), .CK(clk), .RN(n4845), .QN(n8962)
         );
  DFFR_X1 id_ex_imm32_q_reg_22_ ( .D(n3833), .CK(clk), .RN(n4846), .Q(n4407), 
        .QN(n8939) );
  DFFR_X1 if_id_instr_q_reg_5_ ( .D(n3832), .CK(clk), .RN(n4876), .Q(n4525), 
        .QN(n8956) );
  DFFR_X1 id_ex_imm32_q_reg_5_ ( .D(n3831), .CK(clk), .RN(n4870), .QN(n8820)
         );
  DFFR_X1 id_ex_imm32_q_reg_21_ ( .D(n3830), .CK(clk), .RN(n4869), .Q(n4175), 
        .QN(n8941) );
  DFFR_X1 if_id_instr_q_reg_3_ ( .D(n3828), .CK(clk), .RN(n4876), .Q(n4318), 
        .QN(n8955) );
  DFFR_X1 id_ex_imm32_q_reg_3_ ( .D(n3827), .CK(clk), .RN(n4870), .QN(n8819)
         );
  DFFR_X1 id_ex_imm32_q_reg_19_ ( .D(n3826), .CK(clk), .RN(n4846), .Q(n4176), 
        .QN(n8942) );
  DFFR_X1 id_ex_aluCtrl_q_reg_3_ ( .D(n3825), .CK(clk), .RN(n4849), .Q(n4133), 
        .QN(n9047) );
  DFFR_X1 if_id_instr_q_reg_1_ ( .D(n3824), .CK(clk), .RN(n4875), .Q(n4524), 
        .QN(n8944) );
  DFFR_X1 id_ex_imm32_q_reg_1_ ( .D(n3823), .CK(clk), .RN(n4869), .QN(n8818)
         );
  DFFR_X1 id_ex_imm32_q_reg_17_ ( .D(n3822), .CK(clk), .RN(n4846), .Q(n4567), 
        .QN(n8943) );
  DFFR_X1 id_ex_aluCtrl_q_reg_1_ ( .D(n3821), .CK(clk), .RN(n4849), .Q(n4136), 
        .QN(n9051) );
  DFFR_X1 id_ex_setInv_q_reg ( .D(n3820), .CK(clk), .RN(n4873), .Q(setInv_2)
         );
  DFFR_X1 id_ex_rd_q_reg_4_ ( .D(n3819), .CK(clk), .RN(n4873), .Q(rd_2[4]), 
        .QN(n4533) );
  DFFR_X1 id_ex_rd_q_reg_3_ ( .D(n3818), .CK(clk), .RN(n4841), .Q(rd_2[3]), 
        .QN(n4324) );
  DFFR_X1 id_ex_rd_q_reg_2_ ( .D(n3817), .CK(clk), .RN(n4873), .Q(rd_2[2]), 
        .QN(n4095) );
  DFFR_X1 id_ex_rd_q_reg_1_ ( .D(n3816), .CK(clk), .RN(n4877), .Q(rd_2[1]), 
        .QN(n4322) );
  DFFR_X1 id_ex_rd_q_reg_0_ ( .D(n3815), .CK(clk), .RN(n4873), .Q(rd_2[0]), 
        .QN(n4094) );
  DFFR_X1 id_ex_aluCtrl_q_reg_0_ ( .D(n3814), .CK(clk), .RN(n4866), .Q(n4121), 
        .QN(n9048) );
  DFFR_X1 ex_mem_fp_q_reg ( .D(n3763), .CK(clk), .RN(n4862), .Q(n4627), .QN(
        n8817) );
  DFFR_X1 ex_mem_rd_q_reg_0_ ( .D(n3761), .CK(clk), .RN(n4850), .Q(rd_3[0]), 
        .QN(n4319) );
  DFFR_X1 ex_mem_rd_q_reg_1_ ( .D(n3759), .CK(clk), .RN(n4865), .Q(rd_3[1]), 
        .QN(n4093) );
  DFFR_X1 ex_mem_rd_q_reg_2_ ( .D(n3757), .CK(clk), .RN(n4850), .Q(rd_3[2]), 
        .QN(n4081) );
  DFFR_X1 ex_mem_busA_q_reg_31_ ( .D(n3755), .CK(clk), .RN(n4860), .Q(n4359)
         );
  DFFR_X1 ex_mem_busA_q_reg_20_ ( .D(n3754), .CK(clk), .RN(n4860), .Q(n4579)
         );
  DFFR_X1 ex_mem_busA_q_reg_15_ ( .D(n3753), .CK(clk), .RN(n4860), .Q(n4578)
         );
  DFFR_X1 ex_mem_busA_q_reg_10_ ( .D(n3752), .CK(clk), .RN(n4856), .Q(n4492)
         );
  DFFR_X1 ex_mem_busA_q_reg_0_ ( .D(n3751), .CK(clk), .RN(n4859), .Q(n4673), 
        .QN(n8816) );
  DFFR_X1 ex_mem_rd_q_reg_4_ ( .D(n3750), .CK(clk), .RN(n4850), .Q(rd_3[4]), 
        .QN(n4320) );
  DFFR_X1 ex_mem_rd_q_reg_3_ ( .D(n3748), .CK(clk), .RN(n4866), .Q(rd_3[3]), 
        .QN(n4092) );
  DFFR_X1 ex_mem_op0_q_reg ( .D(n9177), .CK(clk), .RN(n4865), .Q(op0_3), .QN(
        n4651) );
  DFFR_X1 ex_mem_link_q_reg ( .D(n3745), .CK(clk), .RN(n4865), .Q(n4631), .QN(
        n8815) );
  DFFR_X1 ex_mem_jr_q_reg ( .D(n3743), .CK(clk), .RN(n4865), .Q(n4090), .QN(
        n8903) );
  DFFR_X1 ex_mem_branch_q_reg ( .D(n3742), .CK(clk), .RN(n4857), .QN(n8986) );
  DFFR_X1 ex_mem_jump_q_reg ( .D(n3741), .CK(clk), .RN(n4850), .QN(n8985) );
  DFFR_X1 ex_mem_memRd_q_reg ( .D(n3740), .CK(clk), .RN(n4850), .Q(n4362), 
        .QN(n8814) );
  DFFR_X1 ex_mem_imm32_q_reg_31_ ( .D(n3738), .CK(clk), .RN(n4853), .QN(n8850)
         );
  DFFR_X1 ex_mem_imm32_q_reg_30_ ( .D(n3737), .CK(clk), .RN(n4862), .QN(n8853)
         );
  DFFR_X1 ex_mem_imm32_q_reg_29_ ( .D(n3736), .CK(clk), .RN(n4862), .QN(n8855)
         );
  DFFR_X1 ex_mem_imm32_q_reg_28_ ( .D(n9173), .CK(clk), .RN(n4853), .Q(n4540), 
        .QN(n8967) );
  DFFR_X1 ex_mem_imm32_q_reg_27_ ( .D(n3734), .CK(clk), .RN(n4862), .QN(n8858)
         );
  DFFR_X1 ex_mem_imm32_q_reg_26_ ( .D(n9172), .CK(clk), .RN(n4853), .Q(n4541), 
        .QN(n8969) );
  DFFR_X1 ex_mem_imm32_q_reg_25_ ( .D(n3732), .CK(clk), .RN(n4862), .QN(n8861)
         );
  DFFR_X1 ex_mem_imm32_q_reg_24_ ( .D(n3731), .CK(clk), .RN(n4853), .Q(n4542), 
        .QN(n8862) );
  DFFR_X1 ex_mem_imm32_q_reg_23_ ( .D(n3730), .CK(clk), .RN(n4862), .QN(n8865)
         );
  DFFR_X1 ex_mem_imm32_q_reg_22_ ( .D(n3729), .CK(clk), .RN(n4853), .Q(n4464), 
        .QN(n8866) );
  DFFR_X1 ex_mem_imm32_q_reg_21_ ( .D(n3728), .CK(clk), .RN(n4862), .QN(n8869)
         );
  DFFR_X1 ex_mem_imm32_q_reg_20_ ( .D(n9171), .CK(clk), .RN(n4853), .Q(n4462), 
        .QN(n8971) );
  DFFR_X1 ex_mem_imm32_q_reg_19_ ( .D(n3726), .CK(clk), .RN(n4853), .QN(n8873)
         );
  DFFR_X1 ex_mem_imm32_q_reg_18_ ( .D(n9170), .CK(clk), .RN(n4871), .Q(n4463), 
        .QN(n8973) );
  DFFR_X1 ex_mem_imm32_q_reg_17_ ( .D(n3724), .CK(clk), .RN(n4853), .QN(n8876)
         );
  DFFR_X1 ex_mem_imm32_q_reg_16_ ( .D(n9169), .CK(clk), .RN(n4875), .QN(n8975)
         );
  DFFR_X1 ex_mem_imm32_q_reg_15_ ( .D(n3722), .CK(clk), .RN(n4854), .Q(n4465), 
        .QN(n8879) );
  DFFR_X1 ex_mem_imm32_q_reg_14_ ( .D(n3721), .CK(clk), .RN(n4864), .QN(n8880)
         );
  DFFR_X1 ex_mem_imm32_q_reg_13_ ( .D(n3720), .CK(clk), .RN(n4854), .Q(n4466), 
        .QN(n8883) );
  DFFR_X1 ex_mem_imm32_q_reg_12_ ( .D(n3719), .CK(clk), .RN(n4874), .QN(n8884)
         );
  DFFR_X1 ex_mem_imm32_q_reg_11_ ( .D(n3718), .CK(clk), .RN(n4854), .Q(n4403), 
        .QN(n8887) );
  DFFR_X1 ex_mem_imm32_q_reg_10_ ( .D(n3717), .CK(clk), .RN(n4863), .QN(n8888)
         );
  DFFR_X1 ex_mem_imm32_q_reg_9_ ( .D(n3716), .CK(clk), .RN(n4862), .Q(n4404), 
        .QN(n8891) );
  DFFR_X1 ex_mem_imm32_q_reg_8_ ( .D(n9176), .CK(clk), .RN(n4853), .QN(n8961)
         );
  DFFR_X1 ex_mem_imm32_q_reg_7_ ( .D(n3714), .CK(clk), .RN(n4862), .Q(n4405), 
        .QN(n8894) );
  DFFR_X1 ex_mem_imm32_q_reg_6_ ( .D(n9175), .CK(clk), .RN(n4853), .QN(n8963)
         );
  DFFR_X1 ex_mem_imm32_q_reg_5_ ( .D(n3712), .CK(clk), .RN(n4862), .Q(n4406), 
        .QN(n8897) );
  DFFR_X1 ex_mem_imm32_q_reg_4_ ( .D(n9174), .CK(clk), .RN(n4853), .QN(n8965)
         );
  DFFR_X1 ex_mem_imm32_q_reg_3_ ( .D(n3710), .CK(clk), .RN(n4862), .Q(n4402), 
        .QN(n8813) );
  DFFR_X1 ex_mem_imm32_q_reg_2_ ( .D(n3709), .CK(clk), .RN(n4853), .Q(n4408), 
        .QN(n8899) );
  DFFR_X1 ex_mem_imm32_q_reg_1_ ( .D(n3708), .CK(clk), .RN(n4872), .QN(n8812)
         );
  DFFR_X1 ex_mem_imm32_q_reg_0_ ( .D(n3707), .CK(clk), .RN(n4854), .Q(n4137), 
        .QN(n8901) );
  DFFR_X1 ex_mem_busB_q_reg_31_ ( .D(n3706), .CK(clk), .RN(n4866), .QN(n8811)
         );
  DFFR_X1 ex_mem_busB_q_reg_30_ ( .D(n3705), .CK(clk), .RN(n4854), .QN(n8810)
         );
  DFFR_X1 ex_mem_busB_q_reg_28_ ( .D(n3704), .CK(clk), .RN(n4861), .QN(n8809)
         );
  DFFR_X1 ex_mem_busB_q_reg_26_ ( .D(n3703), .CK(clk), .RN(n4861), .QN(n8808)
         );
  DFFR_X1 ex_mem_busB_q_reg_24_ ( .D(n3702), .CK(clk), .RN(n4861), .Q(n4682), 
        .QN(n8807) );
  DFFR_X1 ex_mem_busB_q_reg_23_ ( .D(n3701), .CK(clk), .RN(n4855), .QN(n8806)
         );
  DFFR_X1 ex_mem_busB_q_reg_16_ ( .D(n3700), .CK(clk), .RN(n4855), .Q(n4681), 
        .QN(n8805) );
  DFFR_X1 ex_mem_busB_q_reg_13_ ( .D(n3699), .CK(clk), .RN(n4861), .Q(n4701), 
        .QN(n8804) );
  DFFR_X1 ex_mem_busB_q_reg_11_ ( .D(n3698), .CK(clk), .RN(n4861), .Q(n4700), 
        .QN(n8803) );
  DFFR_X1 ex_mem_busB_q_reg_7_ ( .D(n3697), .CK(clk), .RN(n4854), .Q(n4699), 
        .QN(n8802) );
  DFFR_X1 ex_mem_busB_q_reg_1_ ( .D(n3696), .CK(clk), .RN(n4855), .Q(n4680), 
        .QN(n8801) );
  DFFR_X1 id_ex_instr_q_reg_1_ ( .D(n3693), .CK(clk), .RN(n4872), .QN(n8800)
         );
  DFFR_X1 ex_mem_instr_q_reg_1_ ( .D(n3692), .CK(clk), .RN(n4864), .Q(
        memInstr[1]), .QN(n8799) );
  DFFR_X1 id_ex_instr_q_reg_3_ ( .D(n3689), .CK(clk), .RN(n4873), .QN(n8915)
         );
  DFFR_X1 ex_mem_instr_q_reg_3_ ( .D(n3688), .CK(clk), .RN(n4865), .Q(
        memInstr[3]), .QN(n8798) );
  DFFR_X1 id_ex_instr_q_reg_5_ ( .D(n3685), .CK(clk), .RN(n4873), .QN(n8926)
         );
  DFFR_X1 ex_mem_instr_q_reg_5_ ( .D(n3684), .CK(clk), .RN(n4865), .Q(
        memInstr[5]), .QN(n8797) );
  DFFR_X1 id_ex_instr_q_reg_26_ ( .D(n3683), .CK(clk), .RN(n4843), .QN(n8929)
         );
  DFFR_X1 ex_mem_instr_q_reg_26_ ( .D(n3682), .CK(clk), .RN(n4850), .Q(
        memInstr[26]), .QN(n8796) );
  DFFR_X1 id_ex_instr_q_reg_27_ ( .D(n3681), .CK(clk), .RN(n4872), .QN(n8930)
         );
  DFFR_X1 ex_mem_instr_q_reg_27_ ( .D(n3680), .CK(clk), .RN(n4864), .Q(
        memInstr[27]), .QN(n8795) );
  DFFR_X1 id_ex_instr_q_reg_28_ ( .D(n3679), .CK(clk), .RN(n4843), .QN(n8928)
         );
  DFFR_X1 ex_mem_instr_q_reg_28_ ( .D(n3678), .CK(clk), .RN(n4850), .Q(
        memInstr[28]), .QN(n8794) );
  DFFR_X1 id_ex_instr_q_reg_29_ ( .D(n3677), .CK(clk), .RN(n4872), .QN(n8918)
         );
  DFFR_X1 ex_mem_instr_q_reg_29_ ( .D(n3676), .CK(clk), .RN(n4865), .Q(
        memInstr[29]), .QN(n8793) );
  DFFR_X1 id_ex_instr_q_reg_30_ ( .D(n3675), .CK(clk), .RN(n4873), .QN(n8917)
         );
  DFFR_X1 ex_mem_instr_q_reg_30_ ( .D(n3674), .CK(clk), .RN(n4865), .Q(
        memInstr[30]), .QN(n8792) );
  DFFR_X1 id_ex_memWr_q_reg ( .D(n3673), .CK(clk), .RN(n4842), .QN(n8791) );
  DFFR_X1 ex_mem_memWr_q_reg ( .D(n3672), .CK(clk), .RN(n4865), .Q(memWr), 
        .QN(n8790) );
  DFFR_X1 id_ex_regWr_q_reg ( .D(n3671), .CK(clk), .RN(n4843), .QN(n4610) );
  DFFR_X1 ex_mem_regWr_q_reg ( .D(n3670), .CK(clk), .RN(n4866), .QN(n4360) );
  DFFR_X1 if_id_incPC_q_reg_0_ ( .D(n3665), .CK(clk), .RN(n4865), .QN(n8789)
         );
  DFFR_X1 id_ex_incPC_q_reg_0_ ( .D(n3664), .CK(clk), .RN(n4845), .QN(n8788)
         );
  DFFR_X1 ex_mem_incPC_q_reg_0_ ( .D(n3663), .CK(clk), .RN(n4852), .Q(
        reg31Val_3[0]), .QN(n4532) );
  DFFR_X1 id_ex_zeroExt_q_reg ( .D(n3661), .CK(clk), .RN(n4874), .Q(zeroExt_2), 
        .QN(n4087) );
  DFFR_X1 id_ex_instr_q_reg_25_ ( .D(n3660), .CK(clk), .RN(n4872), .QN(n8931)
         );
  DFFR_X1 ex_mem_instr_q_reg_25_ ( .D(n3659), .CK(clk), .RN(n4864), .Q(
        memInstr[25]), .QN(n8787) );
  DFFR_X1 id_ex_instr_q_reg_24_ ( .D(n3658), .CK(clk), .RN(n4843), .Q(n4330), 
        .QN(n8786) );
  DFFR_X1 ex_mem_instr_q_reg_24_ ( .D(n3657), .CK(clk), .RN(n4851), .Q(
        memInstr[24]), .QN(n8785) );
  DFFR_X1 id_ex_instr_q_reg_23_ ( .D(n3656), .CK(clk), .RN(n4872), .QN(n8919)
         );
  DFFR_X1 ex_mem_instr_q_reg_23_ ( .D(n3655), .CK(clk), .RN(n4864), .Q(
        memInstr[23]), .QN(n8784) );
  DFFR_X1 id_ex_instr_q_reg_22_ ( .D(n3654), .CK(clk), .RN(n4843), .QN(n8920)
         );
  DFFR_X1 ex_mem_instr_q_reg_22_ ( .D(n3653), .CK(clk), .RN(n4851), .Q(
        memInstr[22]), .QN(n8783) );
  DFFR_X1 id_ex_instr_q_reg_21_ ( .D(n3652), .CK(clk), .RN(n4872), .QN(n8921)
         );
  DFFR_X1 ex_mem_instr_q_reg_21_ ( .D(n3651), .CK(clk), .RN(n4864), .Q(
        memInstr[21]), .QN(n8782) );
  DFFR_X1 id_ex_instr_q_reg_20_ ( .D(n3650), .CK(clk), .RN(n4843), .QN(n8922)
         );
  DFFR_X1 ex_mem_instr_q_reg_20_ ( .D(n3649), .CK(clk), .RN(n4851), .Q(
        memInstr[20]), .QN(n8781) );
  DFFR_X1 id_ex_instr_q_reg_19_ ( .D(n3648), .CK(clk), .RN(n4843), .QN(n8924)
         );
  DFFR_X1 ex_mem_instr_q_reg_19_ ( .D(n3647), .CK(clk), .RN(n4851), .Q(
        memInstr[19]), .QN(n8780) );
  DFFR_X1 id_ex_instr_q_reg_18_ ( .D(n3646), .CK(clk), .RN(n4872), .QN(n8923)
         );
  DFFR_X1 ex_mem_instr_q_reg_18_ ( .D(n3645), .CK(clk), .RN(n4864), .Q(
        memInstr[18]), .QN(n8779) );
  DFFR_X1 id_ex_instr_q_reg_17_ ( .D(n3644), .CK(clk), .RN(n4843), .QN(n8925)
         );
  DFFR_X1 ex_mem_instr_q_reg_17_ ( .D(n3643), .CK(clk), .RN(n4851), .Q(
        memInstr[17]), .QN(n8778) );
  DFFR_X1 id_ex_instr_q_reg_16_ ( .D(n3642), .CK(clk), .RN(n4872), .QN(n8909)
         );
  DFFR_X1 ex_mem_instr_q_reg_16_ ( .D(n3641), .CK(clk), .RN(n4864), .Q(
        memInstr[16]), .QN(n8777) );
  DFFR_X1 id_ex_instr_q_reg_15_ ( .D(n3640), .CK(clk), .RN(n4843), .QN(n8911)
         );
  DFFR_X1 ex_mem_instr_q_reg_15_ ( .D(n3639), .CK(clk), .RN(n4851), .Q(
        memInstr[15]), .QN(n8776) );
  DFFR_X1 id_ex_instr_q_reg_14_ ( .D(n3638), .CK(clk), .RN(n4872), .QN(n8912)
         );
  DFFR_X1 ex_mem_instr_q_reg_14_ ( .D(n3637), .CK(clk), .RN(n4864), .Q(
        memInstr[14]), .QN(n8775) );
  DFFR_X1 id_ex_instr_q_reg_13_ ( .D(n3636), .CK(clk), .RN(n4843), .QN(n8913)
         );
  DFFR_X1 ex_mem_instr_q_reg_13_ ( .D(n3635), .CK(clk), .RN(n4851), .Q(
        memInstr[13]), .QN(n8774) );
  DFFR_X1 id_ex_instr_q_reg_12_ ( .D(n3634), .CK(clk), .RN(n4872), .QN(n8914)
         );
  DFFR_X1 ex_mem_instr_q_reg_12_ ( .D(n3633), .CK(clk), .RN(n4864), .Q(
        memInstr[12]), .QN(n8773) );
  DFFR_X1 id_ex_instr_q_reg_11_ ( .D(n3632), .CK(clk), .RN(n4844), .QN(n8772)
         );
  DFFR_X1 ex_mem_instr_q_reg_11_ ( .D(n3631), .CK(clk), .RN(n4851), .Q(
        memInstr[11]), .QN(n8771) );
  DFFR_X1 id_ex_instr_q_reg_10_ ( .D(n3630), .CK(clk), .RN(n4872), .QN(n8770)
         );
  DFFR_X1 ex_mem_instr_q_reg_10_ ( .D(n3629), .CK(clk), .RN(n4864), .Q(
        memInstr[10]), .QN(n8769) );
  DFFR_X1 id_ex_instr_q_reg_9_ ( .D(n3628), .CK(clk), .RN(n4873), .Q(n4544), 
        .QN(n8768) );
  DFFR_X1 ex_mem_instr_q_reg_9_ ( .D(n3627), .CK(clk), .RN(n4865), .Q(
        memInstr[9]), .QN(n8767) );
  DFFR_X1 id_ex_instr_q_reg_8_ ( .D(n3626), .CK(clk), .RN(n4843), .Q(n4131), 
        .QN(n8766) );
  DFFR_X1 ex_mem_instr_q_reg_8_ ( .D(n3625), .CK(clk), .RN(n4850), .Q(
        memInstr[8]), .QN(n8765) );
  DFFR_X1 id_ex_instr_q_reg_7_ ( .D(n3624), .CK(clk), .RN(n4873), .QN(n8910)
         );
  DFFR_X1 ex_mem_instr_q_reg_7_ ( .D(n3623), .CK(clk), .RN(n4865), .Q(
        memInstr[7]), .QN(n8764) );
  DFFR_X1 id_ex_instr_q_reg_6_ ( .D(n3622), .CK(clk), .RN(n4843), .QN(n8927)
         );
  DFFR_X1 ex_mem_instr_q_reg_6_ ( .D(n3621), .CK(clk), .RN(n4850), .Q(
        memInstr[6]), .QN(n8763) );
  DFFR_X1 id_ex_valid_q_reg ( .D(n3620), .CK(clk), .RN(n4844), .Q(valid_2), 
        .QN(n4361) );
  DFFR_X1 ex_mem_valid_q_reg ( .D(n3619), .CK(clk), .RN(n4849), .Q(valid_3), 
        .QN(n4612) );
  DFFR_X1 id_ex_busB_sel_q_reg_1_ ( .D(n3618), .CK(clk), .RN(n4846), .Q(n4140), 
        .QN(n9057) );
  DFFR_X1 id_ex_busA_sel_q_reg_1_ ( .D(n3617), .CK(clk), .RN(n4848), .Q(n4373), 
        .QN(n9052) );
  DFFR_X1 id_ex_busB_sel_q_reg_0_ ( .D(n3616), .CK(clk), .RN(n4869), .Q(n4139), 
        .QN(n9058) );
  DFFR_X1 ex_mem_busB_q_reg_0_ ( .D(n3615), .CK(clk), .RN(n4861), .Q(n4679), 
        .QN(n8762) );
  DFFR_X1 id_ex_busA_sel_q_reg_0_ ( .D(n3614), .CK(clk), .RN(n4867), .Q(n4156), 
        .QN(n9053) );
  DFFR_X1 ex_mem_busA_q_reg_1_ ( .D(n3613), .CK(clk), .RN(n4856), .Q(n4672), 
        .QN(n8761) );
  DFFR_X1 if_id_incPC_q_reg_1_ ( .D(n3611), .CK(clk), .RN(n4874), .QN(n8760)
         );
  DFFR_X1 id_ex_incPC_q_reg_1_ ( .D(n3610), .CK(clk), .RN(n4871), .QN(n8759)
         );
  DFFR_X1 ex_mem_incPC_q_reg_1_ ( .D(n3609), .CK(clk), .RN(n4863), .Q(
        reg31Val_3[1]), .QN(n4368) );
  DFFR_X1 ex_mem_busA_q_reg_21_ ( .D(n3607), .CK(clk), .RN(n4856), .Q(n4358)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_22_ ( .D(n9161), .CK(clk), .RN(n4857), .Q(
        memAddr[22]), .QN(n9028) );
  DFFR_X1 ex_mem_busA_q_reg_22_ ( .D(n3604), .CK(clk), .RN(n4860), .Q(n4357)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_9_ ( .D(n3603), .CK(clk), .RN(n4859), .Q(
        memAddr[9]), .QN(n9004) );
  DFFR_X1 ex_mem_busB_q_reg_9_ ( .D(n3601), .CK(clk), .RN(n4854), .Q(n4678), 
        .QN(n8758) );
  DFFR_X1 ex_mem_aluRes_q_reg_17_ ( .D(n3600), .CK(clk), .RN(n4858), .Q(
        memAddr[17]), .QN(n9018) );
  DFFR_X1 ex_mem_busA_q_reg_17_ ( .D(n3598), .CK(clk), .RN(n4860), .Q(n4577)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_12_ ( .D(n3597), .CK(clk), .RN(n4858), .Q(
        memAddr[12]), .QN(n9008) );
  DFFR_X1 ex_mem_busA_q_reg_12_ ( .D(n3595), .CK(clk), .RN(n4856), .Q(n4491)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_29_ ( .D(n9167), .CK(clk), .RN(n4859), .Q(
        memAddr[29]), .QN(n9045) );
  DFFR_X1 ex_mem_busA_q_reg_29_ ( .D(n3592), .CK(clk), .RN(n4856), .Q(n4356)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_8_ ( .D(n3591), .CK(clk), .RN(n4857), .Q(
        memAddr[8]), .QN(n9002) );
  DFFR_X1 ex_mem_busA_q_reg_8_ ( .D(n3589), .CK(clk), .RN(n4861), .Q(n4490) );
  DFFR_X1 ex_mem_aluRes_q_reg_25_ ( .D(n9164), .CK(clk), .RN(n4859), .Q(
        memAddr[25]), .QN(n9037) );
  DFFR_X1 ex_mem_busA_q_reg_25_ ( .D(n3586), .CK(clk), .RN(n4856), .Q(n4355)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_18_ ( .D(n9157), .CK(clk), .RN(n4858), .Q(
        memAddr[18]), .QN(n9020) );
  DFFR_X1 ex_mem_busA_q_reg_18_ ( .D(n3583), .CK(clk), .RN(n4856), .Q(n4576)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_27_ ( .D(n9166), .CK(clk), .RN(n4859), .Q(
        memAddr[27]), .QN(n9041) );
  DFFR_X1 ex_mem_busA_q_reg_27_ ( .D(n3580), .CK(clk), .RN(n4856), .Q(n4354)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_4_ ( .D(n3579), .CK(clk), .RN(n4857), .Q(
        memAddr[4]), .QN(n8995) );
  DFFR_X1 ex_mem_busB_q_reg_4_ ( .D(n3577), .CK(clk), .RN(n4867), .Q(n4698), 
        .QN(n8757) );
  DFFR_X1 ex_mem_aluRes_q_reg_19_ ( .D(n9158), .CK(clk), .RN(n4857), .Q(
        memAddr[19]), .QN(n9022) );
  DFFR_X1 ex_mem_busA_q_reg_19_ ( .D(n3574), .CK(clk), .RN(n4860), .Q(n4575)
         );
  DFFR_X1 if_id_incPC_q_reg_19_ ( .D(n3572), .CK(clk), .RN(n4842), .QN(n8755)
         );
  DFFR_X1 id_ex_incPC_q_reg_19_ ( .D(n3571), .CK(clk), .RN(n4844), .QN(n8754)
         );
  DFFR_X1 ex_mem_incPC_q_reg_19_ ( .D(n3570), .CK(clk), .RN(n4852), .Q(n4458), 
        .QN(n8872) );
  DFFR_X1 if_id_incPC_q_reg_20_ ( .D(n3568), .CK(clk), .RN(n4842), .QN(n8752)
         );
  DFFR_X1 id_ex_incPC_q_reg_20_ ( .D(n3567), .CK(clk), .RN(n4844), .QN(n8751)
         );
  DFFR_X1 ex_mem_incPC_q_reg_20_ ( .D(n3566), .CK(clk), .RN(n4852), .Q(n4279), 
        .QN(n8870) );
  DFFR_X1 if_id_incPC_q_reg_21_ ( .D(n3564), .CK(clk), .RN(n4874), .QN(n8749)
         );
  DFFR_X1 id_ex_incPC_q_reg_21_ ( .D(n3563), .CK(clk), .RN(n4871), .QN(n8748)
         );
  DFFR_X1 ex_mem_incPC_q_reg_21_ ( .D(n3562), .CK(clk), .RN(n4863), .Q(n4457), 
        .QN(n8868) );
  DFFR_X1 if_id_incPC_q_reg_23_ ( .D(n3560), .CK(clk), .RN(n4874), .QN(n8746)
         );
  DFFR_X1 id_ex_incPC_q_reg_23_ ( .D(n3559), .CK(clk), .RN(n4871), .QN(n8745)
         );
  DFFR_X1 ex_mem_incPC_q_reg_23_ ( .D(n3558), .CK(clk), .RN(n4863), .Q(n4456), 
        .QN(n8864) );
  DFFR_X1 if_id_incPC_q_reg_24_ ( .D(n3556), .CK(clk), .RN(n4842), .QN(n8743)
         );
  DFFR_X1 id_ex_incPC_q_reg_24_ ( .D(n3555), .CK(clk), .RN(n4844), .QN(n8742)
         );
  DFFR_X1 ex_mem_incPC_q_reg_24_ ( .D(n3554), .CK(clk), .RN(n4852), .Q(n4325), 
        .QN(n8863) );
  DFFR_X1 if_id_incPC_q_reg_25_ ( .D(n3552), .CK(clk), .RN(n4874), .QN(n8740)
         );
  DFFR_X1 id_ex_incPC_q_reg_25_ ( .D(n3551), .CK(clk), .RN(n4871), .QN(n8739)
         );
  DFFR_X1 ex_mem_incPC_q_reg_25_ ( .D(n3550), .CK(clk), .RN(n4863), .Q(n4536), 
        .QN(n8860) );
  DFFR_X1 if_id_incPC_q_reg_26_ ( .D(n3548), .CK(clk), .RN(n4842), .QN(n8737)
         );
  DFFR_X1 id_ex_incPC_q_reg_26_ ( .D(n3547), .CK(clk), .RN(n4844), .QN(n8736)
         );
  DFFR_X1 ex_mem_incPC_q_reg_26_ ( .D(n3546), .CK(clk), .RN(n4852), .Q(n4327), 
        .QN(n8859) );
  DFFR_X1 if_id_incPC_q_reg_27_ ( .D(n3544), .CK(clk), .RN(n4874), .QN(n8734)
         );
  DFFR_X1 id_ex_incPC_q_reg_27_ ( .D(n3543), .CK(clk), .RN(n4871), .QN(n8733)
         );
  DFFR_X1 ex_mem_incPC_q_reg_27_ ( .D(n3542), .CK(clk), .RN(n4863), .Q(n4535), 
        .QN(n8857) );
  DFFR_X1 if_id_incPC_q_reg_28_ ( .D(n3540), .CK(clk), .RN(n4842), .QN(n8731)
         );
  DFFR_X1 id_ex_incPC_q_reg_28_ ( .D(n3539), .CK(clk), .RN(n4844), .QN(n8730)
         );
  DFFR_X1 ex_mem_incPC_q_reg_28_ ( .D(n3538), .CK(clk), .RN(n4852), .Q(n4326), 
        .QN(n8856) );
  DFFR_X1 if_id_incPC_q_reg_29_ ( .D(n3536), .CK(clk), .RN(n4874), .QN(n8728)
         );
  DFFR_X1 id_ex_incPC_q_reg_29_ ( .D(n3535), .CK(clk), .RN(n4871), .QN(n8727)
         );
  DFFR_X1 ex_mem_incPC_q_reg_29_ ( .D(n3534), .CK(clk), .RN(n4863), .Q(n4534), 
        .QN(n8854) );
  DFFR_X1 if_id_incPC_q_reg_30_ ( .D(n3532), .CK(clk), .RN(n4875), .QN(n8725)
         );
  DFFR_X1 id_ex_incPC_q_reg_30_ ( .D(n3531), .CK(clk), .RN(n4871), .QN(n8724)
         );
  DFFR_X1 ex_mem_incPC_q_reg_30_ ( .D(n3530), .CK(clk), .RN(n4863), .Q(n4526), 
        .QN(n8852) );
  DFFR_X1 ex_mem_busA_q_reg_30_ ( .D(n3528), .CK(clk), .RN(n4856), .Q(n4353)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_2_ ( .D(n3527), .CK(clk), .RN(n4857), .Q(
        memAddr[2]), .QN(n8991) );
  DFFR_X1 ex_mem_busA_q_reg_2_ ( .D(n3525), .CK(clk), .RN(n4860), .Q(n4489) );
  DFFR_X1 if_id_incPC_q_reg_2_ ( .D(n3523), .CK(clk), .RN(n4842), .QN(n8723)
         );
  DFFR_X1 id_ex_incPC_q_reg_2_ ( .D(n3522), .CK(clk), .RN(n4844), .QN(n8722)
         );
  DFFR_X1 ex_mem_incPC_q_reg_2_ ( .D(n3521), .CK(clk), .RN(n4852), .Q(n4109), 
        .QN(n8900) );
  DFFR_X1 ex_mem_busB_q_reg_2_ ( .D(n3519), .CK(clk), .RN(n4873), .Q(n4697), 
        .QN(n8721) );
  DFFR_X1 ex_mem_aluRes_q_reg_5_ ( .D(n3518), .CK(clk), .RN(n4859), .Q(
        memAddr[5]), .QN(n8996) );
  DFFR_X1 ex_mem_busB_q_reg_5_ ( .D(n3516), .CK(clk), .RN(n4854), .Q(n4696), 
        .QN(n8720) );
  DFFR_X1 ex_mem_aluRes_q_reg_6_ ( .D(n3515), .CK(clk), .RN(n4857), .Q(
        memAddr[6]), .QN(n8998) );
  DFFR_X1 ex_mem_busA_q_reg_6_ ( .D(n3513), .CK(clk), .RN(n4860), .Q(n4488) );
  DFFR_X1 ex_mem_aluRes_q_reg_14_ ( .D(n3512), .CK(clk), .RN(n4858), .Q(
        memAddr[14]), .QN(n9011) );
  DFFR_X1 ex_mem_busA_q_reg_14_ ( .D(n3510), .CK(clk), .RN(n4856), .Q(n4487)
         );
  DFFR_X1 if_id_incPC_q_reg_15_ ( .D(n3508), .CK(clk), .RN(n4842), .QN(n8718)
         );
  DFFR_X1 id_ex_incPC_q_reg_15_ ( .D(n3507), .CK(clk), .RN(n4845), .QN(n8717)
         );
  DFFR_X1 ex_mem_incPC_q_reg_15_ ( .D(n3506), .CK(clk), .RN(n4852), .Q(n4276), 
        .QN(n8878) );
  DFFR_X1 if_id_incPC_q_reg_16_ ( .D(n3504), .CK(clk), .RN(n4874), .QN(n8715)
         );
  DFFR_X1 id_ex_incPC_q_reg_16_ ( .D(n3503), .CK(clk), .RN(n4871), .QN(n8714)
         );
  DFFR_X1 ex_mem_incPC_q_reg_16_ ( .D(n3502), .CK(clk), .RN(n4863), .Q(n4453), 
        .QN(n8877) );
  DFFR_X1 if_id_incPC_q_reg_17_ ( .D(n3500), .CK(clk), .RN(n4842), .QN(n8712)
         );
  DFFR_X1 id_ex_incPC_q_reg_17_ ( .D(n3499), .CK(clk), .RN(n4845), .QN(n8711)
         );
  DFFR_X1 ex_mem_incPC_q_reg_17_ ( .D(n3498), .CK(clk), .RN(n4852), .Q(n4459), 
        .QN(n8875) );
  DFFR_X1 if_id_incPC_q_reg_18_ ( .D(n3496), .CK(clk), .RN(n4874), .QN(n8709)
         );
  DFFR_X1 id_ex_incPC_q_reg_18_ ( .D(n3495), .CK(clk), .RN(n4871), .QN(n8708)
         );
  DFFR_X1 ex_mem_incPC_q_reg_18_ ( .D(n3494), .CK(clk), .RN(n4863), .Q(n4280), 
        .QN(n8874) );
  DFFR_X1 if_id_incPC_q_reg_22_ ( .D(n3492), .CK(clk), .RN(n4842), .QN(n8706)
         );
  DFFR_X1 id_ex_incPC_q_reg_22_ ( .D(n3491), .CK(clk), .RN(n4844), .QN(n8705)
         );
  DFFR_X1 ex_mem_incPC_q_reg_22_ ( .D(n3490), .CK(clk), .RN(n4852), .Q(n4278), 
        .QN(n8867) );
  DFFR_X1 ex_mem_busA_q_reg_28_ ( .D(n3487), .CK(clk), .RN(n4860), .Q(n4352)
         );
  DFFR_X1 ex_mem_aluRes_q_reg_3_ ( .D(n3486), .CK(clk), .RN(n4859), .Q(
        memAddr[3]), .QN(n8993) );
  DFFR_X1 ex_mem_busA_q_reg_3_ ( .D(n3484), .CK(clk), .RN(n4855), .Q(n4486) );
  DFFR_X1 if_id_incPC_q_reg_3_ ( .D(n3482), .CK(clk), .RN(n4875), .QN(n8703)
         );
  DFFR_X1 id_ex_incPC_q_reg_3_ ( .D(n3481), .CK(clk), .RN(n4871), .QN(n8702)
         );
  DFFR_X1 ex_mem_incPC_q_reg_3_ ( .D(n3480), .CK(clk), .RN(n4863), .Q(n4174), 
        .QN(n8847) );
  DFFR_X1 if_id_incPC_q_reg_4_ ( .D(n3477), .CK(clk), .RN(n4842), .QN(n8700)
         );
  DFFR_X1 id_ex_incPC_q_reg_4_ ( .D(n3476), .CK(clk), .RN(n4844), .QN(n8699)
         );
  DFFR_X1 ex_mem_incPC_q_reg_4_ ( .D(n3475), .CK(clk), .RN(n4851), .Q(n4401), 
        .QN(n8898) );
  DFFR_X1 ex_mem_busA_q_reg_4_ ( .D(n3473), .CK(clk), .RN(n4860), .Q(n4485) );
  DFFR_X1 if_id_incPC_q_reg_5_ ( .D(n3471), .CK(clk), .RN(n4875), .QN(n8697)
         );
  DFFR_X1 id_ex_incPC_q_reg_5_ ( .D(n3470), .CK(clk), .RN(n4871), .QN(n8696)
         );
  DFFR_X1 ex_mem_incPC_q_reg_5_ ( .D(n3469), .CK(clk), .RN(n4863), .Q(n4173), 
        .QN(n8896) );
  DFFR_X1 ex_mem_busA_q_reg_5_ ( .D(n3467), .CK(clk), .RN(n4855), .Q(n4484) );
  DFFR_X1 if_id_incPC_q_reg_6_ ( .D(n3465), .CK(clk), .RN(n4842), .QN(n8694)
         );
  DFFR_X1 id_ex_incPC_q_reg_6_ ( .D(n3464), .CK(clk), .RN(n4844), .QN(n8693)
         );
  DFFR_X1 ex_mem_incPC_q_reg_6_ ( .D(n3463), .CK(clk), .RN(n4851), .Q(n4400), 
        .QN(n8895) );
  DFFR_X1 if_id_incPC_q_reg_7_ ( .D(n3460), .CK(clk), .RN(n4875), .QN(n8691)
         );
  DFFR_X1 id_ex_incPC_q_reg_7_ ( .D(n3459), .CK(clk), .RN(n4871), .QN(n8690)
         );
  DFFR_X1 ex_mem_incPC_q_reg_7_ ( .D(n3458), .CK(clk), .RN(n4864), .Q(n4172), 
        .QN(n8893) );
  DFFR_X1 ex_mem_busA_q_reg_7_ ( .D(n3456), .CK(clk), .RN(n4855), .Q(n4483) );
  DFFR_X1 if_id_incPC_q_reg_8_ ( .D(n3454), .CK(clk), .RN(n4841), .QN(n8688)
         );
  DFFR_X1 id_ex_incPC_q_reg_8_ ( .D(n3453), .CK(clk), .RN(n4844), .QN(n8687)
         );
  DFFR_X1 ex_mem_incPC_q_reg_8_ ( .D(n3452), .CK(clk), .RN(n4851), .Q(n4399), 
        .QN(n8892) );
  DFFR_X1 if_id_incPC_q_reg_9_ ( .D(n3449), .CK(clk), .RN(n4875), .QN(n8685)
         );
  DFFR_X1 id_ex_incPC_q_reg_9_ ( .D(n3448), .CK(clk), .RN(n4872), .QN(n8684)
         );
  DFFR_X1 ex_mem_incPC_q_reg_9_ ( .D(n3447), .CK(clk), .RN(n4864), .Q(n4171), 
        .QN(n8890) );
  DFFR_X1 ex_mem_busA_q_reg_9_ ( .D(n3445), .CK(clk), .RN(n4855), .Q(n4482) );
  DFFR_X1 if_id_incPC_q_reg_10_ ( .D(n3443), .CK(clk), .RN(n4874), .QN(n8682)
         );
  DFFR_X1 id_ex_incPC_q_reg_10_ ( .D(n3442), .CK(clk), .RN(n4870), .QN(n8681)
         );
  DFFR_X1 ex_mem_incPC_q_reg_10_ ( .D(n3441), .CK(clk), .RN(n4862), .Q(n4398), 
        .QN(n8889) );
  DFFR_X1 if_id_incPC_q_reg_11_ ( .D(n3438), .CK(clk), .RN(n4839), .QN(n8679)
         );
  DFFR_X1 id_ex_incPC_q_reg_11_ ( .D(n3437), .CK(clk), .RN(n4845), .QN(n8678)
         );
  DFFR_X1 ex_mem_incPC_q_reg_11_ ( .D(n3436), .CK(clk), .RN(n4852), .Q(n4170), 
        .QN(n8886) );
  DFFR_X1 ex_mem_busA_q_reg_11_ ( .D(n3434), .CK(clk), .RN(n4859), .Q(n4481)
         );
  DFFR_X1 if_id_incPC_q_reg_12_ ( .D(n3432), .CK(clk), .RN(n4874), .QN(n8676)
         );
  DFFR_X1 id_ex_incPC_q_reg_12_ ( .D(n3431), .CK(clk), .RN(n4870), .QN(n8675)
         );
  DFFR_X1 ex_mem_incPC_q_reg_12_ ( .D(n3430), .CK(clk), .RN(n4862), .Q(n4397), 
        .QN(n8885) );
  DFFR_X1 if_id_incPC_q_reg_13_ ( .D(n3427), .CK(clk), .RN(n4840), .QN(n8673)
         );
  DFFR_X1 id_ex_incPC_q_reg_13_ ( .D(n3426), .CK(clk), .RN(n4845), .QN(n8672)
         );
  DFFR_X1 ex_mem_incPC_q_reg_13_ ( .D(n3425), .CK(clk), .RN(n4852), .Q(n4277), 
        .QN(n8882) );
  DFFR_X1 ex_mem_busA_q_reg_13_ ( .D(n3423), .CK(clk), .RN(n4859), .Q(n4480)
         );
  DFFR_X1 if_id_incPC_q_reg_14_ ( .D(n3421), .CK(clk), .RN(n4874), .QN(n8670)
         );
  DFFR_X1 id_ex_incPC_q_reg_14_ ( .D(n3420), .CK(clk), .RN(n4870), .QN(n8669)
         );
  DFFR_X1 ex_mem_incPC_q_reg_14_ ( .D(n3419), .CK(clk), .RN(n4863), .Q(n4454), 
        .QN(n8881) );
  DFFR_X1 ex_mem_busA_q_reg_16_ ( .D(n3412), .CK(clk), .RN(n4856), .Q(n4574)
         );
  DFFR_X1 ex_mem_busB_q_reg_3_ ( .D(n3409), .CK(clk), .RN(n4854), .Q(n4695), 
        .QN(n8668) );
  DFFR_X1 ex_mem_busA_q_reg_26_ ( .D(n3406), .CK(clk), .RN(n4860), .Q(n4351)
         );
  DFFR_X1 ex_mem_busA_q_reg_24_ ( .D(n3403), .CK(clk), .RN(n4860), .Q(n4350)
         );
  DFFR_X1 ex_mem_busA_q_reg_23_ ( .D(n3401), .CK(clk), .RN(n4856), .Q(n4349)
         );
  DFFR_X1 ex_mem_busB_q_reg_14_ ( .D(n3399), .CK(clk), .RN(n4855), .Q(n4694), 
        .QN(n8667) );
  DFFR_X1 ex_mem_busB_q_reg_6_ ( .D(n3398), .CK(clk), .RN(n4870), .Q(n4693), 
        .QN(n8666) );
  DFFR_X1 if_id_incPC_q_reg_31_ ( .D(n3396), .CK(clk), .RN(n4842), .QN(n8664)
         );
  DFFR_X1 id_ex_incPC_q_reg_31_ ( .D(n3395), .CK(clk), .RN(n4844), .QN(n8663)
         );
  DFFR_X1 ex_mem_incPC_q_reg_31_ ( .D(n3394), .CK(clk), .RN(n4851), .QN(n8851)
         );
  DFFR_X1 ex_mem_busB_q_reg_19_ ( .D(n3392), .CK(clk), .RN(n4861), .Q(n4692), 
        .QN(n8662) );
  DFFR_X1 ex_mem_busB_q_reg_27_ ( .D(n3391), .CK(clk), .RN(n4854), .Q(n4691), 
        .QN(n8661) );
  DFFR_X1 ex_mem_busB_q_reg_18_ ( .D(n3390), .CK(clk), .RN(n4855), .Q(n4690), 
        .QN(n8660) );
  DFFR_X1 ex_mem_busB_q_reg_25_ ( .D(n3389), .CK(clk), .RN(n4854), .Q(n4677), 
        .QN(n8659) );
  DFFR_X1 ex_mem_busB_q_reg_8_ ( .D(n3388), .CK(clk), .RN(n4868), .Q(n4676), 
        .QN(n8658) );
  DFFR_X1 ex_mem_busB_q_reg_29_ ( .D(n3387), .CK(clk), .RN(n4854), .Q(n4689), 
        .QN(n8657) );
  DFFR_X1 ex_mem_busB_q_reg_12_ ( .D(n3386), .CK(clk), .RN(n4855), .Q(n4688), 
        .QN(n8656) );
  DFFR_X1 ex_mem_busB_q_reg_17_ ( .D(n3385), .CK(clk), .RN(n4861), .Q(n4675), 
        .QN(n8655) );
  DFFR_X1 ex_mem_busB_q_reg_22_ ( .D(n3384), .CK(clk), .RN(n4861), .Q(n4687), 
        .QN(n8654) );
  DFFR_X1 ex_mem_aluRes_q_reg_21_ ( .D(n9160), .CK(clk), .RN(n4858), .Q(
        memAddr[21]), .QN(n9026) );
  DFFR_X1 ex_mem_busB_q_reg_21_ ( .D(n3381), .CK(clk), .RN(n4855), .Q(n4686), 
        .QN(n8653) );
  DFFR_X1 id_ex_instr_q_reg_31_ ( .D(n3380), .CK(clk), .RN(n4843), .QN(n8916)
         );
  DFFR_X1 id_ex_memWrData_sel_q_reg_1_ ( .D(n3379), .CK(clk), .RN(n4873), .QN(
        n8652) );
  DFFR_X1 ex_mem_memWrData_sel_q_reg_1_ ( .D(n3378), .CK(clk), .RN(n4850), .Q(
        n4331), .QN(n8848) );
  DFFR_X1 id_ex_memWrData_sel_q_reg_0_ ( .D(n3377), .CK(clk), .RN(n4845), .QN(
        n8651) );
  DFFR_X1 ex_mem_memWrData_sel_q_reg_0_ ( .D(n3376), .CK(clk), .RN(n4865), .Q(
        n4549), .QN(n8849) );
  DFFR_X1 ex_mem_instr_q_reg_31_ ( .D(n3375), .CK(clk), .RN(n4850), .Q(
        memInstr[31]), .QN(n8650) );
  DFFR_X1 ex_mem_busB_q_reg_20_ ( .D(n3374), .CK(clk), .RN(n4861), .Q(n4685), 
        .QN(n8649) );
  DFFR_X1 ex_mem_busB_q_reg_10_ ( .D(n3373), .CK(clk), .RN(n4855), .Q(n4684), 
        .QN(n8648) );
  DFFR_X1 ex_mem_busB_q_reg_15_ ( .D(n3372), .CK(clk), .RN(n4861), .Q(n4683), 
        .QN(n8647) );
  DFFS_X2 hazard_detect_multiplier_fsm_pc_mult_ctrl_reg ( .D(
        hazard_detect_multiplier_fsm_N19), .CK(clk), .SN(n4878), .QN(n7613) );
  DFFS_X2 hazard_detect_multiplier_fsm_mem_wb_mult_ctrl_reg_1_ ( .D(
        hazard_detect_multiplier_fsm_N19), .CK(clk), .SN(n4877), .QN(n7853) );
  DFF_X2 mem_wb_memRdData_q_reg_31_ ( .D(n9066), .CK(clk), .Q(
        wb_dsize_reg_z2[31]), .QN(n4702) );
  DFFS_X2 if_id_instr_q_reg_0_ ( .D(n3897), .CK(clk), .SN(n4877), .Q(n4321), 
        .QN(n7612) );
  DFFS_X2 if_id_instr_q_reg_2_ ( .D(n3896), .CK(clk), .SN(n4877), .Q(n4539), 
        .QN(n7611) );
  DFFS_X2 if_id_instr_q_reg_4_ ( .D(n3895), .CK(clk), .SN(n4877), .Q(n4129), 
        .QN(n7610) );
  DFFS_X2 if_id_valid_q_reg ( .D(n3894), .CK(clk), .SN(n4877), .QN(n4611) );
  DFF_X2 mem_wb_aluRes_q_reg_0_ ( .D(n3813), .CK(clk), .QN(n7609) );
  DFF_X2 mem_wb_aluRes_q_reg_1_ ( .D(n3812), .CK(clk), .QN(n7608) );
  DFF_X2 mem_wb_aluRes_q_reg_7_ ( .D(n3811), .CK(clk), .QN(n7607) );
  DFF_X2 mem_wb_aluRes_q_reg_10_ ( .D(n3810), .CK(clk), .Q(n4621) );
  DFF_X2 mem_wb_aluRes_q_reg_11_ ( .D(n3809), .CK(clk), .Q(n4622) );
  DFF_X2 mem_wb_aluRes_q_reg_13_ ( .D(n3808), .CK(clk), .Q(n4447), .QN(n7606)
         );
  DFF_X2 mem_wb_aluRes_q_reg_15_ ( .D(n3807), .CK(clk), .QN(n7605) );
  DFF_X2 mem_wb_aluRes_q_reg_16_ ( .D(n3806), .CK(clk), .QN(n7604) );
  DFF_X2 mem_wb_aluRes_q_reg_20_ ( .D(n3805), .CK(clk), .QN(n7603) );
  DFF_X2 mem_wb_aluRes_q_reg_23_ ( .D(n3804), .CK(clk), .QN(n7602) );
  DFF_X2 mem_wb_aluRes_q_reg_24_ ( .D(n3803), .CK(clk), .Q(n4613), .QN(n7601)
         );
  DFF_X2 mem_wb_aluRes_q_reg_26_ ( .D(n3802), .CK(clk), .Q(n4450), .QN(n7600)
         );
  DFF_X2 mem_wb_aluRes_q_reg_28_ ( .D(n3801), .CK(clk), .Q(n4449), .QN(n7599)
         );
  DFF_X2 mem_wb_aluRes_q_reg_30_ ( .D(n3800), .CK(clk), .Q(n4623) );
  DFF_X2 mem_wb_aluRes_q_reg_31_ ( .D(n3799), .CK(clk), .Q(n4614), .QN(n7598)
         );
  DFF_X2 mem_wb_memRdData_q_reg_0_ ( .D(n9090), .CK(clk), .Q(
        wb_dsize_reg_z2[0]), .QN(n4632) );
  DFF_X2 mem_wb_memRdData_q_reg_1_ ( .D(n9079), .CK(clk), .Q(
        wb_dsize_reg_z2[1]), .QN(n4644) );
  DFF_X2 mem_wb_memRdData_q_reg_2_ ( .D(n9068), .CK(clk), .Q(
        wb_dsize_reg_z2[2]), .QN(n4643) );
  DFF_X2 mem_wb_memRdData_q_reg_3_ ( .D(n9065), .CK(clk), .Q(
        wb_dsize_reg_z2[3]), .QN(n4642) );
  DFF_X2 mem_wb_memRdData_q_reg_4_ ( .D(n9064), .CK(clk), .Q(
        wb_dsize_reg_z2[4]), .QN(n4641) );
  DFF_X2 mem_wb_memRdData_q_reg_5_ ( .D(n9063), .CK(clk), .Q(
        wb_dsize_reg_z2[5]), .QN(n4640) );
  DFF_X2 mem_wb_memRdData_q_reg_6_ ( .D(n9062), .CK(clk), .Q(
        wb_dsize_reg_z2[6]), .QN(n4639) );
  DFF_X2 mem_wb_memRdData_q_reg_7_ ( .D(n9061), .CK(clk), .Q(
        wb_dsize_reg_z2[7]), .QN(n4638) );
  DFF_X2 mem_wb_memRdData_q_reg_8_ ( .D(n9060), .CK(clk), .Q(
        wb_dsize_reg_z2[8]), .QN(n4636) );
  DFF_X2 mem_wb_memRdData_q_reg_9_ ( .D(n9059), .CK(clk), .Q(
        wb_dsize_reg_z2[9]), .QN(n4635) );
  DFF_X2 mem_wb_memRdData_q_reg_10_ ( .D(n9089), .CK(clk), .Q(
        wb_dsize_reg_z2[10]), .QN(n4649) );
  DFF_X2 mem_wb_memRdData_q_reg_11_ ( .D(n9088), .CK(clk), .Q(
        wb_dsize_reg_z2[11]), .QN(n4648) );
  DFF_X2 mem_wb_memRdData_q_reg_12_ ( .D(n9087), .CK(clk), .Q(
        wb_dsize_reg_z2[12]), .QN(n4647) );
  DFF_X2 mem_wb_memRdData_q_reg_13_ ( .D(n9086), .CK(clk), .Q(
        wb_dsize_reg_z2[13]), .QN(n4646) );
  DFF_X2 mem_wb_memRdData_q_reg_14_ ( .D(n9085), .CK(clk), .Q(
        wb_dsize_reg_z2[14]), .QN(n4645) );
  DFF_X2 mem_wb_memRdData_q_reg_15_ ( .D(n9084), .CK(clk), .Q(
        wb_dsize_reg_z2[15]), .QN(n4637) );
  DFF_X2 mem_wb_memRdData_q_reg_16_ ( .D(n9083), .CK(clk), .Q(
        wb_dsize_reg_z2[16]), .QN(n4724) );
  DFF_X2 mem_wb_memRdData_q_reg_17_ ( .D(n9082), .CK(clk), .Q(
        wb_dsize_reg_z2[17]), .QN(n4723) );
  DFF_X2 mem_wb_memRdData_q_reg_18_ ( .D(n9081), .CK(clk), .Q(
        wb_dsize_reg_z2[18]), .QN(n4722) );
  DFF_X2 mem_wb_memRdData_q_reg_19_ ( .D(n9080), .CK(clk), .Q(
        wb_dsize_reg_z2[19]), .QN(n4721) );
  DFF_X2 mem_wb_memRdData_q_reg_20_ ( .D(n9078), .CK(clk), .Q(
        wb_dsize_reg_z2[20]), .QN(n4720) );
  DFF_X2 mem_wb_memRdData_q_reg_21_ ( .D(n9077), .CK(clk), .Q(
        wb_dsize_reg_z2[21]), .QN(n4719) );
  DFF_X2 mem_wb_memRdData_q_reg_22_ ( .D(n9076), .CK(clk), .Q(
        wb_dsize_reg_z2[22]), .QN(n4718) );
  DFF_X2 mem_wb_memRdData_q_reg_23_ ( .D(n9075), .CK(clk), .Q(
        wb_dsize_reg_z2[23]), .QN(n4717) );
  DFF_X2 mem_wb_memRdData_q_reg_24_ ( .D(n9074), .CK(clk), .Q(
        wb_dsize_reg_z2[24]), .QN(n4674) );
  DFF_X2 mem_wb_memRdData_q_reg_25_ ( .D(n9073), .CK(clk), .Q(
        wb_dsize_reg_z2[25]), .QN(n4703) );
  DFF_X2 mem_wb_memRdData_q_reg_26_ ( .D(n9072), .CK(clk), .Q(
        wb_dsize_reg_z2[26]), .QN(n4367) );
  DFF_X2 mem_wb_memRdData_q_reg_27_ ( .D(n9071), .CK(clk), .Q(
        wb_dsize_reg_z2[27]), .QN(n4366) );
  DFF_X2 mem_wb_memRdData_q_reg_28_ ( .D(n9070), .CK(clk), .Q(
        wb_dsize_reg_z2[28]), .QN(n4365) );
  DFF_X2 mem_wb_memRdData_q_reg_29_ ( .D(n9069), .CK(clk), .Q(
        wb_dsize_reg_z2[29]), .QN(n4364) );
  DFF_X2 mem_wb_memRdData_q_reg_30_ ( .D(n9067), .CK(clk), .Q(
        wb_dsize_reg_z2[30]), .QN(n4363) );
  DFF_X2 ex_mem_dSize_q_reg_0_ ( .D(n3767), .CK(clk), .Q(dSize[0]) );
  DFF_X2 mem_wb_dSize_q_reg_0_ ( .D(n3766), .CK(clk), .Q(n4105), .QN(n7597) );
  DFF_X2 ex_mem_dSize_q_reg_1_ ( .D(n3765), .CK(clk), .Q(dSize[1]) );
  DFF_X2 mem_wb_dSize_q_reg_1_ ( .D(n3764), .CK(clk), .Q(n4086) );
  DFF_X2 mem_wb_fp_q_reg ( .D(n3762), .CK(clk), .Q(n4106) );
  DFF_X2 mem_wb_rd_q_reg_0_ ( .D(n3760), .CK(clk), .Q(rd[0]) );
  DFF_X2 mem_wb_rd_q_reg_1_ ( .D(n3758), .CK(clk), .Q(rd[1]) );
  DFF_X2 mem_wb_rd_q_reg_2_ ( .D(n3756), .CK(clk), .Q(rd[2]) );
  DFF_X2 mem_wb_rd_q_reg_4_ ( .D(n3749), .CK(clk), .Q(rd[4]) );
  DFF_X2 mem_wb_rd_q_reg_3_ ( .D(n3747), .CK(clk), .Q(rd[3]) );
  DFF_X2 mem_wb_link_q_reg ( .D(n3744), .CK(clk), .Q(n4104), .QN(n7596) );
  DFF_X2 mem_wb_memRd_q_reg ( .D(n3739), .CK(clk), .Q(n4670), .QN(n7595) );
  DFFS_X2 id_ex_instr_q_reg_0_ ( .D(n3695), .CK(clk), .SN(n4877), .QN(n7594)
         );
  DFFS_X2 ex_mem_instr_q_reg_0_ ( .D(n3694), .CK(clk), .SN(n4877), .Q(
        memInstr[0]), .QN(n7593) );
  DFFS_X2 id_ex_instr_q_reg_2_ ( .D(n3691), .CK(clk), .SN(n4877), .Q(n4725), 
        .QN(n7592) );
  DFFS_X2 ex_mem_instr_q_reg_2_ ( .D(n3690), .CK(clk), .SN(n4877), .Q(
        memInstr[2]), .QN(n7591) );
  DFFS_X2 id_ex_instr_q_reg_4_ ( .D(n3687), .CK(clk), .SN(n4877), .Q(n4726), 
        .QN(n7590) );
  DFFS_X2 ex_mem_instr_q_reg_4_ ( .D(n3686), .CK(clk), .SN(n4877), .Q(
        memInstr[4]), .QN(n7589) );
  DFFS_X2 id_ex_not_trap_q_reg ( .D(n3668), .CK(clk), .SN(n4876), .Q(
        not_trap_2), .QN(n4650) );
  DFFS_X2 ex_mem_not_trap_q_reg ( .D(n3667), .CK(clk), .SN(n4876), .Q(
        not_trap_3), .QN(n4716) );
  DFFRS_X2 ifetch_dffa_q_reg_0_ ( .D(n9195), .CK(clk), .RN(n3371), .SN(n3370), 
        .QN(n8902) );
  DFF_X2 mem_wb_reg31Val_q_reg_0_ ( .D(n3662), .CK(clk), .Q(reg31Val_0[0]) );
  DFFRS_X2 ifetch_dffa_q_reg_1_ ( .D(n9196), .CK(clk), .RN(n3369), .SN(n3368), 
        .QN(n8871) );
  DFF_X2 mem_wb_reg31Val_q_reg_1_ ( .D(n3608), .CK(clk), .Q(reg31Val_0[1]) );
  DFF_X2 mem_wb_aluRes_q_reg_22_ ( .D(n3605), .CK(clk), .QN(n7588) );
  DFF_X2 mem_wb_aluRes_q_reg_9_ ( .D(n3602), .CK(clk), .Q(n4615), .QN(n7587)
         );
  DFF_X2 mem_wb_aluRes_q_reg_17_ ( .D(n3599), .CK(clk), .Q(n4616), .QN(n7586)
         );
  DFF_X2 mem_wb_aluRes_q_reg_12_ ( .D(n3596), .CK(clk), .Q(n4624) );
  DFF_X2 mem_wb_aluRes_q_reg_29_ ( .D(n3593), .CK(clk), .Q(n4625) );
  DFF_X2 mem_wb_aluRes_q_reg_8_ ( .D(n3590), .CK(clk), .Q(n4617), .QN(n7585)
         );
  DFF_X2 mem_wb_aluRes_q_reg_25_ ( .D(n3587), .CK(clk), .Q(n4618), .QN(n7584)
         );
  DFF_X2 mem_wb_aluRes_q_reg_18_ ( .D(n3584), .CK(clk), .Q(n4619), .QN(n7583)
         );
  DFF_X2 mem_wb_aluRes_q_reg_27_ ( .D(n3581), .CK(clk), .Q(n4626) );
  DFF_X2 mem_wb_aluRes_q_reg_4_ ( .D(n3578), .CK(clk), .Q(n4620), .QN(n7582)
         );
  DFF_X2 mem_wb_aluRes_q_reg_19_ ( .D(n3575), .CK(clk), .QN(n7581) );
  DFFRS_X2 ifetch_dffa_q_reg_19_ ( .D(n3573), .CK(clk), .RN(n3367), .SN(n3366), 
        .Q(n4603), .QN(n8756) );
  DFFRS_X2 ifetch_dffa_q_reg_20_ ( .D(n3569), .CK(clk), .RN(n3365), .SN(n3364), 
        .Q(n4604), .QN(n8753) );
  DFFRS_X2 ifetch_dffa_q_reg_21_ ( .D(n3565), .CK(clk), .RN(n3363), .SN(n3362), 
        .Q(n4605), .QN(n8750) );
  DFFRS_X2 ifetch_dffa_q_reg_23_ ( .D(n3561), .CK(clk), .RN(n3361), .SN(n3360), 
        .Q(n4606), .QN(n8747) );
  DFFRS_X2 ifetch_dffa_q_reg_24_ ( .D(n3557), .CK(clk), .RN(n3359), .SN(n3358), 
        .Q(n4607), .QN(n8744) );
  DFFRS_X2 ifetch_dffa_q_reg_25_ ( .D(n3553), .CK(clk), .RN(n3357), .SN(n3356), 
        .Q(n4608), .QN(n8741) );
  DFFRS_X2 ifetch_dffa_q_reg_26_ ( .D(n3549), .CK(clk), .RN(n3355), .SN(n3354), 
        .Q(n4609), .QN(n8738) );
  DFFRS_X2 ifetch_dffa_q_reg_27_ ( .D(n3545), .CK(clk), .RN(n3353), .SN(n3352), 
        .Q(n4599), .QN(n8735) );
  DFFRS_X2 ifetch_dffa_q_reg_28_ ( .D(n3541), .CK(clk), .RN(n3351), .SN(n3350), 
        .Q(n4600), .QN(n8732) );
  DFFRS_X2 ifetch_dffa_q_reg_29_ ( .D(n3537), .CK(clk), .RN(n3349), .SN(n3348), 
        .Q(n4601), .QN(n8729) );
  DFFRS_X2 ifetch_dffa_q_reg_30_ ( .D(n3533), .CK(clk), .RN(n3347), .SN(n3346), 
        .Q(n4602), .QN(n8726) );
  DFF_X2 mem_wb_reg31Val_q_reg_30_ ( .D(n3529), .CK(clk), .Q(reg31Val_0[30]), 
        .QN(n4411) );
  DFF_X2 mem_wb_aluRes_q_reg_2_ ( .D(n3526), .CK(clk), .QN(n7580) );
  DFFRS_X2 ifetch_dffa_q_reg_2_ ( .D(n3524), .CK(clk), .RN(n3345), .SN(n3344), 
        .Q(n4556) );
  DFF_X2 mem_wb_reg31Val_q_reg_2_ ( .D(n3520), .CK(clk), .Q(reg31Val_0[2]) );
  DFF_X2 mem_wb_aluRes_q_reg_5_ ( .D(n3517), .CK(clk), .QN(n7579) );
  DFF_X2 mem_wb_aluRes_q_reg_6_ ( .D(n3514), .CK(clk), .QN(n7578) );
  DFF_X2 mem_wb_aluRes_q_reg_14_ ( .D(n3511), .CK(clk), .Q(n4448), .QN(n7577)
         );
  DFFRS_X2 ifetch_dffa_q_reg_15_ ( .D(n3509), .CK(clk), .RN(n3343), .SN(n3342), 
        .Q(n4522), .QN(n8719) );
  DFFRS_X2 ifetch_dffa_q_reg_16_ ( .D(n3505), .CK(clk), .RN(n3341), .SN(n3340), 
        .Q(n4595), .QN(n8716) );
  DFFRS_X2 ifetch_dffa_q_reg_17_ ( .D(n3501), .CK(clk), .RN(n3339), .SN(n3338), 
        .Q(n4596), .QN(n8713) );
  DFFRS_X2 ifetch_dffa_q_reg_18_ ( .D(n3497), .CK(clk), .RN(n3337), .SN(n3336), 
        .Q(n4597), .QN(n8710) );
  DFFRS_X2 ifetch_dffa_q_reg_22_ ( .D(n3493), .CK(clk), .RN(n3335), .SN(n3334), 
        .Q(n4598), .QN(n8707) );
  DFF_X2 mem_wb_reg31Val_q_reg_29_ ( .D(n3489), .CK(clk), .Q(reg31Val_0[29]), 
        .QN(n4409) );
  DFF_X2 mem_wb_reg31Val_q_reg_28_ ( .D(n3488), .CK(clk), .Q(reg31Val_0[28]), 
        .QN(n4410) );
  DFF_X2 mem_wb_aluRes_q_reg_3_ ( .D(n3485), .CK(clk), .QN(n7576) );
  DFFRS_X2 ifetch_dffa_q_reg_3_ ( .D(n3483), .CK(clk), .RN(n3333), .SN(n3332), 
        .Q(n4510), .QN(n8704) );
  DFF_X2 mem_wb_reg31Val_q_reg_3_ ( .D(n3479), .CK(clk), .Q(reg31Val_0[3]) );
  DFFRS_X2 ifetch_dffa_q_reg_4_ ( .D(n3478), .CK(clk), .RN(n3331), .SN(n3330), 
        .Q(n4511), .QN(n8701) );
  DFF_X2 mem_wb_reg31Val_q_reg_4_ ( .D(n3474), .CK(clk), .Q(reg31Val_0[4]) );
  DFFRS_X2 ifetch_dffa_q_reg_5_ ( .D(n3472), .CK(clk), .RN(n3329), .SN(n3328), 
        .Q(n4512), .QN(n8698) );
  DFF_X2 mem_wb_reg31Val_q_reg_5_ ( .D(n3468), .CK(clk), .Q(reg31Val_0[5]) );
  DFFRS_X2 ifetch_dffa_q_reg_6_ ( .D(n3466), .CK(clk), .RN(n3327), .SN(n3326), 
        .Q(n4513), .QN(n8695) );
  DFF_X2 mem_wb_reg31Val_q_reg_6_ ( .D(n3462), .CK(clk), .Q(reg31Val_0[6]) );
  DFFRS_X2 ifetch_dffa_q_reg_7_ ( .D(n3461), .CK(clk), .RN(n3325), .SN(n3324), 
        .Q(n4514), .QN(n8692) );
  DFF_X2 mem_wb_reg31Val_q_reg_7_ ( .D(n3457), .CK(clk), .Q(reg31Val_0[7]) );
  DFFRS_X2 ifetch_dffa_q_reg_8_ ( .D(n3455), .CK(clk), .RN(n3323), .SN(n3322), 
        .Q(n4515), .QN(n8689) );
  DFF_X2 mem_wb_reg31Val_q_reg_8_ ( .D(n3451), .CK(clk), .Q(reg31Val_0[8]), 
        .QN(n4391) );
  DFFRS_X2 ifetch_dffa_q_reg_9_ ( .D(n3450), .CK(clk), .RN(n3321), .SN(n3320), 
        .Q(n4516), .QN(n8686) );
  DFF_X2 mem_wb_reg31Val_q_reg_9_ ( .D(n3446), .CK(clk), .Q(reg31Val_0[9]), 
        .QN(n4390) );
  DFFRS_X2 ifetch_dffa_q_reg_10_ ( .D(n3444), .CK(clk), .RN(n3319), .SN(n3318), 
        .Q(n4517), .QN(n8683) );
  DFF_X2 mem_wb_reg31Val_q_reg_10_ ( .D(n3440), .CK(clk), .Q(reg31Val_0[10])
         );
  DFFRS_X2 ifetch_dffa_q_reg_11_ ( .D(n3439), .CK(clk), .RN(n3317), .SN(n3316), 
        .Q(n4518), .QN(n8680) );
  DFF_X2 mem_wb_reg31Val_q_reg_11_ ( .D(n3435), .CK(clk), .Q(reg31Val_0[11])
         );
  DFFRS_X2 ifetch_dffa_q_reg_12_ ( .D(n3433), .CK(clk), .RN(n3315), .SN(n3314), 
        .Q(n4519), .QN(n8677) );
  DFF_X2 mem_wb_reg31Val_q_reg_12_ ( .D(n3429), .CK(clk), .Q(reg31Val_0[12])
         );
  DFFRS_X2 ifetch_dffa_q_reg_13_ ( .D(n3428), .CK(clk), .RN(n3313), .SN(n3312), 
        .Q(n4520), .QN(n8674) );
  DFF_X2 mem_wb_reg31Val_q_reg_13_ ( .D(n3424), .CK(clk), .Q(reg31Val_0[13])
         );
  DFFRS_X2 ifetch_dffa_q_reg_14_ ( .D(n3422), .CK(clk), .RN(n3311), .SN(n3310), 
        .Q(n4521), .QN(n8671) );
  DFF_X2 mem_wb_reg31Val_q_reg_21_ ( .D(n3418), .CK(clk), .Q(reg31Val_0[21])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_20_ ( .D(n3417), .CK(clk), .Q(reg31Val_0[20])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_19_ ( .D(n3416), .CK(clk), .Q(reg31Val_0[19])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_18_ ( .D(n3415), .CK(clk), .Q(reg31Val_0[18])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_17_ ( .D(n3414), .CK(clk), .Q(reg31Val_0[17])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_16_ ( .D(n3413), .CK(clk), .Q(reg31Val_0[16])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_15_ ( .D(n3411), .CK(clk), .Q(reg31Val_0[15]), 
        .QN(n4441) );
  DFF_X2 mem_wb_reg31Val_q_reg_14_ ( .D(n3410), .CK(clk), .Q(reg31Val_0[14])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_27_ ( .D(n3408), .CK(clk), .Q(reg31Val_0[27]), 
        .QN(n4412) );
  DFF_X2 mem_wb_reg31Val_q_reg_26_ ( .D(n3407), .CK(clk), .Q(reg31Val_0[26]), 
        .QN(n4369) );
  DFF_X2 mem_wb_reg31Val_q_reg_25_ ( .D(n3405), .CK(clk), .Q(reg31Val_0[25])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_24_ ( .D(n3404), .CK(clk), .Q(reg31Val_0[24])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_23_ ( .D(n3402), .CK(clk), .Q(reg31Val_0[23])
         );
  DFF_X2 mem_wb_reg31Val_q_reg_22_ ( .D(n3400), .CK(clk), .Q(reg31Val_0[22])
         );
  DFFRS_X2 ifetch_dffa_q_reg_31_ ( .D(n3397), .CK(clk), .RN(n3309), .SN(n3308), 
        .QN(n8665) );
  DFF_X2 mem_wb_reg31Val_q_reg_31_ ( .D(n3393), .CK(clk), .Q(reg31Val_0[31])
         );
  DFF_X2 mem_wb_aluRes_q_reg_21_ ( .D(n3382), .CK(clk), .QN(n7575) );
  DFFR_X2 if_id_instr_q_reg_30_ ( .D(n3892), .CK(clk), .RN(n4876), .Q(n4554), 
        .QN(n8959) );
  DFFR_X2 if_id_instr_q_reg_26_ ( .D(n3885), .CK(clk), .RN(n4841), .Q(op0_1), 
        .QN(n4323) );
  DFFR_X2 mem_wb_regWr_q_reg ( .D(n3669), .CK(clk), .RN(n4876), .Q(regWr) );
  DFFR_X2 id_ex_fp_q_reg ( .D(n3829), .CK(clk), .RN(n4869), .Q(n4130), .QN(
        n4091) );
  NAND2_X2 U4101 ( .A1(n5481), .A2(n4569), .ZN(n5475) );
  INV_X4 U4102 ( .A(n5481), .ZN(n6333) );
  NAND2_X2 U4103 ( .A1(n5798), .A2(n4593), .ZN(n5799) );
  NAND2_X2 U4104 ( .A1(n6342), .A2(n6341), .ZN(n3896) );
  NAND2_X2 U4105 ( .A1(n6340), .A2(n6339), .ZN(n3895) );
  NAND2_X2 U4106 ( .A1(n6344), .A2(n6343), .ZN(n3897) );
  NAND2_X2 U4107 ( .A1(n6071), .A2(n5882), .ZN(n7841) );
  NAND2_X2 U4108 ( .A1(n7853), .A2(n4558), .ZN(n7125) );
  OAI21_X2 U4109 ( .B1(n6561), .B2(n4169), .A(n6560), .ZN(n6562) );
  OAI21_X2 U4110 ( .B1(n6090), .B2(n6168), .A(n6089), .ZN(n6091) );
  OAI21_X2 U4111 ( .B1(n4110), .B2(n6187), .A(n6188), .ZN(n6431) );
  NAND3_X2 U4112 ( .A1(n6114), .A2(n6115), .A3(n6113), .ZN(n6195) );
  NOR2_X2 U4113 ( .A1(n6159), .A2(n6112), .ZN(n6113) );
  AOI21_X1 U4114 ( .B1(n8349), .B2(n4750), .A(n8348), .ZN(n6112) );
  OAI21_X2 U4115 ( .B1(n6110), .B2(n6190), .A(n6109), .ZN(n6111) );
  OAI21_X2 U4116 ( .B1(n4112), .B2(n6198), .A(n6199), .ZN(n6484) );
  NAND3_X1 U4117 ( .A1(n5344), .A2(n7657), .A3(n4750), .ZN(n5375) );
  NAND3_X1 U4118 ( .A1(n6121), .A2(n4750), .A3(n8348), .ZN(n6118) );
  OAI21_X2 U4119 ( .B1(n6196), .B2(n6195), .A(n6115), .ZN(n6202) );
  OAI21_X2 U4120 ( .B1(n5515), .B2(n5514), .A(n5513), .ZN(n5516) );
  OAI21_X2 U4121 ( .B1(n4252), .B2(n6486), .A(n6510), .ZN(n6511) );
  NAND3_X1 U4122 ( .A1(n6121), .A2(n8364), .A3(n4750), .ZN(n6125) );
  OAI21_X2 U4123 ( .B1(n4114), .B2(n6209), .A(n6210), .ZN(n6739) );
  NAND3_X1 U4124 ( .A1(n6132), .A2(n7723), .A3(n4750), .ZN(n6136) );
  OAI21_X2 U4125 ( .B1(n6130), .B2(n6212), .A(n6129), .ZN(n6131) );
  OAI21_X2 U4126 ( .B1(n4183), .B2(n6220), .A(n6221), .ZN(n6785) );
  OAI21_X2 U4127 ( .B1(n4253), .B2(n6518), .A(n6733), .ZN(n6734) );
  NAND3_X1 U4128 ( .A1(n6143), .A2(n4107), .A3(n7721), .ZN(n6147) );
  OAI21_X2 U4129 ( .B1(n4283), .B2(n6876), .A(n7006), .ZN(n7007) );
  OAI21_X2 U4130 ( .B1(n4293), .B2(n6825), .A(n6844), .ZN(n6845) );
  NAND3_X1 U4131 ( .A1(n4178), .A2(n4753), .A3(n8316), .ZN(n6162) );
  OAI21_X2 U4132 ( .B1(n5584), .B2(n5583), .A(n5538), .ZN(n5539) );
  OAI21_X2 U4133 ( .B1(n6363), .B2(n6362), .A(n6361), .ZN(n6364) );
  OAI21_X2 U4134 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5727) );
  OAI21_X2 U4135 ( .B1(n6747), .B2(n6903), .A(n6746), .ZN(n6912) );
  OAI21_X2 U4136 ( .B1(n4301), .B2(n6770), .A(n6771), .ZN(n6911) );
  NAND3_X2 U4137 ( .A1(n6537), .A2(n4784), .A3(n4561), .ZN(n6538) );
  NAND3_X2 U4138 ( .A1(n4999), .A2(n4998), .A3(n4997), .ZN(n7696) );
  NOR2_X2 U4139 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  NOR2_X2 U4140 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NOR2_X2 U4141 ( .A1(n8968), .A2(n9054), .ZN(n5063) );
  NAND3_X2 U4142 ( .A1(n5109), .A2(n5108), .A3(n5107), .ZN(n7211) );
  NOR2_X2 U4143 ( .A1(n5106), .A2(n5105), .ZN(n5107) );
  NOR2_X2 U4144 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NAND3_X2 U4145 ( .A1(n4985), .A2(n4984), .A3(n4983), .ZN(n7968) );
  NOR2_X2 U4146 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NAND3_X2 U4147 ( .A1(n5104), .A2(n5103), .A3(n5102), .ZN(n5935) );
  NOR2_X2 U4148 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NAND3_X2 U4149 ( .A1(n5177), .A2(n5176), .A3(n5175), .ZN(n7918) );
  NAND3_X2 U4150 ( .A1(n5219), .A2(n4385), .A3(n5218), .ZN(n7659) );
  NAND3_X2 U4151 ( .A1(n5204), .A2(n4382), .A3(n5203), .ZN(n7665) );
  OAI21_X2 U4152 ( .B1(n6563), .B2(n6562), .A(n6564), .ZN(n6708) );
  OAI21_X2 U4153 ( .B1(n6889), .B2(n6888), .A(n7053), .ZN(n7054) );
  OAI21_X2 U4154 ( .B1(n4306), .B2(n6555), .A(n6556), .ZN(n6954) );
  OAI21_X2 U4155 ( .B1(n4316), .B2(n6929), .A(n6930), .ZN(n6968) );
  OAI21_X2 U4156 ( .B1(n4308), .B2(n6908), .A(n6909), .ZN(n7099) );
  OAI21_X2 U4157 ( .B1(n6529), .B2(n6528), .A(n6900), .ZN(n6901) );
  NAND3_X2 U4158 ( .A1(n5097), .A2(n5096), .A3(n5095), .ZN(n7212) );
  NOR2_X2 U4159 ( .A1(n5003), .A2(n5002), .ZN(n5004) );
  NOR2_X2 U4160 ( .A1(n8834), .A2(n4838), .ZN(n5002) );
  OAI21_X2 U4161 ( .B1(n4310), .B2(n7064), .A(n7065), .ZN(n7286) );
  NAND3_X2 U4162 ( .A1(n4994), .A2(n4993), .A3(n4992), .ZN(n7671) );
  NOR2_X2 U4163 ( .A1(n4991), .A2(n4990), .ZN(n4992) );
  NOR3_X2 U4164 ( .A1(n4901), .A2(n4086), .A3(n4105), .ZN(n5171) );
  NOR2_X2 U4165 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NOR2_X2 U4166 ( .A1(n8836), .A2(n4838), .ZN(n5239) );
  NAND3_X1 U4167 ( .A1(n5565), .A2(n4737), .A3(n4750), .ZN(n5561) );
  NAND3_X1 U4168 ( .A1(n5419), .A2(n4737), .A3(n4750), .ZN(n5524) );
  OAI21_X2 U4169 ( .B1(n4752), .B2(n7494), .A(n6096), .ZN(n6098) );
  NAND3_X1 U4170 ( .A1(n5565), .A2(n4750), .A3(n7648), .ZN(n5627) );
  OAI21_X2 U4171 ( .B1(n4211), .B2(n6181), .A(n6182), .ZN(n6405) );
  OAI21_X2 U4172 ( .B1(n4141), .B2(n5705), .A(n5744), .ZN(n5745) );
  OAI21_X2 U4173 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n5694) );
  OAI21_X2 U4174 ( .B1(n4145), .B2(n5569), .A(n5620), .ZN(n5621) );
  OAI21_X2 U4175 ( .B1(n5558), .B2(n5557), .A(n5556), .ZN(n5559) );
  NAND3_X1 U4176 ( .A1(n5419), .A2(n7657), .A3(n4750), .ZN(n5415) );
  OAI21_X2 U4177 ( .B1(n5412), .B2(n5411), .A(n5410), .ZN(n5413) );
  OAI21_X2 U4178 ( .B1(n4752), .B2(n7498), .A(n6116), .ZN(n6117) );
  OAI21_X2 U4179 ( .B1(n4113), .B2(n6203), .A(n6204), .ZN(n6514) );
  NAND3_X2 U4180 ( .A1(n5375), .A2(n5347), .A3(n5346), .ZN(n5376) );
  NOR2_X2 U4181 ( .A1(n6159), .A2(n5345), .ZN(n5346) );
  AOI21_X1 U4182 ( .B1(n7659), .B2(n4750), .A(n7657), .ZN(n5345) );
  OAI21_X2 U4183 ( .B1(n4230), .B2(n6407), .A(n6428), .ZN(n6429) );
  OAI21_X2 U4184 ( .B1(n4260), .B2(n5707), .A(n5740), .ZN(n5741) );
  OAI21_X2 U4185 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5690) );
  OAI21_X2 U4186 ( .B1(n4153), .B2(n5571), .A(n5616), .ZN(n5617) );
  OAI21_X2 U4187 ( .B1(n5554), .B2(n5553), .A(n5552), .ZN(n5555) );
  OAI21_X2 U4188 ( .B1(n4237), .B2(n6433), .A(n6456), .ZN(n6457) );
  OAI21_X2 U4189 ( .B1(n4239), .B2(n6461), .A(n6481), .ZN(n6482) );
  OAI21_X2 U4190 ( .B1(n4249), .B2(n6741), .A(n6761), .ZN(n6762) );
  OAI21_X2 U4191 ( .B1(n4187), .B2(n6019), .A(n6303), .ZN(n6304) );
  OAI21_X2 U4192 ( .B1(n6002), .B2(n6001), .A(n6000), .ZN(n6003) );
  OAI21_X2 U4193 ( .B1(n4212), .B2(n6214), .A(n6215), .ZN(n6764) );
  OAI21_X2 U4194 ( .B1(n4241), .B2(n6766), .A(n6789), .ZN(n6790) );
  OAI21_X2 U4195 ( .B1(n5337), .B2(n5336), .A(n5335), .ZN(n5338) );
  NAND3_X1 U4196 ( .A1(n5344), .A2(n7661), .A3(n4750), .ZN(n5340) );
  OAI21_X2 U4197 ( .B1(n4236), .B2(n6408), .A(n6424), .ZN(n6425) );
  OAI21_X2 U4198 ( .B1(n4228), .B2(n5709), .A(n5736), .ZN(n5737) );
  OAI21_X1 U4199 ( .B1(n5685), .B2(n5684), .A(n5683), .ZN(n5686) );
  OAI21_X2 U4200 ( .B1(n4258), .B2(n5573), .A(n5612), .ZN(n5613) );
  OAI21_X2 U4201 ( .B1(n5550), .B2(n5549), .A(n5548), .ZN(n5551) );
  OAI21_X2 U4202 ( .B1(n4231), .B2(n6434), .A(n6452), .ZN(n6453) );
  NAND3_X2 U4203 ( .A1(n6135), .A2(n6136), .A3(n6134), .ZN(n6217) );
  NOR2_X2 U4204 ( .A1(n6159), .A2(n6133), .ZN(n6134) );
  AOI21_X1 U4205 ( .B1(n4750), .B2(n8326), .A(n7723), .ZN(n6133) );
  OAI21_X2 U4206 ( .B1(n6378), .B2(n6377), .A(n6376), .ZN(n6379) );
  OAI21_X2 U4207 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6508) );
  OAI21_X2 U4208 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(n6756) );
  OAI21_X2 U4209 ( .B1(n4244), .B2(n6742), .A(n6757), .ZN(n6758) );
  OAI21_X2 U4210 ( .B1(n4180), .B2(n6021), .A(n6299), .ZN(n6300) );
  OAI21_X2 U4211 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(n5999) );
  OAI21_X2 U4212 ( .B1(n5370), .B2(n5369), .A(n5368), .ZN(n5405) );
  NAND3_X1 U4213 ( .A1(n6143), .A2(n7723), .A3(n4107), .ZN(n6140) );
  OAI21_X2 U4214 ( .B1(n4184), .B2(n6225), .A(n6226), .ZN(n6817) );
  OAI21_X2 U4215 ( .B1(n4256), .B2(n6819), .A(n6831), .ZN(n6832) );
  OAI21_X2 U4216 ( .B1(n4250), .B2(n6767), .A(n6782), .ZN(n6783) );
  OAI21_X2 U4217 ( .B1(n4242), .B2(n6792), .A(n6808), .ZN(n6809) );
  OAI21_X2 U4218 ( .B1(n4218), .B2(n6409), .A(n6420), .ZN(n6421) );
  OAI21_X2 U4219 ( .B1(n4194), .B2(n5711), .A(n5732), .ZN(n5733) );
  OAI21_X2 U4220 ( .B1(n5681), .B2(n5680), .A(n5679), .ZN(n5682) );
  OAI21_X2 U4221 ( .B1(n4221), .B2(n6488), .A(n6500), .ZN(n6501) );
  OAI21_X2 U4222 ( .B1(n4217), .B2(n5575), .A(n5608), .ZN(n5609) );
  OAI21_X2 U4223 ( .B1(n5546), .B2(n5545), .A(n5544), .ZN(n5547) );
  OAI21_X2 U4224 ( .B1(n4219), .B2(n6435), .A(n6448), .ZN(n6449) );
  NAND3_X2 U4225 ( .A1(n6146), .A2(n6147), .A3(n6145), .ZN(n6228) );
  NOR2_X2 U4226 ( .A1(n6159), .A2(n6144), .ZN(n6145) );
  AOI21_X1 U4227 ( .B1(n4750), .B2(n7722), .A(n7721), .ZN(n6144) );
  OAI21_X2 U4228 ( .B1(n4115), .B2(n6231), .A(n6232), .ZN(n6828) );
  OAI21_X2 U4229 ( .B1(n4263), .B2(n6830), .A(n6866), .ZN(n6867) );
  OAI21_X2 U4230 ( .B1(n4220), .B2(n6463), .A(n6473), .ZN(n6474) );
  OAI21_X2 U4231 ( .B1(n4223), .B2(n6743), .A(n6753), .ZN(n6754) );
  OAI21_X2 U4232 ( .B1(n4196), .B2(n6023), .A(n6295), .ZN(n6296) );
  OAI21_X2 U4233 ( .B1(n5994), .B2(n5993), .A(n5992), .ZN(n5995) );
  OAI21_X2 U4234 ( .B1(n5386), .B2(n5385), .A(n5384), .ZN(n5400) );
  OAI21_X2 U4235 ( .B1(n4185), .B2(n6236), .A(n6237), .ZN(n6870) );
  OAI21_X2 U4236 ( .B1(n4224), .B2(n6768), .A(n6778), .ZN(n6779) );
  OAI21_X2 U4237 ( .B1(n5306), .B2(n5495), .A(n5294), .ZN(n5314) );
  OAI21_X2 U4238 ( .B1(n4190), .B2(n6410), .A(n6437), .ZN(n6438) );
  OAI21_X2 U4239 ( .B1(n4201), .B2(n5713), .A(n5728), .ZN(n5729) );
  OAI21_X2 U4240 ( .B1(n5677), .B2(n5676), .A(n5675), .ZN(n5678) );
  OAI21_X2 U4241 ( .B1(n4227), .B2(n6489), .A(n6495), .ZN(n6496) );
  OAI21_X2 U4242 ( .B1(n4199), .B2(n5577), .A(n5604), .ZN(n5605) );
  OAI21_X2 U4243 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5543) );
  OAI21_X2 U4244 ( .B1(n4264), .B2(n6874), .A(n7002), .ZN(n7003) );
  OAI21_X2 U4245 ( .B1(n6863), .B2(n6862), .A(n6861), .ZN(n6864) );
  OAI21_X2 U4246 ( .B1(n6153), .B2(n6234), .A(n6152), .ZN(n6154) );
  OAI21_X2 U4247 ( .B1(n4213), .B2(n6242), .A(n6243), .ZN(n6995) );
  OAI21_X2 U4248 ( .B1(n6997), .B2(n4266), .A(n7031), .ZN(n7032) );
  OAI21_X2 U4249 ( .B1(n4284), .B2(n7005), .A(n7022), .ZN(n7023) );
  OAI21_X2 U4250 ( .B1(n4226), .B2(n6464), .A(n6469), .ZN(n6470) );
  OAI21_X2 U4251 ( .B1(n5970), .B2(n5434), .A(n5393), .ZN(n5394) );
  OAI21_X2 U4252 ( .B1(n4290), .B2(n6744), .A(n6749), .ZN(n6750) );
  OAI21_X2 U4253 ( .B1(n5990), .B2(n5989), .A(n5988), .ZN(n5991) );
  OAI21_X2 U4254 ( .B1(n4297), .B2(n7001), .A(n7026), .ZN(n7027) );
  OAI21_X2 U4255 ( .B1(n6240), .B2(n6239), .A(n6156), .ZN(n6246) );
  NAND3_X2 U4256 ( .A1(n6161), .A2(n6162), .A3(n6160), .ZN(n6245) );
  NOR2_X2 U4257 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  AOI21_X2 U4258 ( .B1(n8304), .B2(n4753), .A(n8316), .ZN(n6158) );
  OAI21_X2 U4259 ( .B1(n4186), .B2(n6247), .A(n6248), .ZN(n7034) );
  OAI21_X2 U4260 ( .B1(n7036), .B2(n4248), .A(n7249), .ZN(n7250) );
  OAI21_X2 U4261 ( .B1(n7039), .B2(n4288), .A(n7260), .ZN(n7261) );
  OAI21_X2 U4262 ( .B1(n4291), .B2(n6769), .A(n6774), .ZN(n6775) );
  OAI21_X2 U4263 ( .B1(n4292), .B2(n6794), .A(n6799), .ZN(n6800) );
  OAI21_X2 U4264 ( .B1(n4285), .B2(n7009), .A(n7017), .ZN(n7018) );
  OAI21_X2 U4265 ( .B1(n6467), .B2(n6558), .A(n6466), .ZN(n6567) );
  OAI21_X2 U4266 ( .B1(n4299), .B2(n6490), .A(n6491), .ZN(n6566) );
  OAI21_X2 U4267 ( .B1(n6541), .B2(n6540), .A(n6417), .ZN(n6418) );
  NAND3_X2 U4268 ( .A1(n7255), .A2(n7722), .A3(n4100), .ZN(n7327) );
  NOR2_X2 U4269 ( .A1(n8999), .A2(n4837), .ZN(n4973) );
  NOR2_X2 U4270 ( .A1(n8962), .A2(n4838), .ZN(n4972) );
  OAI21_X2 U4271 ( .B1(n4298), .B2(n6465), .A(n6466), .ZN(n6558) );
  OAI21_X2 U4272 ( .B1(n4303), .B2(n6826), .A(n6827), .ZN(n6922) );
  NOR2_X2 U4273 ( .A1(n9042), .A2(n4836), .ZN(n5068) );
  OAI21_X2 U4274 ( .B1(n5602), .B2(n5601), .A(n5600), .ZN(n5603) );
  OAI21_X2 U4275 ( .B1(n6923), .B2(n6922), .A(n6827), .ZN(n6932) );
  OAI21_X2 U4276 ( .B1(n6289), .B2(n6288), .A(n6287), .ZN(n6290) );
  OAI21_X2 U4277 ( .B1(n6772), .B2(n6911), .A(n6771), .ZN(n6890) );
  INV_X4 U4278 ( .A(n4754), .ZN(n4753) );
  NOR2_X2 U4279 ( .A1(n5036), .A2(n4443), .ZN(n5037) );
  NOR2_X2 U4280 ( .A1(n5042), .A2(n4274), .ZN(n5043) );
  NOR2_X2 U4281 ( .A1(n5261), .A2(n4392), .ZN(n5262) );
  NOR2_X2 U4282 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  NOR2_X2 U4283 ( .A1(n8933), .A2(n9054), .ZN(n5272) );
  NAND3_X2 U4284 ( .A1(n5054), .A2(n5053), .A3(n5052), .ZN(n6322) );
  NOR2_X2 U4285 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  NAND3_X2 U4286 ( .A1(n5017), .A2(n5016), .A3(n5015), .ZN(n7906) );
  NOR2_X2 U4287 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  NOR2_X2 U4288 ( .A1(n8943), .A2(n9054), .ZN(n5268) );
  NAND3_X2 U4289 ( .A1(n5049), .A2(n5048), .A3(n5047), .ZN(n5267) );
  NOR2_X2 U4290 ( .A1(n5046), .A2(n5045), .ZN(n5047) );
  NOR2_X2 U4291 ( .A1(n5246), .A2(n4444), .ZN(n5247) );
  OAI21_X1 U4292 ( .B1(n6527), .B2(n4169), .A(n6526), .ZN(n6528) );
  NOR2_X2 U4293 ( .A1(n5039), .A2(n4272), .ZN(n5040) );
  NOR2_X2 U4294 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  NOR2_X2 U4295 ( .A1(n8970), .A2(n4838), .ZN(n5059) );
  INV_X4 U4296 ( .A(n5702), .ZN(n6159) );
  NOR2_X2 U4297 ( .A1(n5236), .A2(n4273), .ZN(n5237) );
  NOR2_X2 U4298 ( .A1(n9050), .A2(n9047), .ZN(n4894) );
  NOR2_X2 U4299 ( .A1(n9048), .A2(n9051), .ZN(n4895) );
  NOR2_X2 U4300 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NOR2_X2 U4301 ( .A1(n8935), .A2(n9054), .ZN(n5227) );
  NOR2_X2 U4302 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  NAND3_X2 U4303 ( .A1(n5215), .A2(n4383), .A3(n5214), .ZN(n7663) );
  OAI22_X2 U4304 ( .A1(n7552), .A2(n8631), .B1(n8632), .B2(n8601), .ZN(n8561)
         );
  OAI21_X2 U4305 ( .B1(n7702), .B2(n7701), .A(n6030), .ZN(n7991) );
  OAI21_X2 U4306 ( .B1(n4166), .B2(n6029), .A(n6282), .ZN(n6283) );
  OAI22_X2 U4307 ( .A1(n7514), .A2(n8640), .B1(n8641), .B2(n8593), .ZN(n8547)
         );
  NAND3_X2 U4308 ( .A1(n5793), .A2(n4440), .A3(n5792), .ZN(n8448) );
  OAI21_X2 U4309 ( .B1(n7689), .B2(n7688), .A(n5718), .ZN(n7910) );
  OAI21_X2 U4310 ( .B1(n4305), .B2(n5717), .A(n5719), .ZN(n7909) );
  OAI21_X2 U4311 ( .B1(n4314), .B2(n6546), .A(n6547), .ZN(n7079) );
  NAND3_X2 U4312 ( .A1(n5087), .A2(n4429), .A3(n5086), .ZN(n8364) );
  OAI21_X2 U4313 ( .B1(n6565), .B2(n6708), .A(n6564), .ZN(n7199) );
  OAI21_X2 U4314 ( .B1(n4307), .B2(n6572), .A(n6573), .ZN(n7198) );
  NAND3_X2 U4315 ( .A1(n5787), .A2(n5786), .A3(n5785), .ZN(n8348) );
  NAND3_X2 U4316 ( .A1(n5057), .A2(n5056), .A3(n5055), .ZN(n5767) );
  OAI21_X2 U4317 ( .B1(n4265), .B2(n5581), .A(n5596), .ZN(n7710) );
  OAI21_X2 U4318 ( .B1(n7889), .B2(n7890), .A(n5594), .ZN(n5595) );
  NOR2_X2 U4319 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  NOR2_X2 U4320 ( .A1(n8974), .A2(n9054), .ZN(n5199) );
  NAND3_X2 U4321 ( .A1(n5795), .A2(n4436), .A3(n5794), .ZN(n8460) );
  OAI21_X2 U4322 ( .B1(n8464), .B2(n8463), .A(n6530), .ZN(n7227) );
  OAI21_X2 U4323 ( .B1(n4313), .B2(n6537), .A(n6538), .ZN(n7226) );
  OAI21_X2 U4324 ( .B1(n7066), .B2(n7286), .A(n7065), .ZN(n7235) );
  OAI21_X2 U4325 ( .B1(n7051), .B2(n7050), .A(n7236), .ZN(n7237) );
  NAND3_X2 U4326 ( .A1(n7276), .A2(n7275), .A3(n7274), .ZN(n7277) );
  AOI22_X2 U4327 ( .A1(n7720), .A2(n8610), .B1(n8584), .B2(n8585), .ZN(n8539)
         );
  NAND3_X2 U4328 ( .A1(n5020), .A2(n5019), .A3(n5018), .ZN(n7682) );
  OAI21_X2 U4329 ( .B1(n6931), .B2(n6968), .A(n6930), .ZN(n7303) );
  OAI21_X2 U4330 ( .B1(n4309), .B2(n6939), .A(n6940), .ZN(n7302) );
  OAI21_X2 U4331 ( .B1(n6910), .B2(n7099), .A(n6909), .ZN(n7313) );
  OAI21_X2 U4332 ( .B1(n4315), .B2(n6916), .A(n6917), .ZN(n7312) );
  OAI21_X2 U4333 ( .B1(n7372), .B2(n7371), .A(n7370), .ZN(n7373) );
  NOR2_X2 U4334 ( .A1(n7576), .A2(n4742), .ZN(n5129) );
  NOR2_X2 U4335 ( .A1(n7585), .A2(n4742), .ZN(n5026) );
  NOR2_X2 U4336 ( .A1(n7587), .A2(n4742), .ZN(n5022) );
  NOR2_X2 U4337 ( .A1(n7605), .A2(n4742), .ZN(n5007) );
  NOR2_X2 U4338 ( .A1(n7475), .A2(n6046), .ZN(n5479) );
  NAND3_X2 U4339 ( .A1(n4927), .A2(n4438), .A3(n4926), .ZN(n7641) );
  NAND3_X2 U4340 ( .A1(n5789), .A2(n4434), .A3(n5788), .ZN(n8349) );
  NOR2_X2 U4341 ( .A1(n4956), .A2(n4955), .ZN(n4957) );
  NOR2_X2 U4342 ( .A1(n8831), .A2(n4838), .ZN(n4955) );
  NAND3_X2 U4343 ( .A1(n5791), .A2(n4435), .A3(n5790), .ZN(n7895) );
  NAND3_X2 U4344 ( .A1(n5784), .A2(n4433), .A3(n5783), .ZN(n8336) );
  NAND3_X2 U4345 ( .A1(n6082), .A2(n6081), .A3(n6080), .ZN(n7726) );
  NAND3_X2 U4346 ( .A1(n5014), .A2(n5013), .A3(n5012), .ZN(n8479) );
  NOR2_X2 U4347 ( .A1(n5011), .A2(n5010), .ZN(n5012) );
  NAND3_X2 U4348 ( .A1(n4921), .A2(n4920), .A3(n4919), .ZN(n7634) );
  AOI21_X2 U4349 ( .B1(n7288), .B2(n7896), .A(n7544), .ZN(n7289) );
  NOR3_X2 U4350 ( .A1(n7433), .A2(n7432), .A3(n7431), .ZN(n7434) );
  NAND3_X2 U4351 ( .A1(n4939), .A2(n4938), .A3(n4937), .ZN(regWrData[0]) );
  AOI22_X2 U4352 ( .A1(wb_dsize_reg_z2[0]), .A2(n5209), .B1(n5171), .B2(
        wb_dsize_reg_z2[24]), .ZN(n4937) );
  AOI21_X2 U4353 ( .B1(reg31Val_0[0]), .B2(n4741), .A(n4935), .ZN(n4939) );
  NAND3_X2 U4354 ( .A1(n4947), .A2(n4946), .A3(n4945), .ZN(regWrData[1]) );
  AOI21_X2 U4355 ( .B1(reg31Val_0[1]), .B2(n4741), .A(n4944), .ZN(n4947) );
  NAND3_X2 U4356 ( .A1(n4943), .A2(n4942), .A3(n4941), .ZN(regWrData[2]) );
  AOI21_X2 U4357 ( .B1(reg31Val_0[2]), .B2(n4741), .A(n4940), .ZN(n4943) );
  NAND3_X2 U4358 ( .A1(n5174), .A2(n5173), .A3(n5172), .ZN(regWrData[4]) );
  AOI21_X2 U4359 ( .B1(reg31Val_0[4]), .B2(n4741), .A(n5169), .ZN(n5174) );
  NAND3_X2 U4360 ( .A1(n4980), .A2(n4979), .A3(n4978), .ZN(regWrData[5]) );
  AOI21_X2 U4361 ( .B1(reg31Val_0[5]), .B2(n4741), .A(n4977), .ZN(n4980) );
  NAND3_X2 U4362 ( .A1(n4971), .A2(n4970), .A3(n4969), .ZN(regWrData[6]) );
  AOI21_X2 U4363 ( .B1(reg31Val_0[6]), .B2(n4741), .A(n4968), .ZN(n4971) );
  NAND3_X2 U4364 ( .A1(n4989), .A2(n4988), .A3(n4987), .ZN(regWrData[7]) );
  AOI21_X2 U4365 ( .B1(reg31Val_0[7]), .B2(n4741), .A(n4986), .ZN(n4989) );
  NAND3_X2 U4366 ( .A1(n4962), .A2(n4961), .A3(n4375), .ZN(regWrData[26]) );
  NAND3_X2 U4367 ( .A1(n4960), .A2(n4959), .A3(n4420), .ZN(regWrData[28]) );
  NAND3_X2 U4368 ( .A1(n5001), .A2(n5000), .A3(n4421), .ZN(regWrData[30]) );
  NAND3_X2 U4369 ( .A1(n4949), .A2(n4948), .A3(n4428), .ZN(regWrData[31]) );
  OAI21_X2 U4370 ( .B1(n4754), .B2(n7553), .A(n5700), .ZN(n5703) );
  OAI21_X2 U4371 ( .B1(n4754), .B2(n7549), .A(n7192), .ZN(n5567) );
  OAI21_X2 U4372 ( .B1(n5563), .B2(n5562), .A(n5561), .ZN(n5564) );
  NAND3_X2 U4373 ( .A1(n6104), .A2(n6105), .A3(n6103), .ZN(n6184) );
  NOR2_X2 U4374 ( .A1(n6159), .A2(n6102), .ZN(n6103) );
  AOI21_X2 U4375 ( .B1(n7895), .B2(n4750), .A(n8448), .ZN(n6102) );
  OAI21_X2 U4376 ( .B1(n6100), .B2(n6179), .A(n6099), .ZN(n6101) );
  NAND3_X2 U4377 ( .A1(n6094), .A2(n6095), .A3(n6093), .ZN(n6174) );
  NOR2_X2 U4378 ( .A1(n6159), .A2(n6092), .ZN(n6093) );
  AOI21_X2 U4379 ( .B1(n7726), .B2(n4750), .A(n8460), .ZN(n6092) );
  OAI21_X2 U4380 ( .B1(n7512), .B2(n4752), .A(n4088), .ZN(n5421) );
  NAND3_X2 U4381 ( .A1(n6015), .A2(n6083), .A3(n6014), .ZN(n6084) );
  NOR2_X2 U4382 ( .A1(n6159), .A2(n6013), .ZN(n6014) );
  AOI21_X2 U4383 ( .B1(n7634), .B2(n4750), .A(n7641), .ZN(n6013) );
  OAI21_X2 U4384 ( .B1(n5753), .B2(n5752), .A(n5751), .ZN(n6008) );
  OAI21_X2 U4385 ( .B1(n4752), .B2(n7553), .A(n5748), .ZN(n5750) );
  OAI21_X2 U4386 ( .B1(n5629), .B2(n5628), .A(n5627), .ZN(n5695) );
  OAI21_X2 U4387 ( .B1(n4752), .B2(n7549), .A(n5624), .ZN(n5626) );
  OAI21_X2 U4388 ( .B1(n6185), .B2(n6184), .A(n6105), .ZN(n6191) );
  OAI21_X2 U4389 ( .B1(n4752), .B2(n7495), .A(n6106), .ZN(n6108) );
  OAI21_X2 U4390 ( .B1(n6085), .B2(n6084), .A(n6083), .ZN(n6169) );
  OAI21_X2 U4391 ( .B1(n4752), .B2(n7551), .A(n6086), .ZN(n6088) );
  OAI21_X2 U4392 ( .B1(n4144), .B2(n5527), .A(n5556), .ZN(n5557) );
  OAI21_X2 U4393 ( .B1(n5519), .B2(n5518), .A(n5517), .ZN(n5520) );
  OAI21_X2 U4394 ( .B1(n4210), .B2(n6177), .A(n6178), .ZN(n6366) );
  OAI21_X2 U4395 ( .B1(n6172), .B2(n6307), .A(n6171), .ZN(n6173) );
  OAI21_X2 U4396 ( .B1(n6189), .B2(n6431), .A(n6188), .ZN(n6460) );
  OAI21_X2 U4397 ( .B1(n4111), .B2(n6192), .A(n6193), .ZN(n6459) );
  OAI21_X2 U4398 ( .B1(n4143), .B2(n5423), .A(n5517), .ZN(n5518) );
  OAI21_X2 U4399 ( .B1(n4148), .B2(n6017), .A(n6165), .ZN(n6166) );
  OAI21_X2 U4400 ( .B1(n4147), .B2(n5754), .A(n6004), .ZN(n6005) );
  OAI21_X2 U4401 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(n5747) );
  OAI21_X2 U4402 ( .B1(n4146), .B2(n5630), .A(n5691), .ZN(n5692) );
  OAI21_X2 U4403 ( .B1(n5622), .B2(n5621), .A(n5620), .ZN(n5623) );
  OAI21_X2 U4404 ( .B1(n5377), .B2(n5376), .A(n5375), .ZN(n5414) );
  OAI21_X2 U4405 ( .B1(n7513), .B2(n4752), .A(n5378), .ZN(n5379) );
  OAI21_X2 U4406 ( .B1(n6167), .B2(n6166), .A(n6165), .ZN(n6308) );
  OAI21_X2 U4407 ( .B1(n4149), .B2(n6170), .A(n6171), .ZN(n6307) );
  OAI21_X2 U4408 ( .B1(n6404), .B2(n6403), .A(n6402), .ZN(n6427) );
  OAI21_X2 U4409 ( .B1(n4161), .B2(n5529), .A(n5552), .ZN(n5553) );
  NAND3_X2 U4410 ( .A1(n6124), .A2(n6125), .A3(n6123), .ZN(n6206) );
  NOR2_X2 U4411 ( .A1(n6159), .A2(n6122), .ZN(n6123) );
  AOI21_X2 U4412 ( .B1(n4753), .B2(n8364), .A(n8336), .ZN(n6122) );
  OAI21_X2 U4413 ( .B1(n6119), .B2(n6201), .A(n6118), .ZN(n6120) );
  OAI21_X2 U4414 ( .B1(n6205), .B2(n6514), .A(n6204), .ZN(n6740) );
  OAI21_X2 U4415 ( .B1(n4235), .B2(n6369), .A(n6402), .ZN(n6403) );
  OAI21_X2 U4416 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(n6480) );
  OAI21_X2 U4417 ( .B1(n4164), .B2(n5425), .A(n5513), .ZN(n5514) );
  OAI21_X2 U4418 ( .B1(n5408), .B2(n5407), .A(n5406), .ZN(n5409) );
  OAI21_X2 U4419 ( .B1(n4243), .B2(n6516), .A(n6736), .ZN(n6737) );
  OAI21_X2 U4420 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6513) );
  OAI21_X2 U4421 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(n6760) );
  OAI21_X2 U4422 ( .B1(n4179), .B2(n5756), .A(n6000), .ZN(n6001) );
  OAI21_X2 U4423 ( .B1(n5742), .B2(n5741), .A(n5740), .ZN(n5743) );
  OAI21_X2 U4424 ( .B1(n4154), .B2(n5632), .A(n5687), .ZN(n5688) );
  OAI21_X2 U4425 ( .B1(n5618), .B2(n5617), .A(n5616), .ZN(n5619) );
  OAI21_X2 U4426 ( .B1(n5373), .B2(n5372), .A(n5371), .ZN(n5374) );
  OAI21_X2 U4427 ( .B1(n5380), .B2(n4151), .A(n5410), .ZN(n5411) );
  NAND3_X2 U4428 ( .A1(n6132), .A2(n8364), .A3(n4750), .ZN(n6129) );
  OAI21_X2 U4429 ( .B1(n6207), .B2(n6206), .A(n6125), .ZN(n6213) );
  OAI21_X2 U4430 ( .B1(n4233), .B2(n6309), .A(n6370), .ZN(n6371) );
  OAI21_X2 U4431 ( .B1(n6305), .B2(n6304), .A(n6303), .ZN(n6306) );
  OAI21_X2 U4432 ( .B1(n5349), .B2(n4103), .A(n5371), .ZN(n5372) );
  OAI21_X2 U4433 ( .B1(n6401), .B2(n6400), .A(n6399), .ZN(n6423) );
  OAI21_X2 U4434 ( .B1(n4245), .B2(n5531), .A(n5548), .ZN(n5549) );
  OAI21_X2 U4435 ( .B1(n4240), .B2(n6487), .A(n6505), .ZN(n6506) );
  OAI21_X2 U4436 ( .B1(n6216), .B2(n6764), .A(n6215), .ZN(n6786) );
  OAI21_X2 U4437 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6812) );
  OAI21_X2 U4438 ( .B1(n6787), .B2(n4255), .A(n6813), .ZN(n6814) );
  OAI21_X2 U4439 ( .B1(n4234), .B2(n6375), .A(n6399), .ZN(n6400) );
  OAI21_X2 U4440 ( .B1(n7515), .B2(n4752), .A(n5322), .ZN(n5323) );
  OAI21_X2 U4441 ( .B1(n6454), .B2(n6453), .A(n6452), .ZN(n6476) );
  OAI21_X2 U4442 ( .B1(n4238), .B2(n6462), .A(n6477), .ZN(n6478) );
  NAND3_X2 U4443 ( .A1(n5299), .A2(n7661), .A3(n4750), .ZN(n5319) );
  OAI21_X2 U4444 ( .B1(n4269), .B2(n5427), .A(n5509), .ZN(n5510) );
  OAI21_X2 U4445 ( .B1(n5403), .B2(n5402), .A(n5401), .ZN(n5404) );
  OAI21_X2 U4446 ( .B1(n4261), .B2(n5758), .A(n5996), .ZN(n5997) );
  OAI21_X2 U4447 ( .B1(n5738), .B2(n5737), .A(n5736), .ZN(n5739) );
  OAI21_X2 U4448 ( .B1(n4214), .B2(n5634), .A(n5683), .ZN(n5684) );
  OAI21_X2 U4449 ( .B1(n5614), .B2(n5613), .A(n5612), .ZN(n5615) );
  OAI21_X2 U4450 ( .B1(n5382), .B2(n4167), .A(n5406), .ZN(n5407) );
  OAI21_X2 U4451 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6781) );
  OAI21_X2 U4452 ( .B1(n4188), .B2(n6311), .A(n6376), .ZN(n6377) );
  OAI21_X2 U4453 ( .B1(n6301), .B2(n6300), .A(n6299), .ZN(n6302) );
  OAI21_X2 U4454 ( .B1(n5351), .B2(n4163), .A(n5368), .ZN(n5369) );
  OAI21_X2 U4455 ( .B1(n5333), .B2(n5332), .A(n5331), .ZN(n5334) );
  OAI21_X2 U4456 ( .B1(n5297), .B2(n5296), .A(n5295), .ZN(n5298) );
  NAND3_X2 U4457 ( .A1(n5702), .A2(n5319), .A3(n5302), .ZN(n5320) );
  NOR2_X2 U4458 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  AOI21_X2 U4459 ( .B1(n4753), .B2(n7661), .A(n7663), .ZN(n5301) );
  NOR2_X2 U4460 ( .A1(n7661), .A2(n4750), .ZN(n5300) );
  OAI21_X2 U4461 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(n6419) );
  OAI21_X2 U4462 ( .B1(n4192), .B2(n5533), .A(n5544), .ZN(n5545) );
  OAI21_X2 U4463 ( .B1(n5507), .B2(n5506), .A(n5505), .ZN(n5508) );
  OAI21_X2 U4464 ( .B1(n4251), .B2(n6821), .A(n6835), .ZN(n6836) );
  OAI21_X2 U4465 ( .B1(n6810), .B2(n6809), .A(n6808), .ZN(n6811) );
  OAI21_X2 U4466 ( .B1(n6141), .B2(n6223), .A(n6140), .ZN(n6142) );
  OAI21_X2 U4467 ( .B1(n6227), .B2(n6817), .A(n6226), .ZN(n6829) );
  OAI21_X2 U4468 ( .B1(n4189), .B2(n6381), .A(n6396), .ZN(n6397) );
  OAI21_X2 U4469 ( .B1(n5317), .B2(n5316), .A(n5315), .ZN(n5318) );
  OAI21_X2 U4470 ( .B1(n5324), .B2(n4150), .A(n5335), .ZN(n5336) );
  OAI21_X2 U4471 ( .B1(n6450), .B2(n6449), .A(n6448), .ZN(n6472) );
  OAI21_X2 U4472 ( .B1(n4117), .B2(n6823), .A(n6839), .ZN(n6840) );
  OAI21_X2 U4473 ( .B1(n4216), .B2(n5429), .A(n5505), .ZN(n5506) );
  OAI21_X2 U4474 ( .B1(n4222), .B2(n6520), .A(n6730), .ZN(n6731) );
  OAI21_X2 U4475 ( .B1(n6502), .B2(n6501), .A(n6500), .ZN(n6503) );
  OAI21_X2 U4476 ( .B1(n6732), .B2(n6731), .A(n6730), .ZN(n6752) );
  OAI21_X2 U4477 ( .B1(n4195), .B2(n5760), .A(n5992), .ZN(n5993) );
  OAI21_X2 U4478 ( .B1(n5734), .B2(n5733), .A(n5732), .ZN(n5735) );
  OAI21_X2 U4479 ( .B1(n4193), .B2(n5636), .A(n5679), .ZN(n5680) );
  OAI21_X2 U4480 ( .B1(n5610), .B2(n5609), .A(n5608), .ZN(n5611) );
  OAI21_X2 U4481 ( .B1(n4157), .B2(n5383), .A(n5401), .ZN(n5402) );
  OAI21_X2 U4482 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(n6860) );
  OAI21_X2 U4483 ( .B1(n4257), .B2(n6834), .A(n6861), .ZN(n6862) );
  OAI21_X2 U4484 ( .B1(n6229), .B2(n6228), .A(n6147), .ZN(n6235) );
  OAI21_X2 U4485 ( .B1(n4232), .B2(n6872), .A(n6998), .ZN(n6999) );
  OAI21_X2 U4486 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6869) );
  OAI21_X2 U4487 ( .B1(n4181), .B2(n6313), .A(n6382), .ZN(n6383) );
  OAI21_X2 U4488 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(n6298) );
  OAI21_X2 U4489 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6802) );
  OAI21_X2 U4490 ( .B1(n4116), .B2(n6793), .A(n6803), .ZN(n6804) );
  OAI21_X2 U4491 ( .B1(n5353), .B2(n4158), .A(n5384), .ZN(n5385) );
  OAI21_X2 U4492 ( .B1(n5669), .B2(n5356), .A(n5328), .ZN(n5329) );
  OAI21_X2 U4493 ( .B1(n4142), .B2(n5304), .A(n5315), .ZN(n5316) );
  OAI21_X2 U4494 ( .B1(n6841), .B2(n6840), .A(n6839), .ZN(n6855) );
  OAI21_X2 U4495 ( .B1(n4123), .B2(n6838), .A(n6856), .ZN(n6857) );
  OAI21_X2 U4496 ( .B1(n4198), .B2(n5535), .A(n5540), .ZN(n5541) );
  OAI21_X2 U4497 ( .B1(n5503), .B2(n5502), .A(n5501), .ZN(n5504) );
  OAI21_X2 U4498 ( .B1(n6439), .B2(n6438), .A(n6437), .ZN(n6440) );
  OAI21_X2 U4499 ( .B1(n4225), .B2(n6436), .A(n6444), .ZN(n6445) );
  OAI21_X2 U4500 ( .B1(n6238), .B2(n6870), .A(n6237), .ZN(n6996) );
  OAI21_X2 U4501 ( .B1(n7000), .B2(n6999), .A(n6998), .ZN(n7030) );
  OAI21_X2 U4502 ( .B1(n4182), .B2(n6387), .A(n6411), .ZN(n6412) );
  NAND3_X2 U4503 ( .A1(n5280), .A2(n4750), .A3(n5796), .ZN(n5281) );
  OAI21_X2 U4504 ( .B1(n5313), .B2(n5312), .A(n5311), .ZN(n5330) );
  OAI21_X2 U4505 ( .B1(n5326), .B2(n4165), .A(n5331), .ZN(n5332) );
  OAI21_X2 U4506 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n6468) );
  OAI21_X2 U4507 ( .B1(n4197), .B2(n5431), .A(n5501), .ZN(n5502) );
  OAI21_X2 U4508 ( .B1(n6497), .B2(n6496), .A(n6495), .ZN(n6498) );
  OAI21_X2 U4509 ( .B1(n4289), .B2(n6522), .A(n6727), .ZN(n6728) );
  OAI21_X2 U4510 ( .B1(n6729), .B2(n6728), .A(n6727), .ZN(n6748) );
  OAI21_X2 U4511 ( .B1(n5730), .B2(n5729), .A(n5728), .ZN(n5731) );
  OAI21_X2 U4512 ( .B1(n4202), .B2(n5762), .A(n5988), .ZN(n5989) );
  OAI21_X2 U4513 ( .B1(n5606), .B2(n5605), .A(n5604), .ZN(n5607) );
  OAI21_X2 U4514 ( .B1(n4200), .B2(n5638), .A(n5675), .ZN(n5676) );
  OAI21_X2 U4515 ( .B1(n5367), .B2(n5366), .A(n5365), .ZN(n5398) );
  OAI21_X2 U4516 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7259) );
  OAI21_X2 U4517 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6294) );
  OAI21_X2 U4518 ( .B1(n4204), .B2(n6315), .A(n6388), .ZN(n6389) );
  OAI21_X2 U4519 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n6798) );
  NAND3_X2 U4520 ( .A1(n5072), .A2(n7540), .A3(n5071), .ZN(n5077) );
  NOR2_X2 U4521 ( .A1(n7988), .A2(n6274), .ZN(n5072) );
  NOR3_X2 U4522 ( .A1(n6268), .A2(n8335), .A3(n6266), .ZN(n5071) );
  NAND3_X2 U4523 ( .A1(n7539), .A2(n7538), .A3(n5663), .ZN(n5075) );
  NAND3_X2 U4524 ( .A1(n7537), .A2(n7536), .A3(n6320), .ZN(n5058) );
  NOR2_X2 U4525 ( .A1(n8512), .A2(n8511), .ZN(n5080) );
  NAND3_X2 U4526 ( .A1(n5288), .A2(n7212), .A3(n4099), .ZN(n5294) );
  OAI21_X2 U4527 ( .B1(n4191), .B2(n5355), .A(n5365), .ZN(n5366) );
  OAI21_X2 U4528 ( .B1(n4159), .B2(n5305), .A(n5311), .ZN(n5313) );
  OAI21_X2 U4529 ( .B1(n6846), .B2(n6845), .A(n6844), .ZN(n6850) );
  OAI21_X2 U4530 ( .B1(n4125), .B2(n6842), .A(n6851), .ZN(n6852) );
  OAI21_X2 U4531 ( .B1(n6532), .B2(n6531), .A(n6394), .ZN(n6395) );
  OAI21_X2 U4532 ( .B1(n4281), .B2(n6416), .A(n6417), .ZN(n6540) );
  OAI21_X2 U4533 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5500) );
  OAI21_X2 U4534 ( .B1(n4247), .B2(n5537), .A(n5538), .ZN(n5583) );
  OAI21_X2 U4535 ( .B1(n4246), .B2(n5715), .A(n5724), .ZN(n5725) );
  OAI21_X2 U4536 ( .B1(n5673), .B2(n5672), .A(n5671), .ZN(n5674) );
  OAI21_X2 U4537 ( .B1(n4118), .B2(n5579), .A(n5600), .ZN(n5601) );
  OAI21_X2 U4538 ( .B1(n4282), .B2(n6442), .A(n6443), .ZN(n6549) );
  NAND3_X2 U4539 ( .A1(n5391), .A2(n7212), .A3(n4108), .ZN(n5393) );
  OAI21_X2 U4540 ( .B1(n7037), .B2(n4311), .A(n7252), .ZN(n7253) );
  OAI21_X2 U4541 ( .B1(n7028), .B2(n7027), .A(n7026), .ZN(n7029) );
  OAI21_X2 U4542 ( .B1(n6163), .B2(n6245), .A(n6162), .ZN(n8305) );
  NOR2_X2 U4543 ( .A1(n8306), .A2(n4753), .ZN(n6073) );
  NOR2_X2 U4544 ( .A1(n7528), .A2(n4752), .ZN(n6074) );
  OAI21_X2 U4545 ( .B1(n6249), .B2(n7034), .A(n6248), .ZN(n7245) );
  OAI21_X2 U4546 ( .B1(n7251), .B2(n7250), .A(n7249), .ZN(n7333) );
  OAI21_X2 U4547 ( .B1(n4286), .B2(n7040), .A(n7263), .ZN(n7264) );
  OAI21_X2 U4548 ( .B1(n7019), .B2(n7018), .A(n7017), .ZN(n7020) );
  OAI21_X2 U4549 ( .B1(n4262), .B2(n6393), .A(n6394), .ZN(n6531) );
  NOR3_X2 U4550 ( .A1(n6275), .A2(n6273), .A3(n6267), .ZN(n5081) );
  NOR3_X2 U4551 ( .A1(n5058), .A2(n6322), .A3(n5767), .ZN(n5079) );
  NOR3_X2 U4552 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(n5078) );
  OAI21_X2 U4553 ( .B1(n4160), .B2(n5327), .A(n5328), .ZN(n5356) );
  OAI21_X2 U4554 ( .B1(n6550), .B2(n6549), .A(n6443), .ZN(n6559) );
  NOR2_X2 U4555 ( .A1(n4837), .A2(n9021), .ZN(n5036) );
  NOR2_X2 U4556 ( .A1(n4837), .A2(n9040), .ZN(n5042) );
  NOR2_X2 U4557 ( .A1(n4837), .A2(n9019), .ZN(n5261) );
  NOR2_X2 U4558 ( .A1(n9035), .A2(n4836), .ZN(n5273) );
  NOR2_X2 U4559 ( .A1(n9003), .A2(n4837), .ZN(n5051) );
  NOR2_X2 U4560 ( .A1(n8960), .A2(n9054), .ZN(n5050) );
  OAI21_X2 U4561 ( .B1(n4254), .B2(n5433), .A(n5497), .ZN(n5498) );
  NOR2_X2 U4562 ( .A1(n9017), .A2(n4836), .ZN(n5269) );
  NOR2_X2 U4563 ( .A1(n9005), .A2(n4837), .ZN(n5046) );
  NOR2_X2 U4564 ( .A1(n8822), .A2(n9054), .ZN(n5045) );
  NOR2_X2 U4565 ( .A1(n4837), .A2(n9027), .ZN(n5246) );
  OAI21_X2 U4566 ( .B1(n4296), .B2(n6524), .A(n6724), .ZN(n6725) );
  OAI21_X2 U4567 ( .B1(n6492), .B2(n6566), .A(n6491), .ZN(n6493) );
  NOR2_X2 U4568 ( .A1(n4837), .A2(n9025), .ZN(n5039) );
  NOR2_X2 U4569 ( .A1(n9023), .A2(n4836), .ZN(n5060) );
  OAI21_X2 U4570 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6904) );
  OAI21_X2 U4571 ( .B1(n4300), .B2(n6745), .A(n6746), .ZN(n6903) );
  OAI21_X2 U4572 ( .B1(n5986), .B2(n5985), .A(n5984), .ZN(n5987) );
  OAI21_X2 U4573 ( .B1(n4215), .B2(n6027), .A(n6287), .ZN(n6288) );
  NOR2_X2 U4574 ( .A1(n9010), .A2(n4837), .ZN(n4996) );
  NOR2_X2 U4575 ( .A1(n8830), .A2(n4838), .ZN(n4995) );
  OAI21_X2 U4576 ( .B1(n4259), .B2(n5764), .A(n5984), .ZN(n5985) );
  OAI21_X2 U4577 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n7056) );
  OAI21_X2 U4578 ( .B1(n4270), .B2(n5640), .A(n5671), .ZN(n5672) );
  NOR2_X2 U4579 ( .A1(n9038), .A2(n4836), .ZN(n5064) );
  NOR2_X2 U4580 ( .A1(n4837), .A2(n9029), .ZN(n5236) );
  OAI21_X2 U4581 ( .B1(n7254), .B2(n7253), .A(n7252), .ZN(n7350) );
  NOR2_X2 U4582 ( .A1(n6159), .A2(n6073), .ZN(n6077) );
  AOI21_X2 U4583 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n7331) );
  NOR2_X2 U4584 ( .A1(n4771), .A2(n7527), .ZN(n7325) );
  OAI21_X2 U4585 ( .B1(n7329), .B2(n7328), .A(n7327), .ZN(n7330) );
  NOR2_X2 U4586 ( .A1(n4771), .A2(n7500), .ZN(n8315) );
  OAI21_X2 U4587 ( .B1(n7246), .B2(n7245), .A(n8313), .ZN(n7337) );
  OAI21_X2 U4588 ( .B1(n7265), .B2(n7264), .A(n7263), .ZN(n7342) );
  OAI21_X2 U4589 ( .B1(n4229), .B2(n6317), .A(n6361), .ZN(n6362) );
  NAND2_X2 U4590 ( .A1(n5082), .A2(n7546), .ZN(n8494) );
  INV_X4 U4591 ( .A(n8493), .ZN(n7531) );
  INV_X4 U4592 ( .A(n8494), .ZN(n7532) );
  INV_X4 U4593 ( .A(n8492), .ZN(n7530) );
  NOR2_X2 U4594 ( .A1(n8990), .A2(n4836), .ZN(n5106) );
  NOR2_X2 U4595 ( .A1(n8818), .A2(n9054), .ZN(n5105) );
  NOR2_X2 U4596 ( .A1(n9032), .A2(n4836), .ZN(n5228) );
  NOR2_X2 U4597 ( .A1(n8485), .A2(n7423), .ZN(n7384) );
  NOR2_X2 U4598 ( .A1(n9056), .A2(n4836), .ZN(n5149) );
  NOR2_X2 U4599 ( .A1(n8839), .A2(n4838), .ZN(n5148) );
  NOR2_X2 U4600 ( .A1(n8994), .A2(n4836), .ZN(n5134) );
  NOR2_X2 U4601 ( .A1(n8819), .A2(n4838), .ZN(n5133) );
  NOR2_X2 U4602 ( .A1(n8997), .A2(n4837), .ZN(n4982) );
  NOR2_X2 U4603 ( .A1(n8820), .A2(n9054), .ZN(n4981) );
  NOR2_X2 U4604 ( .A1(n8992), .A2(n4836), .ZN(n5101) );
  NOR2_X2 U4605 ( .A1(n8840), .A2(n4838), .ZN(n5100) );
  NAND3_X2 U4606 ( .A1(n4967), .A2(n4966), .A3(n4965), .ZN(n7988) );
  NAND3_X2 U4607 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n7977) );
  NOR2_X2 U4608 ( .A1(n4973), .A2(n4972), .ZN(n4974) );
  AOI21_X2 U4609 ( .B1(n4468), .B2(n8364), .A(n7532), .ZN(n5178) );
  OAI21_X2 U4610 ( .B1(n4302), .B2(n6880), .A(n6992), .ZN(n6993) );
  OAI22_X2 U4611 ( .A1(n7496), .A2(n8624), .B1(n8590), .B2(n8591), .ZN(n8564)
         );
  OAI22_X2 U4612 ( .A1(n7500), .A2(n8614), .B1(n8615), .B2(n8589), .ZN(n8552)
         );
  OAI22_X2 U4613 ( .A1(n7512), .A2(n8637), .B1(n8638), .B2(n8597), .ZN(n8544)
         );
  OAI22_X2 U4614 ( .A1(n7504), .A2(n8609), .B1(n8539), .B2(n8540), .ZN(n8555)
         );
  NOR2_X2 U4615 ( .A1(n8371), .A2(n4128), .ZN(n5652) );
  OAI22_X2 U4616 ( .A1(n7499), .A2(n8618), .B1(n8619), .B2(n8587), .ZN(n8570)
         );
  OAI22_X2 U4617 ( .A1(n7497), .A2(n8621), .B1(n8576), .B2(n8577), .ZN(n8567)
         );
  OAI21_X2 U4618 ( .B1(n4152), .B2(n8605), .A(n5926), .ZN(n6329) );
  NAND3_X2 U4619 ( .A1(n4455), .A2(n4784), .A3(n5592), .ZN(n5594) );
  OAI21_X2 U4620 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(n8542) );
  NOR2_X2 U4621 ( .A1(n9015), .A2(n4836), .ZN(n5200) );
  OAI21_X2 U4622 ( .B1(n4304), .B2(n7042), .A(n7268), .ZN(n7269) );
  OAI21_X2 U4623 ( .B1(n7270), .B2(n7269), .A(n7268), .ZN(n7271) );
  NAND3_X2 U4624 ( .A1(n8499), .A2(n6253), .A3(n6252), .ZN(n6255) );
  NOR2_X2 U4625 ( .A1(n9046), .A2(n4837), .ZN(n5003) );
  AOI21_X2 U4626 ( .B1(n4737), .B2(n7523), .A(n7532), .ZN(n5443) );
  NAND3_X2 U4627 ( .A1(n5091), .A2(n8494), .A3(n5090), .ZN(n8452) );
  NOR2_X2 U4628 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  NOR2_X2 U4629 ( .A1(n8966), .A2(n4838), .ZN(n5067) );
  NAND2_X2 U4630 ( .A1(n8541), .A2(n8542), .ZN(n8543) );
  AOI21_X2 U4631 ( .B1(n7243), .B2(n6936), .A(n6935), .ZN(n6937) );
  NOR2_X2 U4632 ( .A1(n7241), .A2(n6934), .ZN(n6935) );
  NOR2_X2 U4633 ( .A1(n5946), .A2(n4128), .ZN(n5947) );
  NOR2_X2 U4634 ( .A1(n5945), .A2(n7393), .ZN(n5948) );
  AOI211_X2 U4635 ( .C1(n7525), .C2(n5140), .A(n8405), .B(n8392), .ZN(n5944)
         );
  INV_X4 U4636 ( .A(n8476), .ZN(n7558) );
  NAND3_X2 U4637 ( .A1(n5123), .A2(n8494), .A3(n5122), .ZN(n8472) );
  NAND3_X2 U4638 ( .A1(n5128), .A2(n8494), .A3(n5127), .ZN(n8473) );
  NOR2_X2 U4639 ( .A1(n7918), .A2(n7525), .ZN(n8391) );
  NOR2_X2 U4640 ( .A1(n9001), .A2(n4837), .ZN(n4991) );
  NOR2_X2 U4641 ( .A1(n8821), .A2(n4838), .ZN(n4990) );
  INV_X4 U4642 ( .A(n4079), .ZN(n4836) );
  AOI21_X2 U4643 ( .B1(n7273), .B2(n6894), .A(n6893), .ZN(n6895) );
  NOR2_X2 U4644 ( .A1(n6892), .A2(n7362), .ZN(n6893) );
  NAND3_X2 U4645 ( .A1(n5099), .A2(n8494), .A3(n5098), .ZN(n8381) );
  NOR2_X2 U4646 ( .A1(n8333), .A2(n7558), .ZN(n8380) );
  NOR2_X2 U4647 ( .A1(n5464), .A2(n4736), .ZN(n5465) );
  NOR2_X2 U4648 ( .A1(n5944), .A2(n7393), .ZN(n5449) );
  NOR2_X2 U4649 ( .A1(n5946), .A2(n4734), .ZN(n5450) );
  NOR2_X2 U4650 ( .A1(n5644), .A2(n4128), .ZN(n5447) );
  AOI21_X2 U4651 ( .B1(n7387), .B2(n7560), .A(n7386), .ZN(n7388) );
  NOR2_X2 U4652 ( .A1(n8486), .A2(n7547), .ZN(n7386) );
  NOR2_X2 U4653 ( .A1(n8318), .A2(n8317), .ZN(n8515) );
  OAI21_X2 U4654 ( .B1(n8154), .B2(n8155), .A(n6072), .ZN(n5882) );
  OAI21_X2 U4655 ( .B1(n4805), .B2(n7663), .A(n4804), .ZN(n6039) );
  NOR2_X2 U4656 ( .A1(n7488), .A2(n7216), .ZN(n5954) );
  OAI21_X2 U4657 ( .B1(n4805), .B2(n7659), .A(n4804), .ZN(n5955) );
  OAI21_X2 U4658 ( .B1(n4805), .B2(n7665), .A(n4804), .ZN(n5936) );
  NOR2_X2 U4659 ( .A1(n5829), .A2(n4563), .ZN(n5830) );
  NOR2_X2 U4660 ( .A1(n4734), .A2(n6263), .ZN(n5829) );
  OAI21_X2 U4661 ( .B1(n4805), .B2(n7661), .A(n4804), .ZN(n5831) );
  AOI21_X2 U4662 ( .B1(n7551), .B2(n4077), .A(n4082), .ZN(n5981) );
  NOR2_X2 U4663 ( .A1(n4738), .A2(n5974), .ZN(n5980) );
  NAND3_X2 U4664 ( .A1(n5221), .A2(n4386), .A3(n5220), .ZN(n7657) );
  AOI21_X2 U4665 ( .B1(n5962), .B2(n7977), .A(n5961), .ZN(n5966) );
  OAI21_X2 U4666 ( .B1(n4805), .B2(n7657), .A(n4804), .ZN(n5962) );
  NOR2_X2 U4667 ( .A1(n8361), .A2(n7216), .ZN(n5961) );
  OAI22_X2 U4668 ( .A1(n7502), .A2(n8611), .B1(n8612), .B2(n8583), .ZN(n8584)
         );
  NOR2_X2 U4669 ( .A1(n5944), .A2(n4128), .ZN(n5820) );
  NOR2_X2 U4670 ( .A1(n5945), .A2(n4734), .ZN(n5821) );
  NAND3_X2 U4671 ( .A1(n5780), .A2(n4431), .A3(n5779), .ZN(n7722) );
  OAI21_X2 U4672 ( .B1(n4082), .B2(n5454), .A(n6322), .ZN(n5457) );
  OAI21_X2 U4673 ( .B1(n4805), .B2(n6322), .A(n4804), .ZN(n5455) );
  NOR2_X2 U4674 ( .A1(n7912), .A2(n4738), .ZN(n5453) );
  OAI21_X2 U4675 ( .B1(n8380), .B2(n8473), .A(n8382), .ZN(n6263) );
  NOR2_X2 U4676 ( .A1(n9044), .A2(n4837), .ZN(n4956) );
  AOI21_X2 U4677 ( .B1(n7553), .B2(n4077), .A(n4082), .ZN(n5813) );
  NOR2_X2 U4678 ( .A1(n8427), .A2(n7216), .ZN(n5811) );
  NOR2_X2 U4679 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  NOR2_X2 U4680 ( .A1(n5651), .A2(n4734), .ZN(n5653) );
  NOR2_X2 U4681 ( .A1(n8379), .A2(n4128), .ZN(n5647) );
  NOR2_X2 U4682 ( .A1(n6277), .A2(n4734), .ZN(n5648) );
  OAI21_X2 U4683 ( .B1(n4082), .B2(n5187), .A(n5267), .ZN(n5190) );
  OAI21_X2 U4684 ( .B1(n4805), .B2(n5267), .A(n4804), .ZN(n5188) );
  OAI21_X2 U4685 ( .B1(n5593), .B2(n5592), .A(n5594), .ZN(n7889) );
  NOR2_X2 U4686 ( .A1(n7571), .A2(n4078), .ZN(n5593) );
  OAI21_X2 U4687 ( .B1(n4088), .B2(n6324), .A(n8545), .ZN(n8594) );
  NOR2_X2 U4688 ( .A1(n8379), .A2(n7393), .ZN(n5112) );
  NOR2_X2 U4689 ( .A1(n8402), .A2(n4128), .ZN(n5113) );
  NOR2_X2 U4690 ( .A1(n8362), .A2(n4734), .ZN(n5110) );
  NOR2_X2 U4691 ( .A1(n8416), .A2(n4128), .ZN(n5144) );
  NOR2_X2 U4692 ( .A1(n5644), .A2(n4734), .ZN(n5139) );
  NOR2_X2 U4693 ( .A1(n8379), .A2(n4734), .ZN(n5485) );
  NOR2_X2 U4694 ( .A1(n6277), .A2(n4736), .ZN(n5486) );
  NOR3_X2 U4695 ( .A1(n5159), .A2(n5158), .A3(n5157), .ZN(n7526) );
  NOR2_X2 U4696 ( .A1(n5651), .A2(n7393), .ZN(n5158) );
  NOR2_X2 U4697 ( .A1(n8444), .A2(n4317), .ZN(n5157) );
  NOR2_X2 U4698 ( .A1(n7429), .A2(n7216), .ZN(n7217) );
  OAI21_X2 U4699 ( .B1(n4082), .B2(n7210), .A(n7211), .ZN(n7215) );
  OAI21_X2 U4700 ( .B1(n7211), .B2(n4805), .A(n4804), .ZN(n7213) );
  NOR2_X2 U4701 ( .A1(n7207), .A2(n4738), .ZN(n7208) );
  AOI21_X2 U4702 ( .B1(n7423), .B2(n5586), .A(n6159), .ZN(n5589) );
  NOR2_X2 U4703 ( .A1(n8401), .A2(n7216), .ZN(n5153) );
  OAI21_X2 U4704 ( .B1(n4805), .B2(n7648), .A(n4804), .ZN(n5154) );
  AOI21_X2 U4705 ( .B1(n7641), .B2(n8629), .A(n8630), .ZN(n8580) );
  NOR2_X2 U4706 ( .A1(n8444), .A2(n4128), .ZN(n5802) );
  NOR2_X2 U4707 ( .A1(n8428), .A2(n4734), .ZN(n6278) );
  NOR2_X2 U4708 ( .A1(n9014), .A2(n4837), .ZN(n5011) );
  NOR2_X2 U4709 ( .A1(n8837), .A2(n4838), .ZN(n5010) );
  OAI21_X2 U4710 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(n6285) );
  OAI21_X2 U4711 ( .B1(n4162), .B2(n6319), .A(n6530), .ZN(n8464) );
  OAI21_X2 U4712 ( .B1(n6256), .B2(n6255), .A(n6254), .ZN(n6261) );
  NAND3_X2 U4713 ( .A1(n5094), .A2(n5093), .A3(n5092), .ZN(n8306) );
  NOR2_X2 U4714 ( .A1(n4505), .A2(n5446), .ZN(n5945) );
  OAI21_X2 U4715 ( .B1(n8378), .B2(n7563), .A(n5445), .ZN(n5446) );
  NOR2_X2 U4716 ( .A1(n5656), .A2(n4738), .ZN(n5657) );
  NOR2_X2 U4717 ( .A1(n5976), .A2(n5978), .ZN(n5658) );
  NOR2_X2 U4718 ( .A1(n7505), .A2(n7216), .ZN(n5659) );
  OAI21_X2 U4719 ( .B1(n7909), .B2(n5720), .A(n5719), .ZN(n5721) );
  OAI21_X2 U4720 ( .B1(n4268), .B2(n5766), .A(n6030), .ZN(n7702) );
  OAI21_X2 U4721 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n7287) );
  OAI21_X2 U4722 ( .B1(n7549), .B2(n8636), .A(n8543), .ZN(n8602) );
  NOR2_X2 U4723 ( .A1(n8427), .A2(n4738), .ZN(n5490) );
  NOR2_X2 U4724 ( .A1(n5488), .A2(n5978), .ZN(n5489) );
  NOR2_X2 U4725 ( .A1(n7526), .A2(n7216), .ZN(n5491) );
  INV_X4 U4726 ( .A(n5975), .ZN(n7219) );
  OAI21_X2 U4727 ( .B1(n7710), .B2(n7711), .A(n5596), .ZN(n5597) );
  OAI21_X2 U4728 ( .B1(n4267), .B2(n5642), .A(n5718), .ZN(n7689) );
  NOR2_X2 U4729 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND3_X2 U4730 ( .A1(n5778), .A2(n5777), .A3(n5776), .ZN(n7721) );
  NOR2_X2 U4731 ( .A1(n8371), .A2(n7393), .ZN(n5165) );
  NOR2_X2 U4732 ( .A1(n8341), .A2(n4128), .ZN(n5166) );
  AOI21_X2 U4733 ( .B1(n8472), .B2(n7558), .A(n7564), .ZN(n5156) );
  NAND3_X2 U4734 ( .A1(n5119), .A2(n4430), .A3(n5118), .ZN(n8326) );
  NOR2_X2 U4735 ( .A1(n8370), .A2(n7216), .ZN(n5469) );
  OAI21_X2 U4736 ( .B1(n4805), .B2(n7617), .A(n4804), .ZN(n5470) );
  NOR2_X2 U4737 ( .A1(n8987), .A2(n4836), .ZN(n5240) );
  NAND3_X2 U4738 ( .A1(n7367), .A2(n7366), .A3(n7365), .ZN(n7368) );
  OAI21_X2 U4739 ( .B1(n6918), .B2(n7312), .A(n6917), .ZN(n7409) );
  OAI21_X2 U4740 ( .B1(n8380), .B2(n8381), .A(n8382), .ZN(n5941) );
  NAND2_X2 U4741 ( .A1(n6040), .A2(n4091), .ZN(n8324) );
  NAND2_X2 U4742 ( .A1(n7209), .A2(n4091), .ZN(n8323) );
  NOR2_X2 U4743 ( .A1(n5448), .A2(n5447), .ZN(n5452) );
  NOR2_X2 U4744 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NOR2_X2 U4745 ( .A1(n5945), .A2(n4317), .ZN(n5448) );
  NAND3_X2 U4746 ( .A1(n5782), .A2(n4432), .A3(n5781), .ZN(n7723) );
  AOI21_X2 U4747 ( .B1(n7424), .B2(n4804), .A(n7423), .ZN(n7425) );
  OAI21_X2 U4748 ( .B1(n7429), .B2(n4738), .A(n7428), .ZN(n7433) );
  NOR2_X2 U4749 ( .A1(n8477), .A2(n4469), .ZN(n7431) );
  NOR2_X2 U4750 ( .A1(n4804), .A2(n7430), .ZN(n7432) );
  NOR2_X2 U4751 ( .A1(n7609), .A2(n4742), .ZN(n4935) );
  NOR2_X2 U4752 ( .A1(n7608), .A2(n4742), .ZN(n4944) );
  NOR2_X2 U4753 ( .A1(n7580), .A2(n4742), .ZN(n4940) );
  NOR2_X2 U4754 ( .A1(n7582), .A2(n4742), .ZN(n5169) );
  NOR2_X2 U4755 ( .A1(n7579), .A2(n4742), .ZN(n4977) );
  NOR2_X2 U4756 ( .A1(n7578), .A2(n4742), .ZN(n4968) );
  NOR2_X2 U4757 ( .A1(n7607), .A2(n4742), .ZN(n4986) );
  INV_X4 U4758 ( .A(n4803), .ZN(n4800) );
  AOI21_X2 U4759 ( .B1(n7613), .B2(n4744), .A(n6072), .ZN(n5884) );
  INV_X4 U4760 ( .A(n4803), .ZN(n4799) );
  INV_X4 U4761 ( .A(n4803), .ZN(n4798) );
  NOR2_X2 U4762 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  OAI21_X2 U4763 ( .B1(iAddr[13]), .B2(n6063), .A(n6064), .ZN(n8082) );
  OAI21_X2 U4764 ( .B1(iAddr[11]), .B2(n6060), .A(n6061), .ZN(n8070) );
  OAI21_X2 U4765 ( .B1(iAddr[9]), .B2(n6057), .A(n6058), .ZN(n8058) );
  OAI21_X2 U4766 ( .B1(iAddr[7]), .B2(n6054), .A(n6055), .ZN(n8046) );
  OAI21_X2 U4767 ( .B1(iAddr[5]), .B2(n6051), .A(n6052), .ZN(n8034) );
  OAI21_X2 U4768 ( .B1(iAddr[4]), .B2(n6050), .A(n6049), .ZN(n8029) );
  OAI21_X2 U4769 ( .B1(iAddr[2]), .B2(iAddr[3]), .A(n6048), .ZN(n8025) );
  NOR2_X2 U4770 ( .A1(n7442), .A2(n6046), .ZN(n6047) );
  OAI21_X2 U4771 ( .B1(iAddr[22]), .B2(n6038), .A(n6037), .ZN(n8010) );
  OAI21_X2 U4772 ( .B1(iAddr[17]), .B2(n6034), .A(n6035), .ZN(n8003) );
  INV_X4 U4773 ( .A(n4779), .ZN(n4777) );
  OAI21_X2 U4774 ( .B1(iAddr[15]), .B2(n6031), .A(n6032), .ZN(n7994) );
  NOR2_X2 U4775 ( .A1(n7447), .A2(n6046), .ZN(n5972) );
  AOI21_X2 U4776 ( .B1(n5955), .B2(n7968), .A(n5954), .ZN(n5959) );
  NAND3_X2 U4777 ( .A1(n5938), .A2(n4287), .A3(n5937), .ZN(n7458) );
  AOI222_X1 U4778 ( .A1(n7209), .A2(n7295), .B1(n7960), .B2(n7665), .C1(n6040), 
        .C2(n7962), .ZN(n5938) );
  NOR2_X2 U4779 ( .A1(n7456), .A2(n6046), .ZN(n5940) );
  OAI21_X2 U4780 ( .B1(iAddr[29]), .B2(n5922), .A(n6067), .ZN(n7952) );
  OAI21_X2 U4781 ( .B1(iAddr[28]), .B2(n5918), .A(n5921), .ZN(n7949) );
  OAI21_X2 U4782 ( .B1(iAddr[27]), .B2(n5914), .A(n5917), .ZN(n7946) );
  OAI21_X2 U4783 ( .B1(iAddr[26]), .B2(n5910), .A(n5913), .ZN(n7943) );
  OAI21_X2 U4784 ( .B1(iAddr[25]), .B2(n5906), .A(n5909), .ZN(n7940) );
  OAI21_X2 U4785 ( .B1(iAddr[24]), .B2(n5902), .A(n5905), .ZN(n7937) );
  OAI21_X2 U4786 ( .B1(iAddr[23]), .B2(n5898), .A(n5901), .ZN(n7934) );
  OAI21_X2 U4787 ( .B1(iAddr[21]), .B2(n5892), .A(n5897), .ZN(n7931) );
  OAI21_X2 U4788 ( .B1(iAddr[20]), .B2(n5888), .A(n5891), .ZN(n7928) );
  OAI21_X2 U4789 ( .B1(iAddr[19]), .B2(n5881), .A(n5887), .ZN(n7924) );
  NOR2_X2 U4790 ( .A1(n7462), .A2(n6046), .ZN(n5837) );
  INV_X4 U4791 ( .A(n4779), .ZN(n4776) );
  INV_X4 U4792 ( .A(n4780), .ZN(n4775) );
  NOR2_X2 U4793 ( .A1(n8806), .A2(n4772), .ZN(n7145) );
  NOR2_X2 U4794 ( .A1(n8808), .A2(n4772), .ZN(n7151) );
  NOR2_X2 U4795 ( .A1(n8809), .A2(n4772), .ZN(n7155) );
  NOR2_X2 U4796 ( .A1(n8810), .A2(n4772), .ZN(n7159) );
  NOR2_X2 U4797 ( .A1(n8811), .A2(n4772), .ZN(n7166) );
  INV_X4 U4798 ( .A(n4792), .ZN(n4789) );
  INV_X4 U4799 ( .A(rst), .ZN(n4887) );
  INV_X4 U4800 ( .A(rst), .ZN(n4892) );
  INV_X4 U4801 ( .A(n4821), .ZN(n4819) );
  NAND2_X2 U4802 ( .A1(n7805), .A2(n4824), .ZN(n7763) );
  AOI21_X2 U4803 ( .B1(n7750), .B2(n7740), .A(n4820), .ZN(n7747) );
  INV_X4 U4804 ( .A(rst), .ZN(n4881) );
  INV_X4 U4805 ( .A(n4823), .ZN(n4813) );
  INV_X4 U4806 ( .A(n4823), .ZN(n4814) );
  INV_X4 U4807 ( .A(n4823), .ZN(n4812) );
  INV_X4 U4808 ( .A(n4821), .ZN(n4817) );
  NOR2_X2 U4809 ( .A1(n7634), .A2(n7628), .ZN(n7194) );
  INV_X4 U4810 ( .A(n4781), .ZN(n4774) );
  INV_X4 U4811 ( .A(n5967), .ZN(n7507) );
  INV_X4 U4812 ( .A(n6046), .ZN(n7506) );
  AOI211_X2 U4813 ( .C1(n7427), .C2(n7700), .A(n5983), .B(n5982), .ZN(n7987)
         );
  NOR2_X2 U4814 ( .A1(n5980), .A2(n5979), .ZN(n7986) );
  NOR2_X2 U4815 ( .A1(n7541), .A2(n5981), .ZN(n5983) );
  OAI21_X2 U4816 ( .B1(n8533), .B2(n8534), .A(n8535), .ZN(n7664) );
  NAND3_X2 U4817 ( .A1(n5662), .A2(n4470), .A3(n5661), .ZN(n7695) );
  AOI21_X2 U4818 ( .B1(n6712), .B2(n4794), .A(n6711), .ZN(n6713) );
  AOI21_X2 U4819 ( .B1(n6710), .B2(n7896), .A(n7533), .ZN(n6711) );
  NOR2_X2 U4820 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND3_X2 U4821 ( .A1(n5775), .A2(n4477), .A3(n5774), .ZN(n7720) );
  AOI21_X2 U4822 ( .B1(n6945), .B2(n4794), .A(n6944), .ZN(n6946) );
  AOI21_X2 U4823 ( .B1(n6943), .B2(n7896), .A(n7535), .ZN(n6944) );
  AOI21_X2 U4824 ( .B1(n6956), .B2(n7896), .A(n7519), .ZN(n6957) );
  AOI21_X2 U4825 ( .B1(n6970), .B2(n7896), .A(n7517), .ZN(n6971) );
  NOR2_X2 U4826 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  NOR2_X2 U4827 ( .A1(n4128), .A2(n6263), .ZN(n5462) );
  NOR2_X2 U4828 ( .A1(n8341), .A2(n4734), .ZN(n5461) );
  NAND3_X2 U4829 ( .A1(n5773), .A2(n5772), .A3(n5771), .ZN(n8304) );
  OAI21_X2 U4830 ( .B1(n7894), .B2(n8304), .A(n7896), .ZN(n6991) );
  NAND3_X2 U4831 ( .A1(n5650), .A2(n4471), .A3(n5649), .ZN(n7700) );
  NOR2_X2 U4832 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  NAND3_X2 U4833 ( .A1(n5646), .A2(n4476), .A3(n5645), .ZN(n7699) );
  AOI21_X2 U4834 ( .B1(n7083), .B2(n4794), .A(n7082), .ZN(n7084) );
  AOI21_X2 U4835 ( .B1(n7081), .B2(n7896), .A(n7518), .ZN(n7082) );
  AOI21_X2 U4836 ( .B1(n7427), .B2(n7888), .A(n5191), .ZN(n5192) );
  AOI21_X2 U4837 ( .B1(n7101), .B2(n7896), .A(n7511), .ZN(n7102) );
  NOR2_X2 U4838 ( .A1(n5111), .A2(n5110), .ZN(n5115) );
  NOR2_X2 U4839 ( .A1(n5113), .A2(n5112), .ZN(n5114) );
  NOR2_X2 U4840 ( .A1(n6277), .A2(n4317), .ZN(n5111) );
  AOI21_X2 U4841 ( .B1(n4312), .B2(n5800), .A(n5144), .ZN(n5145) );
  NOR2_X2 U4842 ( .A1(n5139), .A2(n5138), .ZN(n5143) );
  NOR2_X2 U4843 ( .A1(n5946), .A2(n7393), .ZN(n5138) );
  AOI21_X2 U4844 ( .B1(n6577), .B2(n4794), .A(n6576), .ZN(n6578) );
  AOI21_X2 U4845 ( .B1(n6575), .B2(n7896), .A(n7534), .ZN(n6576) );
  AOI21_X2 U4846 ( .B1(n7200), .B2(n7896), .A(n7542), .ZN(n7201) );
  NAND3_X2 U4847 ( .A1(n4122), .A2(n4472), .A3(n5487), .ZN(n7685) );
  NOR2_X2 U4848 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  AOI21_X2 U4849 ( .B1(n5154), .B2(n5767), .A(n5153), .ZN(n5164) );
  NOR2_X2 U4850 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NOR2_X2 U4851 ( .A1(n8416), .A2(n7393), .ZN(n5801) );
  NOR2_X2 U4852 ( .A1(n6279), .A2(n6278), .ZN(n6281) );
  NOR2_X2 U4853 ( .A1(n6277), .A2(n4128), .ZN(n6279) );
  OAI21_X2 U4854 ( .B1(n7238), .B2(n7237), .A(n7236), .ZN(n7239) );
  OAI21_X2 U4855 ( .B1(n4587), .B2(n7277), .A(n7370), .ZN(n7371) );
  OAI21_X2 U4856 ( .B1(n7894), .B2(n8306), .A(n7896), .ZN(n7279) );
  INV_X4 U4857 ( .A(n7293), .ZN(n7492) );
  NOR3_X2 U4858 ( .A1(n5659), .A2(n5658), .A3(n5657), .ZN(n7693) );
  AOI21_X2 U4859 ( .B1(n5664), .B2(n4804), .A(n5663), .ZN(n5666) );
  OAI21_X2 U4860 ( .B1(n7294), .B2(n7293), .A(n7292), .ZN(n7296) );
  NAND3_X2 U4861 ( .A1(n5770), .A2(n5769), .A3(n5768), .ZN(n8316) );
  OAI21_X2 U4862 ( .B1(n4805), .B2(n7623), .A(n4804), .ZN(n5492) );
  AOI21_X2 U4863 ( .B1(n7304), .B2(n7896), .A(n7543), .ZN(n7305) );
  AOI21_X2 U4864 ( .B1(n5942), .B2(n4312), .A(n4563), .ZN(n5943) );
  AOI21_X2 U4865 ( .B1(n7314), .B2(n7896), .A(n7510), .ZN(n7315) );
  NAND3_X2 U4866 ( .A1(n4473), .A2(n5168), .A3(n5167), .ZN(n7888) );
  NOR2_X2 U4867 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  AOI21_X2 U4868 ( .B1(n5470), .B2(n7671), .A(n5469), .ZN(n5474) );
  INV_X4 U4869 ( .A(rst), .ZN(n4883) );
  AOI21_X2 U4870 ( .B1(n8323), .B2(n7674), .A(n8333), .ZN(n7380) );
  OAI21_X2 U4871 ( .B1(n7674), .B2(n7547), .A(n7896), .ZN(n7382) );
  INV_X4 U4872 ( .A(rst), .ZN(n4884) );
  AOI21_X2 U4873 ( .B1(n7413), .B2(n7896), .A(n7522), .ZN(n7414) );
  NOR2_X2 U4874 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  NOR2_X2 U4875 ( .A1(n4128), .A2(n5941), .ZN(n5441) );
  NOR2_X2 U4876 ( .A1(n8402), .A2(n4734), .ZN(n5440) );
  INV_X4 U4877 ( .A(rst), .ZN(n4882) );
  NAND3_X2 U4878 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(regWrData[3]) );
  AOI21_X2 U4879 ( .B1(reg31Val_0[3]), .B2(n4741), .A(n5129), .ZN(n5132) );
  NOR2_X2 U4880 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  NOR2_X2 U4881 ( .A1(n5210), .A2(n4391), .ZN(n5025) );
  NOR2_X2 U4882 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  NOR2_X2 U4883 ( .A1(n5210), .A2(n4390), .ZN(n5021) );
  NOR2_X2 U4884 ( .A1(n5007), .A2(n5006), .ZN(n5008) );
  NOR2_X2 U4885 ( .A1(n5210), .A2(n4441), .ZN(n5006) );
  NAND3_X2 U4886 ( .A1(n5198), .A2(n5197), .A3(n4376), .ZN(regWrData[16]) );
  NAND3_X2 U4887 ( .A1(n5208), .A2(n5207), .A3(n4379), .ZN(regWrData[17]) );
  NAND3_X2 U4888 ( .A1(n5206), .A2(n5205), .A3(n4378), .ZN(regWrData[18]) );
  NAND3_X2 U4889 ( .A1(n5035), .A2(n5034), .A3(n4425), .ZN(regWrData[19]) );
  NAND3_X2 U4890 ( .A1(n4964), .A2(n4963), .A3(n4423), .ZN(regWrData[20]) );
  NAND3_X2 U4891 ( .A1(n5033), .A2(n5032), .A3(n4424), .ZN(regWrData[21]) );
  NAND3_X2 U4892 ( .A1(n5085), .A2(n5084), .A3(n4426), .ZN(regWrData[22]) );
  NAND3_X2 U4893 ( .A1(n5117), .A2(n5116), .A3(n4427), .ZN(regWrData[23]) );
  NAND3_X2 U4894 ( .A1(n5196), .A2(n5195), .A3(n4377), .ZN(regWrData[24]) );
  NAND3_X2 U4895 ( .A1(n5213), .A2(n5212), .A3(n4380), .ZN(regWrData[25]) );
  NAND3_X2 U4896 ( .A1(n5031), .A2(n5030), .A3(n4422), .ZN(regWrData[27]) );
  NAND3_X2 U4897 ( .A1(n4954), .A2(n4953), .A3(n4419), .ZN(regWrData[29]) );
  OAI21_X2 U4898 ( .B1(n8902), .B2(n7123), .A(n7122), .ZN(iAddr[0]) );
  OAI21_X2 U4899 ( .B1(n8871), .B2(n7123), .A(n7113), .ZN(iAddr[1]) );
  OAI21_X2 U4900 ( .B1(n4360), .B2(n7127), .A(n7126), .ZN(n3669) );
  NAND3_X2 U4901 ( .A1(regWr), .A2(n7853), .A3(n4558), .ZN(n7126) );
  INV_X4 U4902 ( .A(n4892), .ZN(n4878) );
  NOR3_X2 U4903 ( .A1(n8125), .A2(n8126), .A3(n8127), .ZN(n6070) );
  NOR2_X2 U4904 ( .A1(n5973), .A2(n5972), .ZN(n7975) );
  NOR2_X2 U4905 ( .A1(n7658), .A2(n7982), .ZN(n5960) );
  OAI21_X2 U4906 ( .B1(n8723), .B2(n4810), .A(n6695), .ZN(n3523) );
  NOR2_X2 U4907 ( .A1(n7982), .A2(n7664), .ZN(n5939) );
  NOR2_X2 U4908 ( .A1(n7660), .A2(n7982), .ZN(n5836) );
  OAI21_X2 U4909 ( .B1(n9045), .B2(n4772), .A(n7070), .ZN(n9167) );
  OAI21_X2 U4910 ( .B1(n8760), .B2(n4810), .A(n7114), .ZN(n3611) );
  INV_X4 U4911 ( .A(n4881), .ZN(n4844) );
  OAI21_X2 U4912 ( .B1(n8789), .B2(n4810), .A(n7124), .ZN(n3665) );
  INV_X4 U4913 ( .A(n4880), .ZN(n4842) );
  INV_X4 U4914 ( .A(n4881), .ZN(n4843) );
  NOR2_X2 U4915 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NOR2_X2 U4916 ( .A1(n9029), .A2(n7164), .ZN(n7144) );
  NOR2_X2 U4917 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NOR2_X2 U4918 ( .A1(n9038), .A2(n7164), .ZN(n7150) );
  INV_X4 U4919 ( .A(n4886), .ZN(n4861) );
  NOR2_X2 U4920 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  NOR2_X2 U4921 ( .A1(n9042), .A2(n7164), .ZN(n7154) );
  NOR2_X2 U4922 ( .A1(n7159), .A2(n7158), .ZN(n7160) );
  NOR2_X2 U4923 ( .A1(n9046), .A2(n7164), .ZN(n7158) );
  NOR2_X2 U4924 ( .A1(n7166), .A2(n7165), .ZN(n7167) );
  NOR2_X2 U4925 ( .A1(n8987), .A2(n7164), .ZN(n7165) );
  INV_X4 U4926 ( .A(n4890), .ZN(n4872) );
  INV_X4 U4927 ( .A(n4887), .ZN(n4863) );
  INV_X4 U4928 ( .A(n4891), .ZN(n4874) );
  INV_X4 U4929 ( .A(n4887), .ZN(n4864) );
  INV_X4 U4930 ( .A(n4890), .ZN(n4871) );
  OAI21_X2 U4931 ( .B1(n4772), .B2(n4651), .A(n7169), .ZN(n9177) );
  INV_X4 U4932 ( .A(n4886), .ZN(n4860) );
  INV_X4 U4933 ( .A(n4887), .ZN(n4862) );
  OAI21_X2 U4934 ( .B1(n8817), .B2(n4772), .A(n7191), .ZN(n3763) );
  INV_X4 U4935 ( .A(n4892), .ZN(n4877) );
  INV_X4 U4936 ( .A(n4891), .ZN(n4875) );
  INV_X4 U4937 ( .A(n4881), .ZN(n4845) );
  INV_X4 U4938 ( .A(n4888), .ZN(n4856) );
  INV_X4 U4939 ( .A(n4890), .ZN(n4873) );
  INV_X4 U4940 ( .A(n4891), .ZN(n4876) );
  INV_X4 U4941 ( .A(n4880), .ZN(n4841) );
  INV_X4 U4942 ( .A(n4889), .ZN(n4869) );
  INV_X4 U4943 ( .A(n4889), .ZN(n4868) );
  INV_X4 U4944 ( .A(n4882), .ZN(n4847) );
  INV_X4 U4945 ( .A(n4882), .ZN(n4848) );
  NOR2_X2 U4946 ( .A1(n7726), .A2(n7641), .ZN(n7193) );
  NAND3_X2 U4947 ( .A1(n7225), .A2(n7224), .A3(n7223), .ZN(n3965) );
  NOR2_X2 U4948 ( .A1(n5480), .A2(n5479), .ZN(n7668) );
  NAND3_X2 U4949 ( .A1(n7440), .A2(n7439), .A3(n7438), .ZN(n3978) );
  NOR2_X2 U4950 ( .A1(n7444), .A2(n7443), .ZN(n7446) );
  NOR2_X2 U4951 ( .A1(n7615), .A2(n7442), .ZN(n7443) );
  NOR2_X2 U4952 ( .A1(n4502), .A2(n6953), .ZN(n6960) );
  AOI21_X2 U4953 ( .B1(n6958), .B2(n4794), .A(n6957), .ZN(n6959) );
  NOR2_X2 U4954 ( .A1(n4496), .A2(n6967), .ZN(n6974) );
  AOI21_X2 U4955 ( .B1(n6972), .B2(n4794), .A(n6971), .ZN(n6973) );
  NOR2_X2 U4956 ( .A1(n4503), .A2(n7098), .ZN(n7105) );
  AOI21_X2 U4957 ( .B1(n7103), .B2(n4794), .A(n7102), .ZN(n7104) );
  NOR2_X2 U4958 ( .A1(n4478), .A2(n7197), .ZN(n7204) );
  AOI21_X2 U4959 ( .B1(n7202), .B2(n4794), .A(n7201), .ZN(n7203) );
  AOI211_X2 U4960 ( .C1(n7230), .C2(n4794), .A(n7229), .B(n7228), .ZN(n7231)
         );
  INV_X4 U4961 ( .A(n4883), .ZN(n4851) );
  INV_X4 U4962 ( .A(n4884), .ZN(n4853) );
  NOR3_X2 U4963 ( .A1(n7296), .A2(n4494), .A3(n4295), .ZN(n7297) );
  INV_X4 U4964 ( .A(n4883), .ZN(n4850) );
  NOR2_X2 U4965 ( .A1(n4495), .A2(n7301), .ZN(n7308) );
  NOR2_X2 U4966 ( .A1(n4497), .A2(n7311), .ZN(n7318) );
  AOI21_X2 U4967 ( .B1(n7316), .B2(n4794), .A(n7315), .ZN(n7317) );
  INV_X4 U4968 ( .A(n4884), .ZN(n4852) );
  INV_X4 U4969 ( .A(n4883), .ZN(n4849) );
  AOI21_X2 U4970 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(n7403) );
  NOR2_X2 U4971 ( .A1(n7401), .A2(n7400), .ZN(n7402) );
  INV_X4 U4972 ( .A(n4884), .ZN(n4854) );
  NOR2_X2 U4973 ( .A1(n4501), .A2(n7408), .ZN(n7417) );
  AOI21_X2 U4974 ( .B1(n7415), .B2(n4794), .A(n7414), .ZN(n7416) );
  INV_X4 U4975 ( .A(n4882), .ZN(n4846) );
  AND2_X4 U4976 ( .A1(n7430), .A2(n4083), .ZN(n4076) );
  AND2_X4 U4977 ( .A1(n8482), .A2(n9050), .ZN(n4077) );
  INV_X4 U4978 ( .A(rst), .ZN(n4886) );
  INV_X4 U4979 ( .A(n4889), .ZN(n4870) );
  AND2_X4 U4980 ( .A1(n5225), .A2(n5232), .ZN(n4078) );
  AND2_X4 U4981 ( .A1(n8173), .A2(n4838), .ZN(n4079) );
  AND2_X4 U4982 ( .A1(n8116), .A2(n4087), .ZN(n4080) );
  INV_X4 U4983 ( .A(n7728), .ZN(n4811) );
  INV_X4 U4984 ( .A(n7732), .ZN(n4826) );
  INV_X4 U4985 ( .A(n4821), .ZN(n4818) );
  NAND3_X2 U4986 ( .A1(n9050), .A2(n9051), .A3(n4133), .ZN(n7674) );
  AND2_X4 U4987 ( .A1(n4731), .A2(n4121), .ZN(n4082) );
  INV_X4 U4988 ( .A(n4790), .ZN(n4788) );
  AND3_X4 U4989 ( .A1(n9050), .A2(n4136), .A3(n9047), .ZN(n4083) );
  INV_X4 U4990 ( .A(rst), .ZN(n4880) );
  INV_X4 U4991 ( .A(n4879), .ZN(n4840) );
  INV_X4 U4992 ( .A(n4879), .ZN(n4839) );
  INV_X4 U4993 ( .A(n4885), .ZN(n4857) );
  INV_X16 U4994 ( .A(n4751), .ZN(n4750) );
  NAND3_X2 U4995 ( .A1(n5260), .A2(n5259), .A3(n5258), .ZN(n4084) );
  NAND3_X2 U4996 ( .A1(n5257), .A2(n5256), .A3(n5255), .ZN(n4085) );
  AND3_X4 U4997 ( .A1(n5121), .A2(n4155), .A3(n5120), .ZN(n4088) );
  AND2_X4 U4998 ( .A1(n4820), .A2(n7841), .ZN(n4089) );
  INV_X4 U4999 ( .A(n4826), .ZN(n4822) );
  INV_X4 U5000 ( .A(n4822), .ZN(n4815) );
  INV_X4 U5001 ( .A(n4822), .ZN(n4816) );
  AND2_X4 U5002 ( .A1(n5483), .A2(n6079), .ZN(n4096) );
  INV_X4 U5003 ( .A(n4077), .ZN(n4805) );
  INV_X4 U5004 ( .A(n4082), .ZN(n4804) );
  AND2_X4 U5005 ( .A1(n5475), .A2(n6338), .ZN(n4097) );
  AND2_X4 U5006 ( .A1(n4331), .A2(n4549), .ZN(n4098) );
  INV_X4 U5007 ( .A(n7299), .ZN(n4778) );
  INV_X4 U5008 ( .A(n4778), .ZN(n4772) );
  NAND3_X2 U5009 ( .A1(n5266), .A2(n5265), .A3(n5264), .ZN(n4099) );
  NAND3_X2 U5010 ( .A1(n5254), .A2(n5253), .A3(n5252), .ZN(n4100) );
  AND3_X4 U5011 ( .A1(n9057), .A2(n9054), .A3(n4139), .ZN(n4101) );
  AND3_X4 U5012 ( .A1(n9058), .A2(n4838), .A3(n4140), .ZN(n4102) );
  INV_X4 U5013 ( .A(n4169), .ZN(n7273) );
  AND2_X4 U5014 ( .A1(n4099), .A2(n7661), .ZN(n4103) );
  INV_X4 U5015 ( .A(n6078), .ZN(n4747) );
  INV_X4 U5016 ( .A(n4079), .ZN(n4837) );
  NAND3_X2 U5017 ( .A1(n5278), .A2(n5277), .A3(n5276), .ZN(n4107) );
  NAND3_X2 U5018 ( .A1(n5251), .A2(n5250), .A3(n5249), .ZN(n4108) );
  AND2_X4 U5019 ( .A1(n8460), .A2(n4099), .ZN(n4110) );
  AND2_X4 U5020 ( .A1(n7895), .A2(n4099), .ZN(n4111) );
  AND2_X4 U5021 ( .A1(n8448), .A2(n4099), .ZN(n4112) );
  AND2_X4 U5022 ( .A1(n8349), .A2(n4099), .ZN(n4113) );
  AND2_X4 U5023 ( .A1(n8348), .A2(n4099), .ZN(n4114) );
  AND2_X4 U5024 ( .A1(n7723), .A2(n4099), .ZN(n4115) );
  AND2_X4 U5025 ( .A1(n8349), .A2(n4100), .ZN(n4116) );
  AND2_X4 U5026 ( .A1(n8348), .A2(n4100), .ZN(n4117) );
  AND2_X4 U5027 ( .A1(n7663), .A2(n4770), .ZN(n4118) );
  NAND2_X2 U5028 ( .A1(n7548), .A2(n7211), .ZN(n7393) );
  INV_X4 U5029 ( .A(n7241), .ZN(n7361) );
  OR2_X4 U5030 ( .A1(n8428), .A2(n4317), .ZN(n4122) );
  AND2_X4 U5031 ( .A1(n8336), .A2(n4100), .ZN(n4123) );
  AND2_X4 U5032 ( .A1(n7123), .A2(n7487), .ZN(n4124) );
  AND2_X4 U5033 ( .A1(n8348), .A2(n4108), .ZN(n4125) );
  OAI21_X2 U5034 ( .B1(n5884), .B2(n5883), .A(not_trap_3), .ZN(n7666) );
  AND4_X4 U5035 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n4126)
         );
  INV_X4 U5036 ( .A(n4822), .ZN(n4820) );
  OR2_X4 U5037 ( .A1(n7393), .A2(n5941), .ZN(n4127) );
  NAND2_X2 U5038 ( .A1(n7211), .A2(n5935), .ZN(n4128) );
  INV_X4 U5039 ( .A(n6625), .ZN(n4769) );
  INV_X4 U5040 ( .A(n6625), .ZN(n4768) );
  AND2_X4 U5041 ( .A1(n5483), .A2(n4080), .ZN(n4132) );
  INV_X4 U5042 ( .A(n4543), .ZN(n4831) );
  INV_X4 U5043 ( .A(n4543), .ZN(n4830) );
  AND2_X4 U5044 ( .A1(n8848), .A2(n4549), .ZN(n4134) );
  NOR2_X2 U5045 ( .A1(n8477), .A2(n4130), .ZN(n7554) );
  INV_X4 U5046 ( .A(n4097), .ZN(n4791) );
  INV_X4 U5047 ( .A(n4790), .ZN(n4785) );
  INV_X4 U5048 ( .A(n4790), .ZN(n4786) );
  INV_X4 U5049 ( .A(n4790), .ZN(n4787) );
  INV_X4 U5050 ( .A(n4098), .ZN(n4834) );
  INV_X4 U5051 ( .A(n4098), .ZN(n4835) );
  INV_X4 U5052 ( .A(n4783), .ZN(n4782) );
  INV_X4 U5053 ( .A(n4783), .ZN(n4781) );
  INV_X4 U5054 ( .A(n4783), .ZN(n4780) );
  INV_X4 U5055 ( .A(n4802), .ZN(n4803) );
  INV_X4 U5056 ( .A(rst), .ZN(n4879) );
  INV_X4 U5057 ( .A(n4885), .ZN(n4859) );
  INV_X4 U5058 ( .A(n4885), .ZN(n4858) );
  INV_X4 U5059 ( .A(n4885), .ZN(n4855) );
  INV_X4 U5060 ( .A(n4743), .ZN(n4742) );
  AND2_X4 U5061 ( .A1(n7648), .A2(n4099), .ZN(n4141) );
  AND2_X4 U5062 ( .A1(n4099), .A2(n7665), .ZN(n4142) );
  AND2_X4 U5063 ( .A1(n4099), .A2(n7657), .ZN(n4143) );
  AND2_X4 U5064 ( .A1(n4099), .A2(n7617), .ZN(n4144) );
  AND2_X4 U5065 ( .A1(n4099), .A2(n4737), .ZN(n4145) );
  AND2_X4 U5066 ( .A1(n4099), .A2(n6365), .ZN(n4146) );
  AND2_X4 U5067 ( .A1(n7623), .A2(n4099), .ZN(n4147) );
  NAND3_X2 U5068 ( .A1(n4914), .A2(n4437), .A3(n4913), .ZN(n7628) );
  AND2_X4 U5069 ( .A1(n7628), .A2(n4099), .ZN(n4148) );
  AND2_X4 U5070 ( .A1(n7634), .A2(n4099), .ZN(n4149) );
  AND2_X4 U5071 ( .A1(n7663), .A2(n4099), .ZN(n4150) );
  AND2_X4 U5072 ( .A1(n7659), .A2(n4099), .ZN(n4151) );
  XOR2_X2 U5073 ( .A(n7423), .B(n4381), .Z(n4152) );
  AND2_X4 U5074 ( .A1(n4084), .A2(n7617), .ZN(n4153) );
  NAND3_X2 U5075 ( .A1(n5089), .A2(n4439), .A3(n5088), .ZN(n6365) );
  AND2_X4 U5076 ( .A1(n4084), .A2(n4737), .ZN(n4154) );
  OR2_X4 U5077 ( .A1(n8977), .A2(n4730), .ZN(n4155) );
  NAND3_X2 U5078 ( .A1(n5217), .A2(n4384), .A3(n5216), .ZN(n7661) );
  AND2_X4 U5079 ( .A1(n7663), .A2(n4085), .ZN(n4157) );
  AND2_X4 U5080 ( .A1(n7665), .A2(n4085), .ZN(n4158) );
  AND2_X4 U5081 ( .A1(n4084), .A2(n7212), .ZN(n4159) );
  AND2_X4 U5082 ( .A1(n4085), .A2(n7212), .ZN(n4160) );
  AND2_X4 U5083 ( .A1(n4084), .A2(n7657), .ZN(n4161) );
  AND2_X4 U5084 ( .A1(n7273), .A2(n7360), .ZN(n4162) );
  AND2_X4 U5085 ( .A1(n4084), .A2(n7663), .ZN(n4163) );
  AND2_X4 U5086 ( .A1(n4084), .A2(n7659), .ZN(n4164) );
  AND2_X4 U5087 ( .A1(n4084), .A2(n7665), .ZN(n4165) );
  AND2_X4 U5088 ( .A1(n7244), .A2(n7273), .ZN(n4166) );
  AND2_X4 U5089 ( .A1(n4084), .A2(n7661), .ZN(n4167) );
  XOR2_X2 U5090 ( .A(n7321), .B(n7267), .Z(n4168) );
  NOR2_X2 U5091 ( .A1(zeroExt_2), .A2(n6619), .ZN(n6079) );
  NAND2_X2 U5092 ( .A1(n5225), .A2(n5226), .ZN(n4169) );
  NOR2_X2 U5093 ( .A1(zeroExt_2), .A2(n6622), .ZN(n6078) );
  INV_X4 U5094 ( .A(n4107), .ZN(n4751) );
  INV_X4 U5095 ( .A(n4078), .ZN(n4784) );
  AND2_X4 U5096 ( .A1(n8304), .A2(n4750), .ZN(n4178) );
  AND2_X4 U5097 ( .A1(n7648), .A2(n4084), .ZN(n4179) );
  AND2_X4 U5098 ( .A1(n7648), .A2(n4085), .ZN(n4180) );
  AND2_X4 U5099 ( .A1(n7648), .A2(n4100), .ZN(n4181) );
  AND2_X4 U5100 ( .A1(n7648), .A2(n4108), .ZN(n4182) );
  AND2_X4 U5101 ( .A1(n4099), .A2(n8364), .ZN(n4183) );
  AND2_X4 U5102 ( .A1(n4099), .A2(n8326), .ZN(n4184) );
  AND2_X4 U5103 ( .A1(n4099), .A2(n7722), .ZN(n4185) );
  AND2_X4 U5104 ( .A1(n4099), .A2(n7720), .ZN(n4186) );
  AND2_X4 U5105 ( .A1(n7623), .A2(n4084), .ZN(n4187) );
  AND2_X4 U5106 ( .A1(n7623), .A2(n4085), .ZN(n4188) );
  AND2_X4 U5107 ( .A1(n7623), .A2(n4100), .ZN(n4189) );
  AND2_X4 U5108 ( .A1(n7623), .A2(n4108), .ZN(n4190) );
  AND2_X4 U5109 ( .A1(n4100), .A2(n7212), .ZN(n4191) );
  AND2_X4 U5110 ( .A1(n4100), .A2(n7661), .ZN(n4192) );
  AND2_X4 U5111 ( .A1(n4100), .A2(n7657), .ZN(n4193) );
  AND2_X4 U5112 ( .A1(n4100), .A2(n7617), .ZN(n4194) );
  AND2_X4 U5113 ( .A1(n4100), .A2(n4737), .ZN(n4195) );
  AND2_X4 U5114 ( .A1(n4100), .A2(n6365), .ZN(n4196) );
  AND2_X4 U5115 ( .A1(n4108), .A2(n7665), .ZN(n4197) );
  AND2_X4 U5116 ( .A1(n4108), .A2(n7663), .ZN(n4198) );
  AND2_X4 U5117 ( .A1(n4108), .A2(n7661), .ZN(n4199) );
  AND2_X4 U5118 ( .A1(n4108), .A2(n7659), .ZN(n4200) );
  AND2_X4 U5119 ( .A1(n4108), .A2(n7657), .ZN(n4201) );
  AND2_X4 U5120 ( .A1(n4108), .A2(n7617), .ZN(n4202) );
  AND2_X4 U5121 ( .A1(n4108), .A2(n4737), .ZN(n4203) );
  AND2_X4 U5122 ( .A1(n4108), .A2(n6365), .ZN(n4204) );
  AND2_X4 U5123 ( .A1(n5589), .A2(n5588), .ZN(n4205) );
  AND2_X4 U5124 ( .A1(n7641), .A2(n4099), .ZN(n4210) );
  AND2_X4 U5125 ( .A1(n7726), .A2(n4099), .ZN(n4211) );
  AND2_X4 U5126 ( .A1(n8336), .A2(n4099), .ZN(n4212) );
  AND2_X4 U5127 ( .A1(n7721), .A2(n4099), .ZN(n4213) );
  AND2_X4 U5128 ( .A1(n4085), .A2(n7617), .ZN(n4214) );
  AND2_X4 U5129 ( .A1(n4770), .A2(n7617), .ZN(n4215) );
  AND2_X4 U5130 ( .A1(n7663), .A2(n4100), .ZN(n4216) );
  AND2_X4 U5131 ( .A1(n7659), .A2(n4100), .ZN(n4217) );
  AND2_X4 U5132 ( .A1(n7628), .A2(n4100), .ZN(n4218) );
  AND2_X4 U5133 ( .A1(n7634), .A2(n4100), .ZN(n4219) );
  AND2_X4 U5134 ( .A1(n7641), .A2(n4100), .ZN(n4220) );
  AND2_X4 U5135 ( .A1(n7726), .A2(n4100), .ZN(n4221) );
  AND2_X4 U5136 ( .A1(n8460), .A2(n4100), .ZN(n4222) );
  AND2_X4 U5137 ( .A1(n7895), .A2(n4100), .ZN(n4223) );
  AND2_X4 U5138 ( .A1(n8448), .A2(n4100), .ZN(n4224) );
  AND2_X4 U5139 ( .A1(n7628), .A2(n4108), .ZN(n4225) );
  AND2_X4 U5140 ( .A1(n7634), .A2(n4108), .ZN(n4226) );
  AND2_X4 U5141 ( .A1(n7641), .A2(n4108), .ZN(n4227) );
  AND2_X4 U5142 ( .A1(n4085), .A2(n4737), .ZN(n4228) );
  AND2_X4 U5143 ( .A1(n7266), .A2(n4737), .ZN(n4229) );
  AND2_X4 U5144 ( .A1(n7641), .A2(n4084), .ZN(n4230) );
  AND2_X4 U5145 ( .A1(n7641), .A2(n4085), .ZN(n4231) );
  AND2_X4 U5146 ( .A1(n7723), .A2(n4084), .ZN(n4232) );
  AND2_X4 U5147 ( .A1(n7628), .A2(n4084), .ZN(n4233) );
  AND2_X4 U5148 ( .A1(n7628), .A2(n4085), .ZN(n4234) );
  AND2_X4 U5149 ( .A1(n7634), .A2(n4084), .ZN(n4235) );
  AND2_X4 U5150 ( .A1(n7634), .A2(n4085), .ZN(n4236) );
  AND2_X4 U5151 ( .A1(n7726), .A2(n4084), .ZN(n4237) );
  AND2_X4 U5152 ( .A1(n7726), .A2(n4085), .ZN(n4238) );
  AND2_X4 U5153 ( .A1(n8460), .A2(n4084), .ZN(n4239) );
  AND2_X4 U5154 ( .A1(n8460), .A2(n4085), .ZN(n4240) );
  AND2_X4 U5155 ( .A1(n8348), .A2(n4084), .ZN(n4241) );
  AND2_X4 U5156 ( .A1(n8348), .A2(n4085), .ZN(n4242) );
  AND2_X4 U5157 ( .A1(n8448), .A2(n4084), .ZN(n4243) );
  AND2_X4 U5158 ( .A1(n8448), .A2(n4085), .ZN(n4244) );
  AND2_X4 U5159 ( .A1(n7659), .A2(n4085), .ZN(n4245) );
  AND2_X4 U5160 ( .A1(n7659), .A2(n4770), .ZN(n4246) );
  AND2_X4 U5161 ( .A1(n7665), .A2(n7266), .ZN(n4247) );
  AND2_X4 U5162 ( .A1(n7721), .A2(n4084), .ZN(n4248) );
  AND2_X4 U5163 ( .A1(n8349), .A2(n4084), .ZN(n4249) );
  AND2_X4 U5164 ( .A1(n8349), .A2(n4085), .ZN(n4250) );
  AND2_X4 U5165 ( .A1(n8336), .A2(n4085), .ZN(n4251) );
  AND2_X4 U5166 ( .A1(n7895), .A2(n4084), .ZN(n4252) );
  AND2_X4 U5167 ( .A1(n7895), .A2(n4085), .ZN(n4253) );
  AND2_X4 U5168 ( .A1(n7266), .A2(n7212), .ZN(n4254) );
  AND2_X4 U5169 ( .A1(n8336), .A2(n4084), .ZN(n4255) );
  AND2_X4 U5170 ( .A1(n4084), .A2(n8364), .ZN(n4256) );
  AND2_X4 U5171 ( .A1(n4085), .A2(n8364), .ZN(n4257) );
  AND2_X4 U5172 ( .A1(n4085), .A2(n7657), .ZN(n4258) );
  AND2_X4 U5173 ( .A1(n4770), .A2(n7657), .ZN(n4259) );
  AND2_X4 U5174 ( .A1(n4084), .A2(n6365), .ZN(n4260) );
  AND2_X4 U5175 ( .A1(n4085), .A2(n6365), .ZN(n4261) );
  AND2_X4 U5176 ( .A1(n7266), .A2(n6365), .ZN(n4262) );
  AND2_X4 U5177 ( .A1(n4084), .A2(n8326), .ZN(n4263) );
  AND2_X4 U5178 ( .A1(n4085), .A2(n8326), .ZN(n4264) );
  AND2_X4 U5179 ( .A1(ex_multing_set_product_in_sig_z1[10]), .A2(n4784), .ZN(
        n4265) );
  AND2_X4 U5180 ( .A1(n4084), .A2(n7722), .ZN(n4266) );
  AND2_X4 U5181 ( .A1(n7273), .A2(n6884), .ZN(n4267) );
  AND2_X4 U5182 ( .A1(n7273), .A2(n7046), .ZN(n4268) );
  AND2_X4 U5183 ( .A1(n4085), .A2(n7661), .ZN(n4269) );
  AND2_X4 U5184 ( .A1(n4770), .A2(n7661), .ZN(n4270) );
  XOR2_X2 U5185 ( .A(n6067), .B(iAddr[30]), .Z(n4271) );
  AND2_X4 U5186 ( .A1(n4175), .A2(n4452), .ZN(n4272) );
  AND2_X4 U5187 ( .A1(n4467), .A2(n4452), .ZN(n4273) );
  AND2_X4 U5188 ( .A1(n4177), .A2(n4452), .ZN(n4274) );
  INV_X4 U5189 ( .A(n7123), .ZN(n4744) );
  NAND3_X2 U5190 ( .A1(n5245), .A2(n5244), .A3(n5243), .ZN(n7266) );
  INV_X4 U5191 ( .A(n7266), .ZN(n4771) );
  AND2_X4 U5192 ( .A1(n7648), .A2(n4770), .ZN(n4281) );
  AND2_X4 U5193 ( .A1(n7623), .A2(n4770), .ZN(n4282) );
  AND2_X4 U5194 ( .A1(n4100), .A2(n8364), .ZN(n4283) );
  AND2_X4 U5195 ( .A1(n4100), .A2(n8326), .ZN(n4284) );
  AND2_X4 U5196 ( .A1(n4108), .A2(n8364), .ZN(n4285) );
  AND2_X4 U5197 ( .A1(n4108), .A2(n8326), .ZN(n4286) );
  OR2_X4 U5198 ( .A1(n7207), .A2(n7216), .ZN(n4287) );
  AND2_X4 U5199 ( .A1(n7723), .A2(n4100), .ZN(n4288) );
  AND2_X4 U5200 ( .A1(n7726), .A2(n4108), .ZN(n4289) );
  AND2_X4 U5201 ( .A1(n8460), .A2(n4108), .ZN(n4290) );
  AND2_X4 U5202 ( .A1(n7895), .A2(n4108), .ZN(n4291) );
  AND2_X4 U5203 ( .A1(n8448), .A2(n4108), .ZN(n4292) );
  AND2_X4 U5204 ( .A1(n8349), .A2(n4108), .ZN(n4293) );
  AND2_X4 U5205 ( .A1(n8336), .A2(n4108), .ZN(n4294) );
  AND2_X4 U5206 ( .A1(n7962), .A2(n7490), .ZN(n4295) );
  AND2_X4 U5207 ( .A1(n7641), .A2(n4770), .ZN(n4296) );
  AND2_X4 U5208 ( .A1(n7723), .A2(n4085), .ZN(n4297) );
  AND2_X4 U5209 ( .A1(n7628), .A2(n4770), .ZN(n4298) );
  AND2_X4 U5210 ( .A1(n7634), .A2(n4770), .ZN(n4299) );
  AND2_X4 U5211 ( .A1(n7726), .A2(n4770), .ZN(n4300) );
  AND2_X4 U5212 ( .A1(n8460), .A2(n4770), .ZN(n4301) );
  AND2_X4 U5213 ( .A1(n8348), .A2(n4770), .ZN(n4302) );
  AND2_X4 U5214 ( .A1(n8448), .A2(n4770), .ZN(n4303) );
  AND2_X4 U5215 ( .A1(n7266), .A2(n8364), .ZN(n4304) );
  AND2_X4 U5216 ( .A1(ex_multing_set_product_in_sig_z1[12]), .A2(n4784), .ZN(
        n4305) );
  AND2_X4 U5217 ( .A1(ex_multing_set_product_in_sig_z1[18]), .A2(n4784), .ZN(
        n4306) );
  AND2_X4 U5218 ( .A1(ex_multing_set_product_in_sig_z1[20]), .A2(n4784), .ZN(
        n4307) );
  AND2_X4 U5219 ( .A1(ex_multing_set_product_in_sig_z1[22]), .A2(n4784), .ZN(
        n4308) );
  AND2_X4 U5220 ( .A1(ex_multing_set_product_in_sig_z1[26]), .A2(n4784), .ZN(
        n4309) );
  AND2_X4 U5221 ( .A1(ex_multing_set_product_in_sig_z1[28]), .A2(n4784), .ZN(
        n4310) );
  AND2_X4 U5222 ( .A1(n4085), .A2(n7722), .ZN(n4311) );
  AND2_X4 U5223 ( .A1(n5925), .A2(n5935), .ZN(n4312) );
  AND2_X4 U5224 ( .A1(n4784), .A2(n4561), .ZN(n4313) );
  AND2_X4 U5225 ( .A1(n4784), .A2(n4570), .ZN(n4314) );
  AND2_X4 U5226 ( .A1(n4784), .A2(n4571), .ZN(n4315) );
  AND2_X4 U5227 ( .A1(n4784), .A2(n4572), .ZN(n4316) );
  OAI21_X2 U5228 ( .B1(n6071), .B2(n4898), .A(n5882), .ZN(n7732) );
  NAND2_X2 U5229 ( .A1(n7548), .A2(n5925), .ZN(n4317) );
  INV_X4 U5230 ( .A(n7728), .ZN(n4807) );
  NAND3_X2 U5231 ( .A1(n4744), .A2(n5882), .A3(n5799), .ZN(n7728) );
  INV_X4 U5232 ( .A(n4807), .ZN(n4806) );
  INV_X4 U5233 ( .A(n4089), .ZN(n4827) );
  INV_X4 U5234 ( .A(n7164), .ZN(n4757) );
  INV_X4 U5235 ( .A(n5978), .ZN(n7209) );
  INV_X4 U5236 ( .A(n4735), .ZN(n4736) );
  NAND2_X2 U5237 ( .A1(n4082), .A2(n4091), .ZN(n7896) );
  INV_X4 U5238 ( .A(n7674), .ZN(n4731) );
  INV_X4 U5239 ( .A(n4134), .ZN(n4833) );
  INV_X4 U5240 ( .A(n4134), .ZN(n4832) );
  INV_X4 U5241 ( .A(n7554), .ZN(n4728) );
  INV_X4 U5242 ( .A(n4728), .ZN(n4729) );
  INV_X4 U5243 ( .A(n4803), .ZN(n4801) );
  INV_X4 U5244 ( .A(n4803), .ZN(n4797) );
  INV_X4 U5245 ( .A(n4803), .ZN(n4796) );
  INV_X4 U5246 ( .A(n4782), .ZN(n4773) );
  INV_X4 U5247 ( .A(n4783), .ZN(n4779) );
  INV_X4 U5248 ( .A(rst), .ZN(n4885) );
  INV_X4 U5249 ( .A(n4888), .ZN(n4867) );
  INV_X4 U5250 ( .A(n4888), .ZN(n4866) );
  INV_X4 U5251 ( .A(n4888), .ZN(n4865) );
  OAI21_X2 U5252 ( .B1(n9048), .B2(n4136), .A(n9047), .ZN(n8536) );
  INV_X4 U5253 ( .A(n8536), .ZN(n8605) );
  NAND3_X2 U5254 ( .A1(n4934), .A2(n4933), .A3(n4932), .ZN(n7648) );
  NAND3_X2 U5255 ( .A1(n5224), .A2(n5223), .A3(n5222), .ZN(n7617) );
  XNOR2_X2 U5256 ( .A(n8298), .B(n8299), .ZN(n4374) );
  OR2_X4 U5257 ( .A1(n4369), .A2(n5210), .ZN(n4375) );
  OR2_X4 U5258 ( .A1(n7604), .A2(n4742), .ZN(n4376) );
  OR2_X4 U5259 ( .A1(n7601), .A2(n4742), .ZN(n4377) );
  OR2_X4 U5260 ( .A1(n7583), .A2(n5211), .ZN(n4378) );
  OR2_X4 U5261 ( .A1(n7586), .A2(n4742), .ZN(n4379) );
  OR2_X4 U5262 ( .A1(n7584), .A2(n4742), .ZN(n4380) );
  XOR2_X2 U5263 ( .A(n8605), .B(n7430), .Z(n4381) );
  OR2_X4 U5264 ( .A1(n8982), .A2(n4730), .ZN(n4382) );
  OR2_X4 U5265 ( .A1(n8981), .A2(n4730), .ZN(n4383) );
  OR2_X4 U5266 ( .A1(n8980), .A2(n4730), .ZN(n4384) );
  OR2_X4 U5267 ( .A1(n8979), .A2(n4730), .ZN(n4385) );
  OR2_X4 U5268 ( .A1(n8978), .A2(n4730), .ZN(n4386) );
  XOR2_X2 U5269 ( .A(n8605), .B(n5925), .Z(n4387) );
  XOR2_X2 U5270 ( .A(n6551), .B(n6550), .Z(n4389) );
  NOR3_X2 U5271 ( .A1(n4901), .A2(n7597), .A3(n4086), .ZN(n5170) );
  NOR3_X2 U5272 ( .A1(n4900), .A2(n7595), .A3(n4104), .ZN(n4936) );
  INV_X4 U5273 ( .A(n4102), .ZN(n4733) );
  INV_X4 U5274 ( .A(n4101), .ZN(n4732) );
  AND2_X4 U5275 ( .A1(n4138), .A2(n4452), .ZN(n4392) );
  AND2_X4 U5276 ( .A1(n5625), .A2(n4750), .ZN(n4393) );
  AND2_X4 U5277 ( .A1(n6087), .A2(n4750), .ZN(n4394) );
  AND2_X4 U5278 ( .A1(n5749), .A2(n4107), .ZN(n4395) );
  AND2_X4 U5279 ( .A1(n6097), .A2(n4107), .ZN(n4396) );
  INV_X4 U5280 ( .A(n5210), .ZN(n4741) );
  INV_X4 U5281 ( .A(n5210), .ZN(n4740) );
  INV_X4 U5282 ( .A(n4747), .ZN(n4746) );
  INV_X4 U5283 ( .A(n5029), .ZN(n4739) );
  INV_X4 U5284 ( .A(n6157), .ZN(n4754) );
  NAND3_X2 U5285 ( .A1(n5235), .A2(n5234), .A3(n5233), .ZN(n6157) );
  INV_X4 U5286 ( .A(n4107), .ZN(n4752) );
  AND2_X4 U5287 ( .A1(n4753), .A2(n8306), .ZN(n4416) );
  OR2_X4 U5288 ( .A1(n4409), .A2(n5210), .ZN(n4419) );
  OR2_X4 U5289 ( .A1(n4410), .A2(n5210), .ZN(n4420) );
  OR2_X4 U5290 ( .A1(n4411), .A2(n5210), .ZN(n4421) );
  OR2_X4 U5291 ( .A1(n4412), .A2(n5210), .ZN(n4422) );
  OR2_X4 U5292 ( .A1(n7603), .A2(n4742), .ZN(n4423) );
  OR2_X4 U5293 ( .A1(n7575), .A2(n4742), .ZN(n4424) );
  OR2_X4 U5294 ( .A1(n7581), .A2(n5211), .ZN(n4425) );
  OR2_X4 U5295 ( .A1(n7588), .A2(n5211), .ZN(n4426) );
  OR2_X4 U5296 ( .A1(n7602), .A2(n5211), .ZN(n4427) );
  OR2_X4 U5297 ( .A1(n7598), .A2(n4742), .ZN(n4428) );
  OR2_X4 U5298 ( .A1(n8947), .A2(n4730), .ZN(n4429) );
  OR2_X4 U5299 ( .A1(n9030), .A2(n4730), .ZN(n4430) );
  OR2_X4 U5300 ( .A1(n9036), .A2(n4730), .ZN(n4431) );
  OR2_X4 U5301 ( .A1(n9033), .A2(n4730), .ZN(n4432) );
  OR2_X4 U5302 ( .A1(n8948), .A2(n4730), .ZN(n4433) );
  OR2_X4 U5303 ( .A1(n8949), .A2(n4730), .ZN(n4434) );
  OR2_X4 U5304 ( .A1(n8951), .A2(n4730), .ZN(n4435) );
  OR2_X4 U5305 ( .A1(n8952), .A2(n4730), .ZN(n4436) );
  OR2_X4 U5306 ( .A1(n8984), .A2(n4730), .ZN(n4437) );
  OR2_X4 U5307 ( .A1(n8983), .A2(n4730), .ZN(n4438) );
  OR2_X4 U5308 ( .A1(n8976), .A2(n4730), .ZN(n4439) );
  OR2_X4 U5309 ( .A1(n8950), .A2(n4730), .ZN(n4440) );
  NAND3_X2 U5310 ( .A1(n7596), .A2(n7595), .A3(n4899), .ZN(n5211) );
  INV_X4 U5311 ( .A(n5211), .ZN(n4743) );
  XOR2_X2 U5312 ( .A(n4178), .B(n4416), .Z(n4442) );
  AND2_X4 U5313 ( .A1(n4176), .A2(n4452), .ZN(n4443) );
  AND2_X4 U5314 ( .A1(n4407), .A2(n4452), .ZN(n4444) );
  AND2_X4 U5315 ( .A1(n6107), .A2(n4750), .ZN(n4445) );
  AND2_X4 U5316 ( .A1(n6150), .A2(n4107), .ZN(n4446) );
  INV_X4 U5317 ( .A(n4088), .ZN(n4737) );
  INV_X4 U5318 ( .A(n6079), .ZN(n4749) );
  INV_X4 U5319 ( .A(n4749), .ZN(n4748) );
  OR2_X4 U5320 ( .A1(n7477), .A2(n7476), .ZN(n4451) );
  INV_X4 U5321 ( .A(n4771), .ZN(n4770) );
  INV_X4 U5322 ( .A(n4452), .ZN(n4838) );
  AND2_X4 U5323 ( .A1(n7531), .A2(n7524), .ZN(n4468) );
  XOR2_X2 U5324 ( .A(n8536), .B(n4152), .Z(n4469) );
  OR2_X4 U5325 ( .A1(n8416), .A2(n4734), .ZN(n4470) );
  OR2_X4 U5326 ( .A1(n8428), .A2(n4736), .ZN(n4471) );
  NAND3_X2 U5327 ( .A1(n4908), .A2(n4907), .A3(n4906), .ZN(n7623) );
  NAND3_X2 U5328 ( .A1(n5126), .A2(n5125), .A3(n5124), .ZN(n7479) );
  OR2_X4 U5329 ( .A1(n8362), .A2(n4128), .ZN(n4472) );
  OR2_X4 U5330 ( .A1(n8393), .A2(n4734), .ZN(n4473) );
  OR2_X4 U5331 ( .A1(n5644), .A2(n4317), .ZN(n4476) );
  OR2_X4 U5332 ( .A1(n8946), .A2(n4730), .ZN(n4477) );
  AND2_X4 U5333 ( .A1(n7492), .A2(n7687), .ZN(n4478) );
  AND2_X4 U5334 ( .A1(ex_multing_set_product_in_sig_z1[8]), .A2(n4784), .ZN(
        n4479) );
  AND2_X4 U5335 ( .A1(n7295), .A2(n7491), .ZN(n4494) );
  INV_X4 U5336 ( .A(n6331), .ZN(n4756) );
  INV_X4 U5337 ( .A(n4756), .ZN(n4755) );
  AND2_X4 U5338 ( .A1(n7492), .A2(n7980), .ZN(n4495) );
  AND2_X4 U5339 ( .A1(n7492), .A2(n7675), .ZN(n4496) );
  AND2_X4 U5340 ( .A1(n7492), .A2(n7887), .ZN(n4497) );
  XOR2_X2 U5341 ( .A(n6330), .B(n6329), .Z(n4498) );
  OR2_X4 U5342 ( .A1(n8418), .A2(n7563), .ZN(n4499) );
  OR2_X4 U5343 ( .A1(n7658), .A2(n4728), .ZN(n4500) );
  AND2_X4 U5344 ( .A1(n7492), .A2(n7913), .ZN(n4501) );
  AND2_X4 U5345 ( .A1(n7492), .A2(n7699), .ZN(n4502) );
  AND2_X4 U5346 ( .A1(n7492), .A2(n7709), .ZN(n4503) );
  OR2_X4 U5347 ( .A1(n8486), .A2(n7501), .ZN(n4504) );
  AND2_X4 U5348 ( .A1(n7385), .A2(n7525), .ZN(n4505) );
  INV_X4 U5349 ( .A(n7666), .ZN(n4793) );
  OR2_X4 U5350 ( .A1(n7656), .A2(n4728), .ZN(n4506) );
  AND2_X4 U5351 ( .A1(n4085), .A2(n7720), .ZN(n4507) );
  OR2_X4 U5352 ( .A1(n5944), .A2(n4734), .ZN(n4508) );
  AND2_X4 U5353 ( .A1(n7492), .A2(n7295), .ZN(n4509) );
  INV_X4 U5354 ( .A(n7732), .ZN(n4825) );
  INV_X4 U5355 ( .A(n4825), .ZN(n4823) );
  INV_X4 U5356 ( .A(n4825), .ZN(n4824) );
  INV_X4 U5357 ( .A(n4826), .ZN(n4821) );
  INV_X4 U5358 ( .A(n4080), .ZN(n4730) );
  OR2_X4 U5359 ( .A1(n8401), .A2(n4738), .ZN(n4523) );
  INV_X4 U5360 ( .A(n4806), .ZN(n4809) );
  INV_X4 U5361 ( .A(n4806), .ZN(n4808) );
  INV_X4 U5362 ( .A(n4089), .ZN(n4829) );
  INV_X4 U5363 ( .A(n4089), .ZN(n4828) );
  INV_X4 U5364 ( .A(n4811), .ZN(n4810) );
  AND2_X4 U5365 ( .A1(n8849), .A2(n4331), .ZN(n4543) );
  NAND3_X2 U5366 ( .A1(n5137), .A2(n5136), .A3(n5135), .ZN(n8019) );
  INV_X4 U5367 ( .A(n8019), .ZN(n7525) );
  AND2_X4 U5368 ( .A1(n4744), .A2(n6338), .ZN(n4558) );
  AND2_X4 U5369 ( .A1(n8128), .A2(n8931), .ZN(n4562) );
  OAI21_X2 U5370 ( .B1(n8986), .B2(n4893), .A(n8985), .ZN(n7123) );
  AND2_X4 U5371 ( .A1(n6258), .A2(n7546), .ZN(n4563) );
  INV_X4 U5372 ( .A(n7362), .ZN(n7243) );
  NAND3_X2 U5373 ( .A1(n4952), .A2(n4951), .A3(n4950), .ZN(n7379) );
  INV_X4 U5374 ( .A(n8340), .ZN(n7489) );
  INV_X4 U5375 ( .A(n7393), .ZN(n4735) );
  NAND2_X2 U5376 ( .A1(n7422), .A2(n4083), .ZN(n7216) );
  AND2_X4 U5377 ( .A1(n8018), .A2(n7565), .ZN(n4585) );
  OAI21_X2 U5378 ( .B1(n4747), .B2(n7191), .A(n4783), .ZN(n7677) );
  OR2_X4 U5379 ( .A1(n7660), .A2(n4728), .ZN(n4586) );
  NOR2_X2 U5380 ( .A1(n4805), .A2(n4130), .ZN(n7412) );
  AND2_X4 U5381 ( .A1(n4784), .A2(n4573), .ZN(n4587) );
  INV_X4 U5382 ( .A(n7163), .ZN(n4763) );
  INV_X4 U5383 ( .A(n4763), .ZN(n4761) );
  INV_X4 U5384 ( .A(n4763), .ZN(n4762) );
  NOR3_X2 U5385 ( .A1(n4786), .A2(n9057), .A3(n4139), .ZN(n7163) );
  AND4_X4 U5386 ( .A1(n8129), .A2(n6071), .A3(n4562), .A4(n6070), .ZN(n4591)
         );
  INV_X4 U5387 ( .A(n7162), .ZN(n4760) );
  INV_X4 U5388 ( .A(n4760), .ZN(n4758) );
  INV_X4 U5389 ( .A(n4760), .ZN(n4759) );
  NOR3_X2 U5390 ( .A1(n4785), .A2(n9058), .A3(n4140), .ZN(n7162) );
  INV_X4 U5391 ( .A(n7615), .ZN(n4794) );
  INV_X4 U5392 ( .A(n6332), .ZN(n4745) );
  AND3_X4 U5393 ( .A1(n8129), .A2(n6072), .A3(n4562), .ZN(n4592) );
  INV_X4 U5394 ( .A(n6621), .ZN(n4764) );
  INV_X4 U5395 ( .A(n6621), .ZN(n4765) );
  INV_X4 U5396 ( .A(n6624), .ZN(n4766) );
  INV_X4 U5397 ( .A(n6624), .ZN(n4767) );
  OR2_X4 U5398 ( .A1(n7664), .A2(n4728), .ZN(n4594) );
  INV_X4 U5399 ( .A(n4896), .ZN(n4802) );
  INV_X4 U5400 ( .A(n4803), .ZN(n4795) );
  INV_X4 U5401 ( .A(n4128), .ZN(n6258) );
  INV_X4 U5402 ( .A(n4312), .ZN(n4734) );
  INV_X4 U5403 ( .A(n4097), .ZN(n4792) );
  INV_X4 U5404 ( .A(n4097), .ZN(n4790) );
  INV_X4 U5405 ( .A(n4076), .ZN(n4738) );
  INV_X4 U5406 ( .A(n4778), .ZN(n4783) );
  INV_X4 U5407 ( .A(rst), .ZN(n4891) );
  INV_X4 U5408 ( .A(rst), .ZN(n4890) );
  INV_X4 U5409 ( .A(rst), .ZN(n4889) );
  INV_X4 U5410 ( .A(rst), .ZN(n4888) );
  AOI21_X2 U5411 ( .B1(n8523), .B2(n8515), .A(n8516), .ZN(n8520) );
  AOI22_X2 U5412 ( .A1(n7663), .A2(n8644), .B1(n8537), .B2(n8538), .ZN(n8643)
         );
  OAI21_X2 U5413 ( .B1(n7520), .B2(n8645), .A(n8535), .ZN(n8537) );
  INV_X4 U5414 ( .A(n8562), .ZN(n8630) );
  INV_X4 U5415 ( .A(n8625), .ZN(n8590) );
  INV_X4 U5416 ( .A(n8586), .ZN(n8619) );
  INV_X4 U5417 ( .A(n8588), .ZN(n8615) );
  INV_X4 U5418 ( .A(n8622), .ZN(n8576) );
  INV_X4 U5419 ( .A(n8600), .ZN(n8632) );
  INV_X4 U5420 ( .A(n8592), .ZN(n8641) );
  INV_X4 U5421 ( .A(n8596), .ZN(n8638) );
  INV_X4 U5422 ( .A(n8582), .ZN(n8612) );
  INV_X4 U5423 ( .A(n7796), .ZN(n7745) );
  OR3_X4 U5424 ( .A1(n7798), .A2(n7799), .A3(n7764), .ZN(n7765) );
  INV_X4 U5425 ( .A(n8450), .ZN(n8327) );
  XNOR2_X2 U5426 ( .A(op0_3), .B(n4388), .ZN(n4893) );
  NAND2_X2 U5427 ( .A1(n4895), .A2(n4894), .ZN(n4897) );
  NAND2_X2 U5428 ( .A1(n4744), .A2(n4897), .ZN(n6338) );
  NAND2_X2 U5429 ( .A1(n7125), .A2(n4878), .ZN(n4896) );
  INV_X4 U5430 ( .A(n4897), .ZN(n5798) );
  NAND2_X2 U5431 ( .A1(n4744), .A2(n5798), .ZN(n6071) );
  INV_X4 U5432 ( .A(n6338), .ZN(n6072) );
  NAND2_X2 U5433 ( .A1(n5798), .A2(n4091), .ZN(n7615) );
  NAND2_X2 U5434 ( .A1(regWr), .A2(n4106), .ZN(n4899) );
  NAND2_X2 U5435 ( .A1(n4899), .A2(n4104), .ZN(n5210) );
  NAND2_X2 U5436 ( .A1(reg31Val_0[11]), .A2(n4741), .ZN(n4905) );
  NAND2_X2 U5437 ( .A1(n4743), .A2(n4622), .ZN(n4904) );
  INV_X4 U5438 ( .A(n4899), .ZN(n4900) );
  NAND2_X2 U5439 ( .A1(n4936), .A2(n4086), .ZN(n5029) );
  INV_X4 U5440 ( .A(n5029), .ZN(n5209) );
  NAND2_X2 U5441 ( .A1(wb_dsize_reg_z2[11]), .A2(n4739), .ZN(n4903) );
  INV_X4 U5442 ( .A(n4936), .ZN(n4901) );
  NAND2_X2 U5443 ( .A1(wb_dsize_reg_z2[27]), .A2(n5170), .ZN(n4902) );
  NAND4_X2 U5444 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(
        regWrData[11]) );
  NAND2_X2 U5445 ( .A1(n4080), .A2(n4207), .ZN(n4908) );
  NAND2_X2 U5446 ( .A1(n9052), .A2(n4156), .ZN(n6622) );
  NAND2_X2 U5447 ( .A1(n4746), .A2(memAddr[11]), .ZN(n4907) );
  NAND2_X2 U5448 ( .A1(n9053), .A2(n4373), .ZN(n6619) );
  NAND2_X2 U5449 ( .A1(regWrData[11]), .A2(n6079), .ZN(n4906) );
  NAND2_X2 U5450 ( .A1(reg31Val_0[12]), .A2(n4740), .ZN(n4912) );
  NAND2_X2 U5451 ( .A1(n4743), .A2(n4624), .ZN(n4911) );
  NAND2_X2 U5452 ( .A1(wb_dsize_reg_z2[12]), .A2(n4739), .ZN(n4910) );
  NAND2_X2 U5453 ( .A1(wb_dsize_reg_z2[28]), .A2(n5170), .ZN(n4909) );
  NAND4_X2 U5454 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n4909), .ZN(
        regWrData[12]) );
  NAND2_X2 U5455 ( .A1(n6078), .A2(memAddr[12]), .ZN(n4914) );
  NAND2_X2 U5456 ( .A1(regWrData[12]), .A2(n4748), .ZN(n4913) );
  NAND2_X2 U5457 ( .A1(reg31Val_0[13]), .A2(n4740), .ZN(n4918) );
  NAND2_X2 U5458 ( .A1(n4743), .A2(n4447), .ZN(n4917) );
  NAND2_X2 U5459 ( .A1(wb_dsize_reg_z2[13]), .A2(n4739), .ZN(n4916) );
  NAND2_X2 U5460 ( .A1(wb_dsize_reg_z2[29]), .A2(n5170), .ZN(n4915) );
  NAND4_X2 U5461 ( .A1(n4918), .A2(n4917), .A3(n4916), .A4(n4915), .ZN(
        regWrData[13]) );
  NAND2_X2 U5462 ( .A1(n4080), .A2(n4208), .ZN(n4921) );
  NAND2_X2 U5463 ( .A1(n6078), .A2(memAddr[13]), .ZN(n4920) );
  NAND2_X2 U5464 ( .A1(regWrData[13]), .A2(n6079), .ZN(n4919) );
  NAND2_X2 U5465 ( .A1(reg31Val_0[14]), .A2(n4740), .ZN(n4925) );
  NAND2_X2 U5466 ( .A1(n4743), .A2(n4448), .ZN(n4924) );
  NAND2_X2 U5467 ( .A1(wb_dsize_reg_z2[14]), .A2(n4739), .ZN(n4923) );
  NAND2_X2 U5468 ( .A1(wb_dsize_reg_z2[30]), .A2(n5170), .ZN(n4922) );
  NAND4_X2 U5469 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(
        regWrData[14]) );
  NAND2_X2 U5470 ( .A1(n6078), .A2(memAddr[14]), .ZN(n4927) );
  NAND2_X2 U5471 ( .A1(regWrData[14]), .A2(n4748), .ZN(n4926) );
  NAND2_X2 U5472 ( .A1(reg31Val_0[10]), .A2(n4740), .ZN(n4931) );
  NAND2_X2 U5473 ( .A1(n4743), .A2(n4621), .ZN(n4930) );
  NAND2_X2 U5474 ( .A1(wb_dsize_reg_z2[10]), .A2(n4739), .ZN(n4929) );
  NAND2_X2 U5475 ( .A1(wb_dsize_reg_z2[26]), .A2(n5170), .ZN(n4928) );
  NAND4_X2 U5476 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(
        regWrData[10]) );
  NAND2_X2 U5477 ( .A1(n4080), .A2(n4209), .ZN(n4934) );
  NAND2_X2 U5478 ( .A1(n4746), .A2(memAddr[10]), .ZN(n4933) );
  NAND2_X2 U5479 ( .A1(regWrData[10]), .A2(n4748), .ZN(n4932) );
  NAND2_X2 U5480 ( .A1(n5170), .A2(wb_dsize_reg_z2[16]), .ZN(n4938) );
  NAND2_X2 U5481 ( .A1(n5170), .A2(wb_dsize_reg_z2[18]), .ZN(n4942) );
  AOI22_X2 U5482 ( .A1(wb_dsize_reg_z2[2]), .A2(n5209), .B1(
        wb_dsize_reg_z2[26]), .B2(n5171), .ZN(n4941) );
  NAND2_X2 U5483 ( .A1(n5170), .A2(wb_dsize_reg_z2[17]), .ZN(n4946) );
  AOI22_X2 U5484 ( .A1(wb_dsize_reg_z2[1]), .A2(n5209), .B1(n5171), .B2(
        wb_dsize_reg_z2[25]), .ZN(n4945) );
  NAND2_X2 U5485 ( .A1(n5209), .A2(wb_dsize_reg_z2[31]), .ZN(n4949) );
  NAND2_X2 U5486 ( .A1(reg31Val_0[31]), .A2(n4740), .ZN(n4948) );
  NAND2_X2 U5487 ( .A1(n4080), .A2(n4474), .ZN(n4952) );
  NAND2_X2 U5488 ( .A1(n6078), .A2(memAddr[31]), .ZN(n4951) );
  NAND2_X2 U5489 ( .A1(n4748), .A2(regWrData[31]), .ZN(n4950) );
  NAND2_X2 U5490 ( .A1(n7379), .A2(n4121), .ZN(n8333) );
  NAND2_X2 U5491 ( .A1(n4743), .A2(n4625), .ZN(n4954) );
  NAND2_X2 U5492 ( .A1(n5209), .A2(wb_dsize_reg_z2[29]), .ZN(n4953) );
  INV_X4 U5493 ( .A(regWrData[29]), .ZN(n4958) );
  OAI221_X2 U5494 ( .B1(n4732), .B2(n9045), .C1(n4958), .C2(n4733), .A(n4957), 
        .ZN(n8335) );
  NAND2_X2 U5495 ( .A1(n4743), .A2(n4449), .ZN(n4960) );
  NAND2_X2 U5496 ( .A1(n4739), .A2(wb_dsize_reg_z2[28]), .ZN(n4959) );
  NAND2_X2 U5497 ( .A1(n4743), .A2(n4450), .ZN(n4962) );
  NAND2_X2 U5498 ( .A1(n5209), .A2(wb_dsize_reg_z2[26]), .ZN(n4961) );
  NAND2_X2 U5499 ( .A1(n5209), .A2(wb_dsize_reg_z2[20]), .ZN(n4964) );
  NAND2_X2 U5500 ( .A1(reg31Val_0[20]), .A2(n4740), .ZN(n4963) );
  NAND2_X2 U5501 ( .A1(n4102), .A2(regWrData[14]), .ZN(n4967) );
  NAND2_X2 U5502 ( .A1(n4101), .A2(memAddr[14]), .ZN(n4966) );
  INV_X4 U5503 ( .A(n8646), .ZN(n4965) );
  NAND2_X2 U5504 ( .A1(n5170), .A2(wb_dsize_reg_z2[22]), .ZN(n4970) );
  AOI22_X2 U5505 ( .A1(wb_dsize_reg_z2[6]), .A2(n5209), .B1(
        wb_dsize_reg_z2[30]), .B2(n5171), .ZN(n4969) );
  NAND2_X2 U5506 ( .A1(n4102), .A2(regWrData[6]), .ZN(n4976) );
  NAND2_X2 U5507 ( .A1(n4101), .A2(memAddr[6]), .ZN(n4975) );
  NAND2_X2 U5508 ( .A1(n5170), .A2(wb_dsize_reg_z2[21]), .ZN(n4979) );
  AOI22_X2 U5509 ( .A1(wb_dsize_reg_z2[5]), .A2(n5209), .B1(
        wb_dsize_reg_z2[29]), .B2(n5171), .ZN(n4978) );
  NAND2_X2 U5510 ( .A1(n4102), .A2(regWrData[5]), .ZN(n4985) );
  NAND2_X2 U5511 ( .A1(n4101), .A2(memAddr[5]), .ZN(n4984) );
  NAND2_X2 U5512 ( .A1(n5170), .A2(wb_dsize_reg_z2[23]), .ZN(n4988) );
  AOI22_X2 U5513 ( .A1(wb_dsize_reg_z2[7]), .A2(n5209), .B1(n5171), .B2(
        wb_dsize_reg_z2[31]), .ZN(n4987) );
  NAND2_X2 U5514 ( .A1(n4102), .A2(regWrData[7]), .ZN(n4994) );
  NAND2_X2 U5515 ( .A1(n4101), .A2(memAddr[7]), .ZN(n4993) );
  NAND2_X2 U5516 ( .A1(n4102), .A2(regWrData[13]), .ZN(n4999) );
  NAND2_X2 U5517 ( .A1(n4101), .A2(memAddr[13]), .ZN(n4998) );
  NAND2_X2 U5518 ( .A1(n4743), .A2(n4623), .ZN(n5001) );
  NAND2_X2 U5519 ( .A1(n4739), .A2(wb_dsize_reg_z2[30]), .ZN(n5000) );
  INV_X4 U5520 ( .A(regWrData[30]), .ZN(n5005) );
  OAI221_X2 U5521 ( .B1(n9049), .B2(n4732), .C1(n5005), .C2(n4733), .A(n5004), 
        .ZN(n8325) );
  NAND2_X2 U5522 ( .A1(n5170), .A2(wb_dsize_reg_z2[31]), .ZN(n5009) );
  OAI211_X2 U5523 ( .C1(n5029), .C2(n4637), .A(n5009), .B(n5008), .ZN(
        regWrData[15]) );
  NAND2_X2 U5524 ( .A1(n4102), .A2(regWrData[15]), .ZN(n5014) );
  NAND2_X2 U5525 ( .A1(n4101), .A2(memAddr[15]), .ZN(n5013) );
  AOI22_X2 U5526 ( .A1(n4707), .A2(n4079), .B1(n4413), .B2(n4452), .ZN(n5017)
         );
  NAND2_X2 U5527 ( .A1(n4101), .A2(memAddr[12]), .ZN(n5016) );
  NAND2_X2 U5528 ( .A1(n4102), .A2(regWrData[12]), .ZN(n5015) );
  AOI22_X2 U5529 ( .A1(n4715), .A2(n4079), .B1(n4414), .B2(n4452), .ZN(n5020)
         );
  NAND2_X2 U5530 ( .A1(n4101), .A2(memAddr[11]), .ZN(n5019) );
  NAND2_X2 U5531 ( .A1(n4102), .A2(regWrData[11]), .ZN(n5018) );
  NAND2_X2 U5532 ( .A1(n5170), .A2(wb_dsize_reg_z2[25]), .ZN(n5024) );
  OAI211_X2 U5533 ( .C1(n5029), .C2(n4635), .A(n5024), .B(n5023), .ZN(
        regWrData[9]) );
  NAND2_X2 U5534 ( .A1(n5170), .A2(wb_dsize_reg_z2[24]), .ZN(n5028) );
  OAI211_X2 U5535 ( .C1(n5029), .C2(n4636), .A(n5028), .B(n5027), .ZN(
        regWrData[8]) );
  NAND2_X2 U5536 ( .A1(n4743), .A2(n4626), .ZN(n5031) );
  NAND2_X2 U5537 ( .A1(n4739), .A2(wb_dsize_reg_z2[27]), .ZN(n5030) );
  NAND2_X2 U5538 ( .A1(n4739), .A2(wb_dsize_reg_z2[21]), .ZN(n5033) );
  NAND2_X2 U5539 ( .A1(reg31Val_0[21]), .A2(n4740), .ZN(n5032) );
  NAND2_X2 U5540 ( .A1(n4739), .A2(wb_dsize_reg_z2[19]), .ZN(n5035) );
  NAND2_X2 U5541 ( .A1(reg31Val_0[19]), .A2(n4740), .ZN(n5034) );
  INV_X4 U5542 ( .A(regWrData[19]), .ZN(n5038) );
  OAI221_X2 U5543 ( .B1(n9022), .B2(n4732), .C1(n5038), .C2(n4733), .A(n5037), 
        .ZN(n6275) );
  INV_X4 U5544 ( .A(regWrData[21]), .ZN(n5041) );
  OAI221_X2 U5545 ( .B1(n9026), .B2(n4732), .C1(n5041), .C2(n4733), .A(n5040), 
        .ZN(n6273) );
  INV_X4 U5546 ( .A(regWrData[27]), .ZN(n5044) );
  OAI221_X2 U5547 ( .B1(n9041), .B2(n4732), .C1(n5044), .C2(n4733), .A(n5043), 
        .ZN(n6267) );
  INV_X4 U5548 ( .A(n7906), .ZN(n7537) );
  INV_X4 U5549 ( .A(n7682), .ZN(n7536) );
  NAND2_X2 U5550 ( .A1(n4102), .A2(regWrData[9]), .ZN(n5049) );
  NAND2_X2 U5551 ( .A1(n4101), .A2(memAddr[9]), .ZN(n5048) );
  INV_X4 U5552 ( .A(n5267), .ZN(n6320) );
  NAND2_X2 U5553 ( .A1(n4102), .A2(regWrData[8]), .ZN(n5054) );
  NAND2_X2 U5554 ( .A1(n4101), .A2(memAddr[8]), .ZN(n5053) );
  AOI22_X2 U5555 ( .A1(n4704), .A2(n4079), .B1(n4415), .B2(n4452), .ZN(n5057)
         );
  NAND2_X2 U5556 ( .A1(n4101), .A2(memAddr[10]), .ZN(n5056) );
  NAND2_X2 U5557 ( .A1(n4102), .A2(regWrData[10]), .ZN(n5055) );
  INV_X4 U5558 ( .A(regWrData[20]), .ZN(n5062) );
  OAI221_X2 U5559 ( .B1(n9024), .B2(n4732), .C1(n5062), .C2(n4733), .A(n5061), 
        .ZN(n6274) );
  INV_X4 U5560 ( .A(n7977), .ZN(n7540) );
  INV_X4 U5561 ( .A(regWrData[26]), .ZN(n5066) );
  OAI221_X2 U5562 ( .B1(n9039), .B2(n4732), .C1(n5066), .C2(n4733), .A(n5065), 
        .ZN(n6268) );
  INV_X4 U5563 ( .A(regWrData[28]), .ZN(n5070) );
  OAI221_X2 U5564 ( .B1(n4732), .B2(n9043), .C1(n5070), .C2(n4733), .A(n5069), 
        .ZN(n6266) );
  INV_X4 U5565 ( .A(n8325), .ZN(n5074) );
  INV_X4 U5566 ( .A(n8479), .ZN(n5073) );
  NAND2_X2 U5567 ( .A1(n5074), .A2(n5073), .ZN(n5076) );
  INV_X4 U5568 ( .A(n7968), .ZN(n7539) );
  INV_X4 U5569 ( .A(n7671), .ZN(n7538) );
  INV_X4 U5570 ( .A(n7696), .ZN(n5663) );
  NAND4_X2 U5571 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), .ZN(n5082)
         );
  INV_X4 U5572 ( .A(n8333), .ZN(n7546) );
  INV_X4 U5573 ( .A(n5082), .ZN(n5083) );
  NAND2_X2 U5574 ( .A1(n5083), .A2(n4136), .ZN(n8493) );
  NAND2_X2 U5575 ( .A1(n5083), .A2(n9051), .ZN(n8492) );
  NAND2_X2 U5576 ( .A1(n4739), .A2(wb_dsize_reg_z2[22]), .ZN(n5085) );
  NAND2_X2 U5577 ( .A1(reg31Val_0[22]), .A2(n4740), .ZN(n5084) );
  NAND2_X2 U5578 ( .A1(n6078), .A2(memAddr[22]), .ZN(n5087) );
  NAND2_X2 U5579 ( .A1(n4748), .A2(regWrData[22]), .ZN(n5086) );
  NAND2_X2 U5580 ( .A1(n4746), .A2(memAddr[9]), .ZN(n5089) );
  NAND2_X2 U5581 ( .A1(regWrData[9]), .A2(n4748), .ZN(n5088) );
  NAND2_X2 U5582 ( .A1(n6365), .A2(n7531), .ZN(n5091) );
  NAND2_X2 U5583 ( .A1(n8364), .A2(n7530), .ZN(n5090) );
  NAND2_X2 U5584 ( .A1(n6078), .A2(memAddr[30]), .ZN(n5094) );
  NAND2_X2 U5585 ( .A1(n4712), .A2(n4080), .ZN(n5093) );
  NAND2_X2 U5586 ( .A1(n4748), .A2(regWrData[30]), .ZN(n5092) );
  NAND2_X2 U5587 ( .A1(n4080), .A2(n4371), .ZN(n5097) );
  NAND2_X2 U5588 ( .A1(n4746), .A2(memAddr[1]), .ZN(n5096) );
  NAND2_X2 U5589 ( .A1(regWrData[1]), .A2(n4748), .ZN(n5095) );
  NAND2_X2 U5590 ( .A1(n7212), .A2(n7531), .ZN(n5099) );
  NAND2_X2 U5591 ( .A1(n8306), .A2(n7530), .ZN(n5098) );
  INV_X4 U5592 ( .A(n8474), .ZN(n7564) );
  AOI221_X2 U5593 ( .B1(n8381), .B2(n8391), .C1(n8452), .C2(n7558), .A(n7564), 
        .ZN(n6277) );
  NAND2_X2 U5594 ( .A1(n4102), .A2(regWrData[2]), .ZN(n5104) );
  NAND2_X2 U5595 ( .A1(n4101), .A2(memAddr[2]), .ZN(n5103) );
  INV_X4 U5596 ( .A(n5935), .ZN(n7548) );
  NAND2_X2 U5597 ( .A1(n4102), .A2(regWrData[1]), .ZN(n5109) );
  NAND2_X2 U5598 ( .A1(n4101), .A2(memAddr[1]), .ZN(n5108) );
  INV_X4 U5599 ( .A(n7211), .ZN(n5925) );
  NAND2_X2 U5600 ( .A1(n5115), .A2(n5114), .ZN(n7706) );
  NAND2_X2 U5601 ( .A1(n4739), .A2(wb_dsize_reg_z2[23]), .ZN(n5117) );
  NAND2_X2 U5602 ( .A1(reg31Val_0[23]), .A2(n4741), .ZN(n5116) );
  NAND2_X2 U5603 ( .A1(n4746), .A2(memAddr[23]), .ZN(n5119) );
  NAND2_X2 U5604 ( .A1(n4748), .A2(regWrData[23]), .ZN(n5118) );
  NAND2_X2 U5605 ( .A1(n4746), .A2(memAddr[8]), .ZN(n5121) );
  NAND2_X2 U5606 ( .A1(regWrData[8]), .A2(n6079), .ZN(n5120) );
  NAND2_X2 U5607 ( .A1(n4737), .A2(n7531), .ZN(n5123) );
  NAND2_X2 U5608 ( .A1(n8326), .A2(n7530), .ZN(n5122) );
  NAND2_X2 U5609 ( .A1(n4080), .A2(n4372), .ZN(n5126) );
  NAND2_X2 U5610 ( .A1(n4746), .A2(memAddr[0]), .ZN(n5125) );
  NAND2_X2 U5611 ( .A1(regWrData[0]), .A2(n6079), .ZN(n5124) );
  NAND2_X2 U5612 ( .A1(n7479), .A2(n7531), .ZN(n5128) );
  NAND2_X2 U5613 ( .A1(n7379), .A2(n7530), .ZN(n5127) );
  NAND2_X2 U5614 ( .A1(n5170), .A2(wb_dsize_reg_z2[19]), .ZN(n5131) );
  AOI22_X2 U5615 ( .A1(wb_dsize_reg_z2[3]), .A2(n5209), .B1(
        wb_dsize_reg_z2[27]), .B2(n5171), .ZN(n5130) );
  NAND2_X2 U5616 ( .A1(n4102), .A2(regWrData[3]), .ZN(n5137) );
  NAND2_X2 U5617 ( .A1(n4101), .A2(memAddr[3]), .ZN(n5136) );
  AOI221_X2 U5618 ( .B1(n8451), .B2(n7525), .C1(n8452), .C2(n8391), .A(n8392), 
        .ZN(n5644) );
  AOI221_X2 U5619 ( .B1(n8431), .B2(n7525), .C1(n8432), .C2(n8391), .A(n8392), 
        .ZN(n5946) );
  INV_X4 U5620 ( .A(n8409), .ZN(n5140) );
  INV_X4 U5621 ( .A(n5944), .ZN(n5141) );
  AOI22_X2 U5622 ( .A1(n6254), .A2(n5141), .B1(n8404), .B2(n6258), .ZN(n5142)
         );
  NAND2_X2 U5623 ( .A1(n5143), .A2(n5142), .ZN(n7709) );
  INV_X4 U5624 ( .A(n8392), .ZN(n5445) );
  OAI211_X2 U5625 ( .C1(n8440), .C2(n8019), .A(n8441), .B(n5445), .ZN(n5660)
         );
  NAND2_X2 U5626 ( .A1(n4735), .A2(n5660), .ZN(n5147) );
  INV_X4 U5627 ( .A(n8391), .ZN(n7563) );
  OAI211_X2 U5628 ( .C1(n8417), .C2(n8019), .A(n5445), .B(n4499), .ZN(n5825)
         );
  NAND2_X2 U5629 ( .A1(n6254), .A2(n5825), .ZN(n5146) );
  OAI211_X2 U5630 ( .C1(n8470), .C2(n8019), .A(n8471), .B(n5445), .ZN(n5800)
         );
  NAND3_X2 U5631 ( .A1(n5147), .A2(n5146), .A3(n5145), .ZN(n7686) );
  INV_X4 U5632 ( .A(n7706), .ZN(n8401) );
  NAND2_X2 U5633 ( .A1(n4102), .A2(regWrData[0]), .ZN(n5152) );
  NAND2_X2 U5634 ( .A1(n4101), .A2(memAddr[0]), .ZN(n5151) );
  NAND3_X4 U5635 ( .A1(n5152), .A2(n5151), .A3(n5150), .ZN(n7422) );
  INV_X4 U5636 ( .A(n7422), .ZN(n7430) );
  OAI22_X2 U5637 ( .A1(n8393), .A2(n4128), .B1(n8371), .B2(n4734), .ZN(n5159)
         );
  NAND2_X2 U5638 ( .A1(n8473), .A2(n8391), .ZN(n5155) );
  NAND2_X2 U5639 ( .A1(n5156), .A2(n5155), .ZN(n5806) );
  INV_X4 U5640 ( .A(n5806), .ZN(n5651) );
  INV_X4 U5641 ( .A(n7526), .ZN(n5160) );
  NAND2_X2 U5642 ( .A1(n4076), .A2(n5160), .ZN(n5163) );
  NAND2_X2 U5643 ( .A1(n7707), .A2(n7648), .ZN(n5162) );
  NAND2_X2 U5644 ( .A1(n8475), .A2(n7422), .ZN(n5978) );
  NAND2_X2 U5645 ( .A1(n7430), .A2(n8475), .ZN(n5975) );
  AOI22_X2 U5646 ( .A1(n7209), .A2(n7686), .B1(n7219), .B2(n7709), .ZN(n5161)
         );
  NAND4_X2 U5647 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n7647)
         );
  NAND2_X2 U5648 ( .A1(n6254), .A2(n5806), .ZN(n5168) );
  NAND2_X2 U5649 ( .A1(n5170), .A2(wb_dsize_reg_z2[20]), .ZN(n5173) );
  AOI22_X2 U5650 ( .A1(wb_dsize_reg_z2[4]), .A2(n5209), .B1(
        wb_dsize_reg_z2[28]), .B2(n5171), .ZN(n5172) );
  AOI22_X2 U5651 ( .A1(n4713), .A2(n4079), .B1(n4370), .B2(n4452), .ZN(n5177)
         );
  NAND2_X2 U5652 ( .A1(n4101), .A2(memAddr[4]), .ZN(n5176) );
  NAND2_X2 U5653 ( .A1(n4102), .A2(regWrData[4]), .ZN(n5175) );
  INV_X4 U5654 ( .A(n7918), .ZN(n7524) );
  NAND2_X2 U5655 ( .A1(n7530), .A2(n7524), .ZN(n8489) );
  NAND2_X2 U5656 ( .A1(n6258), .A2(n5800), .ZN(n5186) );
  INV_X4 U5657 ( .A(n8390), .ZN(n5182) );
  NAND2_X2 U5658 ( .A1(n8445), .A2(n7918), .ZN(n5180) );
  INV_X4 U5659 ( .A(n8489), .ZN(n7523) );
  NAND2_X2 U5660 ( .A1(n6365), .A2(n7523), .ZN(n5179) );
  NAND3_X2 U5661 ( .A1(n5180), .A2(n5179), .A3(n5178), .ZN(n6251) );
  INV_X4 U5662 ( .A(n6251), .ZN(n5181) );
  OAI221_X2 U5663 ( .B1(n7563), .B2(n5182), .C1(n8019), .C2(n5181), .A(n5445), 
        .ZN(n5930) );
  NAND2_X2 U5664 ( .A1(n6254), .A2(n5930), .ZN(n5185) );
  NAND2_X2 U5665 ( .A1(n4312), .A2(n5660), .ZN(n5184) );
  NAND2_X2 U5666 ( .A1(n4735), .A2(n5825), .ZN(n5183) );
  NAND4_X2 U5667 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n7887)
         );
  NAND2_X2 U5668 ( .A1(n7219), .A2(n7887), .ZN(n5194) );
  NAND2_X2 U5669 ( .A1(n7209), .A2(n7709), .ZN(n5193) );
  INV_X4 U5670 ( .A(n7216), .ZN(n7427) );
  INV_X4 U5671 ( .A(n6365), .ZN(n7192) );
  MUX2_X2 U5672 ( .A(n4731), .B(n4077), .S(n7192), .Z(n5187) );
  NAND2_X2 U5673 ( .A1(n5188), .A2(n6365), .ZN(n5189) );
  NAND2_X2 U5674 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  NAND4_X2 U5675 ( .A1(n5194), .A2(n4523), .A3(n5193), .A4(n5192), .ZN(n7089)
         );
  MUX2_X2 U5676 ( .A(n6365), .B(n7089), .S(n4091), .Z(n7653) );
  NAND2_X2 U5677 ( .A1(n4739), .A2(wb_dsize_reg_z2[24]), .ZN(n5196) );
  NAND2_X2 U5678 ( .A1(reg31Val_0[24]), .A2(n4741), .ZN(n5195) );
  NAND2_X2 U5679 ( .A1(n4739), .A2(wb_dsize_reg_z2[16]), .ZN(n5198) );
  NAND2_X2 U5680 ( .A1(reg31Val_0[16]), .A2(n4741), .ZN(n5197) );
  INV_X4 U5681 ( .A(regWrData[16]), .ZN(n5202) );
  OAI221_X2 U5682 ( .B1(n9016), .B2(n4732), .C1(n5202), .C2(n4733), .A(n5201), 
        .ZN(n8458) );
  NAND2_X2 U5683 ( .A1(n4746), .A2(memAddr[2]), .ZN(n5204) );
  NAND2_X2 U5684 ( .A1(regWrData[2]), .A2(n6079), .ZN(n5203) );
  NAND2_X2 U5685 ( .A1(n4739), .A2(wb_dsize_reg_z2[18]), .ZN(n5206) );
  NAND2_X2 U5686 ( .A1(reg31Val_0[18]), .A2(n4741), .ZN(n5205) );
  NAND2_X2 U5687 ( .A1(n4739), .A2(wb_dsize_reg_z2[17]), .ZN(n5208) );
  NAND2_X2 U5688 ( .A1(reg31Val_0[17]), .A2(n4741), .ZN(n5207) );
  NAND2_X2 U5689 ( .A1(n4739), .A2(wb_dsize_reg_z2[25]), .ZN(n5213) );
  NAND2_X2 U5690 ( .A1(reg31Val_0[25]), .A2(n4741), .ZN(n5212) );
  NAND2_X2 U5691 ( .A1(n4746), .A2(memAddr[3]), .ZN(n5215) );
  NAND2_X2 U5692 ( .A1(regWrData[3]), .A2(n6079), .ZN(n5214) );
  NAND2_X2 U5693 ( .A1(n4746), .A2(memAddr[4]), .ZN(n5217) );
  NAND2_X2 U5694 ( .A1(regWrData[4]), .A2(n6079), .ZN(n5216) );
  NAND2_X2 U5695 ( .A1(n4746), .A2(memAddr[5]), .ZN(n5219) );
  NAND2_X2 U5696 ( .A1(regWrData[5]), .A2(n6079), .ZN(n5218) );
  NAND2_X2 U5697 ( .A1(n4746), .A2(memAddr[6]), .ZN(n5221) );
  NAND2_X2 U5698 ( .A1(regWrData[6]), .A2(n6079), .ZN(n5220) );
  NAND2_X2 U5699 ( .A1(n4080), .A2(n4206), .ZN(n5224) );
  NAND2_X2 U5700 ( .A1(n4746), .A2(memAddr[7]), .ZN(n5223) );
  NAND2_X2 U5701 ( .A1(regWrData[7]), .A2(n6079), .ZN(n5222) );
  INV_X4 U5702 ( .A(n6071), .ZN(n5481) );
  NAND2_X2 U5703 ( .A1(n5481), .A2(n4135), .ZN(n5231) );
  INV_X4 U5704 ( .A(n5231), .ZN(n5225) );
  NAND2_X2 U5705 ( .A1(n5481), .A2(n4537), .ZN(n5226) );
  NAND2_X2 U5706 ( .A1(n7273), .A2(n6322), .ZN(n5235) );
  INV_X4 U5707 ( .A(n5226), .ZN(n5232) );
  NAND2_X2 U5708 ( .A1(n4078), .A2(n7422), .ZN(n5234) );
  NAND2_X2 U5709 ( .A1(n5231), .A2(n5226), .ZN(n7241) );
  INV_X4 U5710 ( .A(regWrData[24]), .ZN(n5230) );
  OAI221_X2 U5711 ( .B1(n9034), .B2(n4732), .C1(n5230), .C2(n4733), .A(n5229), 
        .ZN(n6270) );
  NAND2_X2 U5712 ( .A1(n5232), .A2(n5231), .ZN(n7362) );
  AOI22_X2 U5713 ( .A1(n7361), .A2(n6270), .B1(n7243), .B2(n8458), .ZN(n5233)
         );
  NAND2_X2 U5714 ( .A1(n4753), .A2(n7479), .ZN(n6897) );
  NAND2_X2 U5715 ( .A1(n7273), .A2(n8479), .ZN(n5245) );
  NAND2_X2 U5716 ( .A1(n4078), .A2(n7671), .ZN(n5244) );
  INV_X4 U5717 ( .A(regWrData[23]), .ZN(n5238) );
  OAI221_X2 U5718 ( .B1(n9031), .B2(n4732), .C1(n5238), .C2(n4733), .A(n5237), 
        .ZN(n6271) );
  INV_X4 U5719 ( .A(regWrData[31]), .ZN(n5242) );
  OAI221_X2 U5720 ( .B1(n8988), .B2(n4732), .C1(n5242), .C2(n4733), .A(n5241), 
        .ZN(n7381) );
  AOI22_X2 U5721 ( .A1(n7243), .A2(n6271), .B1(n7361), .B2(n7381), .ZN(n5243)
         );
  NAND2_X2 U5722 ( .A1(n7273), .A2(n7988), .ZN(n5251) );
  NAND2_X2 U5723 ( .A1(n4078), .A2(n7977), .ZN(n5250) );
  INV_X4 U5724 ( .A(regWrData[22]), .ZN(n5248) );
  OAI221_X2 U5725 ( .B1(n9028), .B2(n4732), .C1(n5248), .C2(n4733), .A(n5247), 
        .ZN(n6272) );
  AOI22_X2 U5726 ( .A1(n7243), .A2(n6272), .B1(n7361), .B2(n8325), .ZN(n5249)
         );
  NAND2_X2 U5727 ( .A1(n4108), .A2(n7479), .ZN(n5968) );
  INV_X4 U5728 ( .A(n5968), .ZN(n5364) );
  NAND2_X2 U5729 ( .A1(n7273), .A2(n7696), .ZN(n5254) );
  NAND2_X2 U5730 ( .A1(n4078), .A2(n7968), .ZN(n5253) );
  AOI22_X2 U5731 ( .A1(n7243), .A2(n6273), .B1(n7361), .B2(n8335), .ZN(n5252)
         );
  NAND2_X2 U5732 ( .A1(n7273), .A2(n7906), .ZN(n5257) );
  NAND2_X2 U5733 ( .A1(n4078), .A2(n7918), .ZN(n5256) );
  AOI22_X2 U5734 ( .A1(n7243), .A2(n6274), .B1(n7361), .B2(n6266), .ZN(n5255)
         );
  NAND2_X2 U5735 ( .A1(n4085), .A2(n7479), .ZN(n5667) );
  INV_X4 U5736 ( .A(n5667), .ZN(n5310) );
  NAND2_X2 U5737 ( .A1(n7273), .A2(n7682), .ZN(n5260) );
  NAND2_X2 U5738 ( .A1(n4078), .A2(n8019), .ZN(n5259) );
  AOI22_X2 U5739 ( .A1(n7243), .A2(n6275), .B1(n7361), .B2(n6267), .ZN(n5258)
         );
  INV_X4 U5740 ( .A(regWrData[18]), .ZN(n5263) );
  OAI221_X2 U5741 ( .B1(n9020), .B2(n4732), .C1(n5263), .C2(n4733), .A(n5262), 
        .ZN(n6276) );
  AOI22_X2 U5742 ( .A1(n7361), .A2(n6268), .B1(n7243), .B2(n6276), .ZN(n5266)
         );
  NAND2_X2 U5743 ( .A1(n4078), .A2(n5935), .ZN(n5265) );
  NAND2_X2 U5744 ( .A1(n7273), .A2(n5767), .ZN(n5264) );
  NAND2_X2 U5745 ( .A1(n4099), .A2(n7212), .ZN(n5286) );
  NAND2_X2 U5746 ( .A1(n7273), .A2(n5267), .ZN(n5278) );
  NAND2_X2 U5747 ( .A1(n4078), .A2(n7211), .ZN(n5277) );
  INV_X4 U5748 ( .A(regWrData[17]), .ZN(n5271) );
  OAI221_X2 U5749 ( .B1(n9018), .B2(n4732), .C1(n5271), .C2(n4733), .A(n5270), 
        .ZN(n5805) );
  INV_X4 U5750 ( .A(regWrData[25]), .ZN(n5275) );
  OAI221_X2 U5751 ( .B1(n9037), .B2(n4732), .C1(n5275), .C2(n4733), .A(n5274), 
        .ZN(n6269) );
  AOI22_X2 U5752 ( .A1(n7243), .A2(n5805), .B1(n7361), .B2(n6269), .ZN(n5276)
         );
  NAND2_X2 U5753 ( .A1(n4750), .A2(n7665), .ZN(n5296) );
  INV_X4 U5754 ( .A(n5296), .ZN(n5279) );
  NAND2_X2 U5755 ( .A1(n7663), .A2(n6157), .ZN(n5297) );
  INV_X4 U5756 ( .A(n5297), .ZN(n5299) );
  XNOR2_X2 U5757 ( .A(n5279), .B(n5299), .ZN(n5282) );
  NAND2_X2 U5758 ( .A1(n4753), .A2(n7212), .ZN(n5586) );
  INV_X4 U5759 ( .A(n5586), .ZN(n5280) );
  INV_X4 U5760 ( .A(n7479), .ZN(n7423) );
  INV_X4 U5761 ( .A(n7665), .ZN(n7520) );
  NAND2_X2 U5762 ( .A1(n7423), .A2(n7520), .ZN(n5796) );
  NAND2_X2 U5763 ( .A1(n5282), .A2(n5281), .ZN(n5285) );
  INV_X4 U5764 ( .A(n5281), .ZN(n5284) );
  INV_X4 U5765 ( .A(n5282), .ZN(n5283) );
  NAND2_X2 U5766 ( .A1(n5284), .A2(n5283), .ZN(n5295) );
  NAND2_X2 U5767 ( .A1(n5285), .A2(n5295), .ZN(n5287) );
  NAND2_X2 U5768 ( .A1(n5286), .A2(n5287), .ZN(n5289) );
  INV_X4 U5769 ( .A(n5287), .ZN(n5288) );
  NAND2_X2 U5770 ( .A1(n5289), .A2(n5294), .ZN(n5306) );
  NAND2_X2 U5771 ( .A1(n4099), .A2(n7479), .ZN(n5493) );
  INV_X4 U5772 ( .A(n5493), .ZN(n5293) );
  NAND2_X2 U5773 ( .A1(n7665), .A2(n4753), .ZN(n5291) );
  NAND3_X2 U5774 ( .A1(n6897), .A2(n7212), .A3(n4750), .ZN(n5290) );
  XNOR2_X2 U5775 ( .A(n5291), .B(n5290), .ZN(n5494) );
  INV_X4 U5776 ( .A(n5494), .ZN(n5292) );
  NAND2_X2 U5777 ( .A1(n5293), .A2(n5292), .ZN(n5495) );
  INV_X4 U5778 ( .A(n5298), .ZN(n5321) );
  NAND2_X2 U5779 ( .A1(n4754), .A2(n4752), .ZN(n5702) );
  INV_X4 U5780 ( .A(n5320), .ZN(n5303) );
  XNOR2_X2 U5781 ( .A(n5321), .B(n5303), .ZN(n5304) );
  NAND2_X2 U5782 ( .A1(n4142), .A2(n5304), .ZN(n5315) );
  XNOR2_X2 U5783 ( .A(n5314), .B(n5316), .ZN(n5305) );
  NAND2_X2 U5784 ( .A1(n4159), .A2(n5305), .ZN(n5311) );
  NAND2_X2 U5785 ( .A1(n4084), .A2(n7479), .ZN(n5598) );
  INV_X4 U5786 ( .A(n5598), .ZN(n5308) );
  XNOR2_X2 U5787 ( .A(n5306), .B(n5495), .ZN(n5599) );
  INV_X4 U5788 ( .A(n5599), .ZN(n5307) );
  NAND2_X2 U5789 ( .A1(n5308), .A2(n5307), .ZN(n5312) );
  XNOR2_X2 U5790 ( .A(n5313), .B(n5312), .ZN(n5668) );
  INV_X4 U5791 ( .A(n5668), .ZN(n5309) );
  NAND2_X2 U5792 ( .A1(n5310), .A2(n5309), .ZN(n5669) );
  INV_X4 U5793 ( .A(n5314), .ZN(n5317) );
  INV_X4 U5794 ( .A(n5318), .ZN(n5337) );
  OAI21_X4 U5795 ( .B1(n5321), .B2(n5320), .A(n5319), .ZN(n5339) );
  NAND2_X2 U5796 ( .A1(n7659), .A2(n4753), .ZN(n5322) );
  INV_X4 U5797 ( .A(n5322), .ZN(n5344) );
  INV_X4 U5798 ( .A(n7661), .ZN(n7515) );
  NAND2_X2 U5799 ( .A1(n5340), .A2(n5323), .ZN(n5341) );
  XNOR2_X2 U5800 ( .A(n5339), .B(n5341), .ZN(n5324) );
  NAND2_X2 U5801 ( .A1(n4150), .A2(n5324), .ZN(n5335) );
  INV_X4 U5802 ( .A(n5336), .ZN(n5325) );
  XNOR2_X2 U5803 ( .A(n5337), .B(n5325), .ZN(n5326) );
  NAND2_X2 U5804 ( .A1(n4165), .A2(n5326), .ZN(n5331) );
  XNOR2_X2 U5805 ( .A(n5330), .B(n5332), .ZN(n5327) );
  NAND2_X2 U5806 ( .A1(n4160), .A2(n5327), .ZN(n5328) );
  INV_X4 U5807 ( .A(n5329), .ZN(n5386) );
  INV_X4 U5808 ( .A(n5330), .ZN(n5333) );
  INV_X4 U5809 ( .A(n5334), .ZN(n5370) );
  INV_X4 U5810 ( .A(n5338), .ZN(n5373) );
  INV_X4 U5811 ( .A(n5339), .ZN(n5342) );
  OAI21_X4 U5812 ( .B1(n5342), .B2(n5341), .A(n5340), .ZN(n5343) );
  INV_X4 U5813 ( .A(n5343), .ZN(n5377) );
  INV_X4 U5814 ( .A(n7659), .ZN(n7514) );
  NAND2_X2 U5815 ( .A1(n4754), .A2(n7514), .ZN(n5347) );
  INV_X4 U5816 ( .A(n5376), .ZN(n5348) );
  XNOR2_X2 U5817 ( .A(n5377), .B(n5348), .ZN(n5349) );
  NAND2_X2 U5818 ( .A1(n4103), .A2(n5349), .ZN(n5371) );
  INV_X4 U5819 ( .A(n5372), .ZN(n5350) );
  XNOR2_X2 U5820 ( .A(n5373), .B(n5350), .ZN(n5351) );
  NAND2_X2 U5821 ( .A1(n4163), .A2(n5351), .ZN(n5368) );
  INV_X4 U5822 ( .A(n5369), .ZN(n5352) );
  XNOR2_X2 U5823 ( .A(n5370), .B(n5352), .ZN(n5353) );
  NAND2_X2 U5824 ( .A1(n4158), .A2(n5353), .ZN(n5384) );
  INV_X4 U5825 ( .A(n5385), .ZN(n5354) );
  XNOR2_X2 U5826 ( .A(n5386), .B(n5354), .ZN(n5355) );
  NAND2_X2 U5827 ( .A1(n4191), .A2(n5355), .ZN(n5365) );
  INV_X4 U5828 ( .A(n5366), .ZN(n5362) );
  NAND2_X2 U5829 ( .A1(n4100), .A2(n7479), .ZN(n5722) );
  INV_X4 U5830 ( .A(n5722), .ZN(n5360) );
  INV_X4 U5831 ( .A(n5356), .ZN(n5358) );
  INV_X4 U5832 ( .A(n5669), .ZN(n5357) );
  XNOR2_X2 U5833 ( .A(n5358), .B(n5357), .ZN(n5723) );
  INV_X4 U5834 ( .A(n5723), .ZN(n5359) );
  NAND2_X2 U5835 ( .A1(n5360), .A2(n5359), .ZN(n5367) );
  INV_X4 U5836 ( .A(n5367), .ZN(n5361) );
  XNOR2_X2 U5837 ( .A(n5362), .B(n5361), .ZN(n5969) );
  INV_X4 U5838 ( .A(n5969), .ZN(n5363) );
  NAND2_X2 U5839 ( .A1(n5364), .A2(n5363), .ZN(n5970) );
  INV_X4 U5840 ( .A(n5398), .ZN(n5388) );
  INV_X4 U5841 ( .A(n5374), .ZN(n5412) );
  NAND2_X2 U5842 ( .A1(n7617), .A2(n4753), .ZN(n5378) );
  INV_X4 U5843 ( .A(n5378), .ZN(n5419) );
  INV_X4 U5844 ( .A(n7657), .ZN(n7513) );
  NAND2_X2 U5845 ( .A1(n5415), .A2(n5379), .ZN(n5416) );
  XNOR2_X2 U5846 ( .A(n5414), .B(n5416), .ZN(n5380) );
  NAND2_X2 U5847 ( .A1(n4151), .A2(n5380), .ZN(n5410) );
  INV_X4 U5848 ( .A(n5411), .ZN(n5381) );
  XNOR2_X2 U5849 ( .A(n5412), .B(n5381), .ZN(n5382) );
  NAND2_X2 U5850 ( .A1(n4167), .A2(n5382), .ZN(n5406) );
  XNOR2_X2 U5851 ( .A(n5405), .B(n5407), .ZN(n5383) );
  NAND2_X2 U5852 ( .A1(n4157), .A2(n5383), .ZN(n5401) );
  XNOR2_X2 U5853 ( .A(n5402), .B(n5400), .ZN(n5396) );
  NAND2_X2 U5854 ( .A1(n7665), .A2(n4100), .ZN(n5395) );
  XNOR2_X2 U5855 ( .A(n5396), .B(n5395), .ZN(n5399) );
  INV_X4 U5856 ( .A(n5399), .ZN(n5387) );
  XNOR2_X2 U5857 ( .A(n5388), .B(n5387), .ZN(n5390) );
  NAND2_X2 U5858 ( .A1(n4108), .A2(n7212), .ZN(n5389) );
  NAND2_X2 U5859 ( .A1(n5390), .A2(n5389), .ZN(n5392) );
  INV_X4 U5860 ( .A(n5390), .ZN(n5391) );
  NAND2_X2 U5861 ( .A1(n5392), .A2(n5393), .ZN(n5434) );
  INV_X4 U5862 ( .A(n5394), .ZN(n5503) );
  INV_X4 U5863 ( .A(n5395), .ZN(n5397) );
  AOI22_X2 U5864 ( .A1(n5399), .A2(n5398), .B1(n5397), .B2(n5396), .ZN(n5507)
         );
  INV_X4 U5865 ( .A(n5400), .ZN(n5403) );
  INV_X4 U5866 ( .A(n5404), .ZN(n5511) );
  INV_X4 U5867 ( .A(n5405), .ZN(n5408) );
  INV_X4 U5868 ( .A(n5409), .ZN(n5515) );
  INV_X4 U5869 ( .A(n5413), .ZN(n5519) );
  INV_X4 U5870 ( .A(n5414), .ZN(n5417) );
  OAI21_X4 U5871 ( .B1(n5417), .B2(n5416), .A(n5415), .ZN(n5418) );
  INV_X4 U5872 ( .A(n5418), .ZN(n5526) );
  INV_X4 U5873 ( .A(n7617), .ZN(n7512) );
  NAND2_X2 U5874 ( .A1(n4754), .A2(n7512), .ZN(n5420) );
  NAND4_X2 U5875 ( .A1(n5421), .A2(n5702), .A3(n5524), .A4(n5420), .ZN(n5525)
         );
  INV_X4 U5876 ( .A(n5525), .ZN(n5422) );
  XNOR2_X2 U5877 ( .A(n5526), .B(n5422), .ZN(n5423) );
  NAND2_X2 U5878 ( .A1(n4143), .A2(n5423), .ZN(n5517) );
  INV_X4 U5879 ( .A(n5518), .ZN(n5424) );
  XNOR2_X2 U5880 ( .A(n5519), .B(n5424), .ZN(n5425) );
  NAND2_X2 U5881 ( .A1(n4164), .A2(n5425), .ZN(n5513) );
  INV_X4 U5882 ( .A(n5514), .ZN(n5426) );
  XNOR2_X2 U5883 ( .A(n5515), .B(n5426), .ZN(n5427) );
  NAND2_X2 U5884 ( .A1(n4269), .A2(n5427), .ZN(n5509) );
  INV_X4 U5885 ( .A(n5510), .ZN(n5428) );
  XNOR2_X2 U5886 ( .A(n5511), .B(n5428), .ZN(n5429) );
  NAND2_X2 U5887 ( .A1(n4216), .A2(n5429), .ZN(n5505) );
  INV_X4 U5888 ( .A(n5506), .ZN(n5430) );
  XNOR2_X2 U5889 ( .A(n5507), .B(n5430), .ZN(n5431) );
  NAND2_X2 U5890 ( .A1(n4197), .A2(n5431), .ZN(n5501) );
  INV_X4 U5891 ( .A(n5502), .ZN(n5432) );
  XNOR2_X2 U5892 ( .A(n5503), .B(n5432), .ZN(n5433) );
  NAND2_X2 U5893 ( .A1(n4254), .A2(n5433), .ZN(n5497) );
  INV_X4 U5894 ( .A(n5498), .ZN(n5438) );
  NAND2_X2 U5895 ( .A1(n7266), .A2(n7479), .ZN(n5477) );
  INV_X4 U5896 ( .A(n5477), .ZN(n5436) );
  XNOR2_X2 U5897 ( .A(n5970), .B(n5434), .ZN(n5478) );
  INV_X4 U5898 ( .A(n5478), .ZN(n5435) );
  NAND2_X2 U5899 ( .A1(n5436), .A2(n5435), .ZN(n5499) );
  INV_X4 U5900 ( .A(n5499), .ZN(n5437) );
  XNOR2_X2 U5901 ( .A(n5438), .B(n5437), .ZN(n6892) );
  OAI22_X2 U5902 ( .A1(n6897), .A2(n4169), .B1(n6892), .B2(n4784), .ZN(n5582)
         );
  INV_X4 U5903 ( .A(n5582), .ZN(n5439) );
  XNOR2_X2 U5904 ( .A(n5439), .B(n4479), .ZN(n7508) );
  OAI221_X2 U5905 ( .B1(n8362), .B2(n4736), .C1(n8379), .C2(n4317), .A(n5442), 
        .ZN(n7676) );
  NAND2_X2 U5906 ( .A1(n4468), .A2(n8326), .ZN(n5444) );
  OAI211_X2 U5907 ( .C1(n8447), .C2(n7524), .A(n5444), .B(n5443), .ZN(n7385)
         );
  NAND2_X2 U5908 ( .A1(n5452), .A2(n5451), .ZN(n7913) );
  INV_X4 U5909 ( .A(n7887), .ZN(n8389) );
  INV_X4 U5910 ( .A(n7888), .ZN(n7912) );
  AOI21_X2 U5911 ( .B1(n7219), .B2(n7913), .A(n5453), .ZN(n5460) );
  MUX2_X2 U5912 ( .A(n4731), .B(n4077), .S(n4088), .Z(n5454) );
  NAND2_X2 U5913 ( .A1(n5455), .A2(n4737), .ZN(n5456) );
  NAND2_X2 U5914 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  AOI21_X2 U5915 ( .B1(n7427), .B2(n7676), .A(n5458), .ZN(n5459) );
  OAI211_X2 U5916 ( .C1(n8389), .C2(n5978), .A(n5460), .B(n5459), .ZN(n6982)
         );
  MUX2_X2 U5917 ( .A(n4737), .B(n6982), .S(n4091), .Z(n7655) );
  OAI221_X2 U5918 ( .B1(n8393), .B2(n4736), .C1(n8371), .C2(n4317), .A(n5463), 
        .ZN(n7670) );
  NAND2_X2 U5919 ( .A1(n6258), .A2(n5660), .ZN(n5468) );
  NAND2_X2 U5920 ( .A1(n4312), .A2(n5825), .ZN(n5467) );
  OAI211_X2 U5921 ( .C1(n8470), .C2(n7525), .A(n8507), .B(n8506), .ZN(n6257)
         );
  INV_X4 U5922 ( .A(n5930), .ZN(n5464) );
  AOI21_X2 U5923 ( .B1(n6254), .B2(n6257), .A(n5465), .ZN(n5466) );
  NAND3_X2 U5924 ( .A1(n5468), .A2(n5467), .A3(n5466), .ZN(n7675) );
  INV_X4 U5925 ( .A(n7670), .ZN(n8370) );
  NAND2_X2 U5926 ( .A1(n4076), .A2(n7676), .ZN(n5473) );
  NAND2_X2 U5927 ( .A1(n7672), .A2(n7617), .ZN(n5472) );
  AOI22_X2 U5928 ( .A1(n7209), .A2(n7913), .B1(n7219), .B2(n7675), .ZN(n5471)
         );
  NAND4_X2 U5929 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n7474)
         );
  INV_X4 U5930 ( .A(n7474), .ZN(n5476) );
  NAND2_X2 U5931 ( .A1(n4791), .A2(n4091), .ZN(n5967) );
  OAI22_X2 U5932 ( .A1(n5476), .A2(n5967), .B1(n7982), .B2(n7616), .ZN(n5480)
         );
  XNOR2_X2 U5933 ( .A(n5478), .B(n5477), .ZN(n6286) );
  MUX2_X2 U5934 ( .A(n7574), .B(n6286), .S(n4078), .Z(n7475) );
  NAND2_X2 U5935 ( .A1(n4791), .A2(n4794), .ZN(n6046) );
  NAND2_X2 U5936 ( .A1(n4791), .A2(n4130), .ZN(n7191) );
  INV_X4 U5937 ( .A(n6333), .ZN(n5482) );
  NAND2_X2 U5938 ( .A1(n4789), .A2(n5482), .ZN(n7299) );
  INV_X4 U5939 ( .A(n7191), .ZN(n5483) );
  INV_X4 U5940 ( .A(n7982), .ZN(n7565) );
  AOI22_X2 U5941 ( .A1(n8404), .A2(n4312), .B1(n8430), .B2(n6258), .ZN(n5484)
         );
  OAI221_X2 U5942 ( .B1(n5644), .B2(n7393), .C1(n5946), .C2(n4317), .A(n5484), 
        .ZN(n7687) );
  INV_X4 U5943 ( .A(n7685), .ZN(n8427) );
  INV_X4 U5944 ( .A(n7687), .ZN(n5488) );
  AOI211_X2 U5945 ( .C1(n7219), .C2(n7686), .A(n5490), .B(n5489), .ZN(n7680)
         );
  AOI221_X2 U5946 ( .B1(n7683), .B2(n7623), .C1(n5492), .C2(n7682), .A(n5491), 
        .ZN(n7681) );
  NAND2_X2 U5947 ( .A1(n5494), .A2(n5493), .ZN(n5496) );
  NAND2_X2 U5948 ( .A1(n5496), .A2(n5495), .ZN(n6934) );
  INV_X4 U5949 ( .A(n5500), .ZN(n5584) );
  INV_X4 U5950 ( .A(n5504), .ZN(n5542) );
  INV_X4 U5951 ( .A(n5508), .ZN(n5546) );
  OAI21_X4 U5952 ( .B1(n5511), .B2(n5510), .A(n5509), .ZN(n5512) );
  INV_X4 U5953 ( .A(n5512), .ZN(n5550) );
  INV_X4 U5954 ( .A(n5516), .ZN(n5554) );
  INV_X4 U5955 ( .A(n5520), .ZN(n5558) );
  NAND2_X2 U5956 ( .A1(n4750), .A2(n4737), .ZN(n5521) );
  NAND2_X2 U5957 ( .A1(n4753), .A2(n6365), .ZN(n5522) );
  NAND2_X2 U5958 ( .A1(n5521), .A2(n5522), .ZN(n5523) );
  INV_X4 U5959 ( .A(n5522), .ZN(n5565) );
  NAND2_X2 U5960 ( .A1(n5523), .A2(n5561), .ZN(n5562) );
  OAI21_X4 U5961 ( .B1(n5526), .B2(n5525), .A(n5524), .ZN(n5560) );
  XNOR2_X2 U5962 ( .A(n5562), .B(n5560), .ZN(n5527) );
  NAND2_X2 U5963 ( .A1(n4144), .A2(n5527), .ZN(n5556) );
  INV_X4 U5964 ( .A(n5557), .ZN(n5528) );
  XNOR2_X2 U5965 ( .A(n5558), .B(n5528), .ZN(n5529) );
  NAND2_X2 U5966 ( .A1(n4161), .A2(n5529), .ZN(n5552) );
  INV_X4 U5967 ( .A(n5553), .ZN(n5530) );
  XNOR2_X2 U5968 ( .A(n5554), .B(n5530), .ZN(n5531) );
  NAND2_X2 U5969 ( .A1(n4245), .A2(n5531), .ZN(n5548) );
  INV_X4 U5970 ( .A(n5549), .ZN(n5532) );
  XNOR2_X2 U5971 ( .A(n5550), .B(n5532), .ZN(n5533) );
  NAND2_X2 U5972 ( .A1(n4192), .A2(n5533), .ZN(n5544) );
  INV_X4 U5973 ( .A(n5545), .ZN(n5534) );
  XNOR2_X2 U5974 ( .A(n5546), .B(n5534), .ZN(n5535) );
  NAND2_X2 U5975 ( .A1(n4198), .A2(n5535), .ZN(n5540) );
  INV_X4 U5976 ( .A(n5541), .ZN(n5536) );
  XNOR2_X2 U5977 ( .A(n5542), .B(n5536), .ZN(n5537) );
  NAND2_X2 U5978 ( .A1(n4247), .A2(n5537), .ZN(n5538) );
  INV_X4 U5979 ( .A(n5539), .ZN(n5602) );
  INV_X4 U5980 ( .A(n5543), .ZN(n5606) );
  INV_X4 U5981 ( .A(n5547), .ZN(n5610) );
  INV_X4 U5982 ( .A(n5551), .ZN(n5614) );
  INV_X4 U5983 ( .A(n5555), .ZN(n5618) );
  INV_X4 U5984 ( .A(n5559), .ZN(n5622) );
  INV_X4 U5985 ( .A(n5560), .ZN(n5563) );
  INV_X4 U5986 ( .A(n5564), .ZN(n5629) );
  INV_X4 U5987 ( .A(n7648), .ZN(n7549) );
  NAND2_X2 U5988 ( .A1(n4752), .A2(n7549), .ZN(n5566) );
  NAND4_X2 U5989 ( .A1(n5567), .A2(n5702), .A3(n5627), .A4(n5566), .ZN(n5628)
         );
  INV_X4 U5990 ( .A(n5628), .ZN(n5568) );
  XNOR2_X2 U5991 ( .A(n5629), .B(n5568), .ZN(n5569) );
  NAND2_X2 U5992 ( .A1(n4145), .A2(n5569), .ZN(n5620) );
  INV_X4 U5993 ( .A(n5621), .ZN(n5570) );
  XNOR2_X2 U5994 ( .A(n5622), .B(n5570), .ZN(n5571) );
  NAND2_X2 U5995 ( .A1(n4153), .A2(n5571), .ZN(n5616) );
  INV_X4 U5996 ( .A(n5617), .ZN(n5572) );
  XNOR2_X2 U5997 ( .A(n5618), .B(n5572), .ZN(n5573) );
  NAND2_X2 U5998 ( .A1(n4258), .A2(n5573), .ZN(n5612) );
  INV_X4 U5999 ( .A(n5613), .ZN(n5574) );
  XNOR2_X2 U6000 ( .A(n5614), .B(n5574), .ZN(n5575) );
  NAND2_X2 U6001 ( .A1(n4217), .A2(n5575), .ZN(n5608) );
  INV_X4 U6002 ( .A(n5609), .ZN(n5576) );
  XNOR2_X2 U6003 ( .A(n5610), .B(n5576), .ZN(n5577) );
  NAND2_X2 U6004 ( .A1(n4199), .A2(n5577), .ZN(n5604) );
  INV_X4 U6005 ( .A(n5605), .ZN(n5578) );
  XNOR2_X2 U6006 ( .A(n5606), .B(n5578), .ZN(n5579) );
  NAND2_X2 U6007 ( .A1(n4118), .A2(n5579), .ZN(n5600) );
  INV_X4 U6008 ( .A(n5601), .ZN(n5580) );
  XNOR2_X2 U6009 ( .A(n5602), .B(n5580), .ZN(n6936) );
  INV_X4 U6010 ( .A(n6936), .ZN(n6554) );
  OAI22_X2 U6011 ( .A1(n4169), .A2(n6934), .B1(n6554), .B2(n4784), .ZN(n5581)
         );
  NAND2_X2 U6012 ( .A1(n4265), .A2(n5581), .ZN(n5596) );
  NAND2_X2 U6013 ( .A1(n4479), .A2(n5582), .ZN(n7890) );
  INV_X4 U6014 ( .A(n5583), .ZN(n5585) );
  XNOR2_X2 U6015 ( .A(n5585), .B(n5584), .ZN(n6924) );
  INV_X4 U6016 ( .A(n6924), .ZN(n5591) );
  INV_X4 U6017 ( .A(n6897), .ZN(n7437) );
  NAND2_X2 U6018 ( .A1(n7437), .A2(n7212), .ZN(n5587) );
  MUX2_X2 U6019 ( .A(n5587), .B(n7212), .S(n4752), .Z(n5588) );
  NAND2_X2 U6020 ( .A1(n7273), .A2(n4205), .ZN(n5590) );
  OAI21_X4 U6021 ( .B1(n5591), .B2(n4784), .A(n5590), .ZN(n5592) );
  INV_X4 U6022 ( .A(n5595), .ZN(n7711) );
  INV_X4 U6023 ( .A(n5597), .ZN(n7688) );
  XNOR2_X2 U6024 ( .A(n5599), .B(n5598), .ZN(n6045) );
  INV_X4 U6025 ( .A(n6045), .ZN(n6884) );
  INV_X4 U6026 ( .A(n5603), .ZN(n5673) );
  INV_X4 U6027 ( .A(n5607), .ZN(n5677) );
  INV_X4 U6028 ( .A(n5611), .ZN(n5681) );
  INV_X4 U6029 ( .A(n5615), .ZN(n5685) );
  INV_X4 U6030 ( .A(n5619), .ZN(n5689) );
  INV_X4 U6031 ( .A(n5623), .ZN(n5693) );
  NAND2_X2 U6032 ( .A1(n7623), .A2(n4753), .ZN(n5624) );
  INV_X4 U6033 ( .A(n5624), .ZN(n5625) );
  NAND2_X2 U6034 ( .A1(n4393), .A2(n7648), .ZN(n5696) );
  NAND2_X2 U6035 ( .A1(n5626), .A2(n5696), .ZN(n5697) );
  XNOR2_X2 U6036 ( .A(n5697), .B(n5695), .ZN(n5630) );
  NAND2_X2 U6037 ( .A1(n4146), .A2(n5630), .ZN(n5691) );
  INV_X4 U6038 ( .A(n5692), .ZN(n5631) );
  XNOR2_X2 U6039 ( .A(n5693), .B(n5631), .ZN(n5632) );
  NAND2_X2 U6040 ( .A1(n4154), .A2(n5632), .ZN(n5687) );
  INV_X4 U6041 ( .A(n5688), .ZN(n5633) );
  XNOR2_X2 U6042 ( .A(n5689), .B(n5633), .ZN(n5634) );
  NAND2_X2 U6043 ( .A1(n4214), .A2(n5634), .ZN(n5683) );
  INV_X4 U6044 ( .A(n5684), .ZN(n5635) );
  XNOR2_X2 U6045 ( .A(n5685), .B(n5635), .ZN(n5636) );
  NAND2_X2 U6046 ( .A1(n4193), .A2(n5636), .ZN(n5679) );
  INV_X4 U6047 ( .A(n5680), .ZN(n5637) );
  XNOR2_X2 U6048 ( .A(n5681), .B(n5637), .ZN(n5638) );
  NAND2_X2 U6049 ( .A1(n4200), .A2(n5638), .ZN(n5675) );
  INV_X4 U6050 ( .A(n5676), .ZN(n5639) );
  XNOR2_X2 U6051 ( .A(n5677), .B(n5639), .ZN(n5640) );
  NAND2_X2 U6052 ( .A1(n4270), .A2(n5640), .ZN(n5671) );
  INV_X4 U6053 ( .A(n5672), .ZN(n5641) );
  XNOR2_X2 U6054 ( .A(n5673), .B(n5641), .ZN(n6883) );
  MUX2_X2 U6055 ( .A(n4460), .B(n6883), .S(n4078), .Z(n5642) );
  NAND2_X2 U6056 ( .A1(n4460), .A2(n4267), .ZN(n5718) );
  INV_X4 U6057 ( .A(n8428), .ZN(n5643) );
  AOI22_X2 U6058 ( .A1(n6258), .A2(n5643), .B1(n8404), .B2(n4735), .ZN(n5646)
         );
  NAND2_X2 U6059 ( .A1(n8430), .A2(n4312), .ZN(n5645) );
  NAND2_X2 U6060 ( .A1(n8430), .A2(n6254), .ZN(n5650) );
  NAND2_X2 U6061 ( .A1(n8443), .A2(n6254), .ZN(n5655) );
  OAI211_X2 U6062 ( .C1(n8444), .C2(n7393), .A(n5655), .B(n5654), .ZN(n5812)
         );
  INV_X4 U6063 ( .A(n5812), .ZN(n7505) );
  INV_X4 U6064 ( .A(n7699), .ZN(n5976) );
  INV_X4 U6065 ( .A(n7700), .ZN(n5656) );
  NAND2_X2 U6066 ( .A1(n4735), .A2(n5800), .ZN(n5662) );
  AOI22_X2 U6067 ( .A1(n6254), .A2(n5660), .B1(n8443), .B2(n6258), .ZN(n5661)
         );
  INV_X4 U6068 ( .A(n7634), .ZN(n7552) );
  NAND2_X2 U6069 ( .A1(n7552), .A2(n4077), .ZN(n5664) );
  AND2_X2 U6070 ( .A1(n7697), .A2(n7634), .ZN(n5665) );
  AOI211_X2 U6071 ( .C1(n7219), .C2(n7695), .A(n5666), .B(n5665), .ZN(n7694)
         );
  NAND2_X2 U6072 ( .A1(n5668), .A2(n5667), .ZN(n5670) );
  NAND2_X2 U6073 ( .A1(n5670), .A2(n5669), .ZN(n7058) );
  INV_X4 U6074 ( .A(n5674), .ZN(n5726) );
  INV_X4 U6075 ( .A(n5678), .ZN(n5730) );
  INV_X4 U6076 ( .A(n5682), .ZN(n5734) );
  INV_X4 U6077 ( .A(n5686), .ZN(n5738) );
  INV_X4 U6078 ( .A(n5690), .ZN(n5742) );
  INV_X4 U6079 ( .A(n5694), .ZN(n5746) );
  INV_X4 U6080 ( .A(n5695), .ZN(n5698) );
  OAI21_X4 U6081 ( .B1(n5698), .B2(n5697), .A(n5696), .ZN(n5699) );
  INV_X4 U6082 ( .A(n5699), .ZN(n5753) );
  INV_X4 U6083 ( .A(n7623), .ZN(n5700) );
  NAND2_X2 U6084 ( .A1(n4393), .A2(n7628), .ZN(n5751) );
  INV_X4 U6085 ( .A(n7628), .ZN(n7553) );
  NAND2_X2 U6086 ( .A1(n4752), .A2(n7553), .ZN(n5701) );
  NAND4_X2 U6087 ( .A1(n5703), .A2(n5702), .A3(n5751), .A4(n5701), .ZN(n5752)
         );
  INV_X4 U6088 ( .A(n5752), .ZN(n5704) );
  XNOR2_X2 U6089 ( .A(n5753), .B(n5704), .ZN(n5705) );
  NAND2_X2 U6090 ( .A1(n4141), .A2(n5705), .ZN(n5744) );
  INV_X4 U6091 ( .A(n5745), .ZN(n5706) );
  XNOR2_X2 U6092 ( .A(n5746), .B(n5706), .ZN(n5707) );
  NAND2_X2 U6093 ( .A1(n4260), .A2(n5707), .ZN(n5740) );
  INV_X4 U6094 ( .A(n5741), .ZN(n5708) );
  XNOR2_X2 U6095 ( .A(n5742), .B(n5708), .ZN(n5709) );
  NAND2_X2 U6096 ( .A1(n4228), .A2(n5709), .ZN(n5736) );
  INV_X4 U6097 ( .A(n5737), .ZN(n5710) );
  XNOR2_X2 U6098 ( .A(n5738), .B(n5710), .ZN(n5711) );
  NAND2_X2 U6099 ( .A1(n4194), .A2(n5711), .ZN(n5732) );
  INV_X4 U6100 ( .A(n5733), .ZN(n5712) );
  XNOR2_X2 U6101 ( .A(n5734), .B(n5712), .ZN(n5713) );
  NAND2_X2 U6102 ( .A1(n4201), .A2(n5713), .ZN(n5728) );
  INV_X4 U6103 ( .A(n5729), .ZN(n5714) );
  XNOR2_X2 U6104 ( .A(n5730), .B(n5714), .ZN(n5715) );
  NAND2_X2 U6105 ( .A1(n4246), .A2(n5715), .ZN(n5724) );
  INV_X4 U6106 ( .A(n5725), .ZN(n5716) );
  XNOR2_X2 U6107 ( .A(n5726), .B(n5716), .ZN(n7059) );
  INV_X4 U6108 ( .A(n7059), .ZN(n6571) );
  OAI22_X2 U6109 ( .A1(n4169), .A2(n7058), .B1(n6571), .B2(n4784), .ZN(n5717)
         );
  NAND2_X2 U6110 ( .A1(n4305), .A2(n5717), .ZN(n5719) );
  INV_X4 U6111 ( .A(n7910), .ZN(n5720) );
  INV_X4 U6112 ( .A(n5721), .ZN(n7701) );
  XNOR2_X2 U6113 ( .A(n5723), .B(n5722), .ZN(n5951) );
  INV_X4 U6114 ( .A(n5951), .ZN(n7046) );
  INV_X4 U6115 ( .A(n5727), .ZN(n5986) );
  INV_X4 U6116 ( .A(n5731), .ZN(n5990) );
  INV_X4 U6117 ( .A(n5735), .ZN(n5994) );
  INV_X4 U6118 ( .A(n5739), .ZN(n5998) );
  INV_X4 U6119 ( .A(n5743), .ZN(n6002) );
  INV_X4 U6120 ( .A(n5747), .ZN(n6006) );
  NAND2_X2 U6121 ( .A1(n7634), .A2(n4753), .ZN(n5748) );
  INV_X4 U6122 ( .A(n5748), .ZN(n5749) );
  NAND2_X2 U6123 ( .A1(n4395), .A2(n7628), .ZN(n6009) );
  NAND2_X2 U6124 ( .A1(n5750), .A2(n6009), .ZN(n6010) );
  XNOR2_X2 U6125 ( .A(n6010), .B(n6008), .ZN(n5754) );
  NAND2_X2 U6126 ( .A1(n4147), .A2(n5754), .ZN(n6004) );
  INV_X4 U6127 ( .A(n6005), .ZN(n5755) );
  XNOR2_X2 U6128 ( .A(n6006), .B(n5755), .ZN(n5756) );
  NAND2_X2 U6129 ( .A1(n4179), .A2(n5756), .ZN(n6000) );
  INV_X4 U6130 ( .A(n6001), .ZN(n5757) );
  XNOR2_X2 U6131 ( .A(n6002), .B(n5757), .ZN(n5758) );
  NAND2_X2 U6132 ( .A1(n4261), .A2(n5758), .ZN(n5996) );
  INV_X4 U6133 ( .A(n5997), .ZN(n5759) );
  XNOR2_X2 U6134 ( .A(n5998), .B(n5759), .ZN(n5760) );
  NAND2_X2 U6135 ( .A1(n4195), .A2(n5760), .ZN(n5992) );
  INV_X4 U6136 ( .A(n5993), .ZN(n5761) );
  XNOR2_X2 U6137 ( .A(n5994), .B(n5761), .ZN(n5762) );
  NAND2_X2 U6138 ( .A1(n4202), .A2(n5762), .ZN(n5988) );
  INV_X4 U6139 ( .A(n5989), .ZN(n5763) );
  XNOR2_X2 U6140 ( .A(n5990), .B(n5763), .ZN(n5764) );
  NAND2_X2 U6141 ( .A1(n4259), .A2(n5764), .ZN(n5984) );
  INV_X4 U6142 ( .A(n5985), .ZN(n5765) );
  XNOR2_X2 U6143 ( .A(n5986), .B(n5765), .ZN(n7045) );
  MUX2_X2 U6144 ( .A(n4461), .B(n7045), .S(n4078), .Z(n5766) );
  NAND2_X2 U6145 ( .A1(n4461), .A2(n4268), .ZN(n6030) );
  INV_X4 U6146 ( .A(n5767), .ZN(n7550) );
  INV_X4 U6147 ( .A(n7379), .ZN(n7547) );
  INV_X4 U6148 ( .A(n8306), .ZN(n7528) );
  NAND2_X2 U6149 ( .A1(n4711), .A2(n4080), .ZN(n5770) );
  NAND2_X2 U6150 ( .A1(memAddr[28]), .A2(n6078), .ZN(n5769) );
  NAND2_X2 U6151 ( .A1(n4748), .A2(regWrData[28]), .ZN(n5768) );
  INV_X4 U6152 ( .A(n8316), .ZN(n7504) );
  NAND2_X2 U6153 ( .A1(n4714), .A2(n4080), .ZN(n5773) );
  NAND2_X2 U6154 ( .A1(memAddr[29]), .A2(n6078), .ZN(n5772) );
  NAND2_X2 U6155 ( .A1(n4748), .A2(regWrData[29]), .ZN(n5771) );
  INV_X4 U6156 ( .A(n8304), .ZN(n7503) );
  NAND2_X2 U6157 ( .A1(n4746), .A2(memAddr[27]), .ZN(n5775) );
  NAND2_X2 U6158 ( .A1(n4748), .A2(regWrData[27]), .ZN(n5774) );
  NAND2_X2 U6159 ( .A1(n4080), .A2(n4475), .ZN(n5778) );
  NAND2_X2 U6160 ( .A1(n4746), .A2(memAddr[26]), .ZN(n5777) );
  NAND2_X2 U6161 ( .A1(n4748), .A2(regWrData[26]), .ZN(n5776) );
  NAND2_X2 U6162 ( .A1(n4746), .A2(memAddr[25]), .ZN(n5780) );
  NAND2_X2 U6163 ( .A1(n4748), .A2(regWrData[25]), .ZN(n5779) );
  NAND2_X2 U6164 ( .A1(n4746), .A2(memAddr[24]), .ZN(n5782) );
  NAND2_X2 U6165 ( .A1(n4748), .A2(regWrData[24]), .ZN(n5781) );
  INV_X4 U6166 ( .A(n8326), .ZN(n7527) );
  INV_X4 U6167 ( .A(n8364), .ZN(n7529) );
  NAND2_X2 U6168 ( .A1(n4746), .A2(memAddr[21]), .ZN(n5784) );
  NAND2_X2 U6169 ( .A1(n4748), .A2(regWrData[21]), .ZN(n5783) );
  INV_X4 U6170 ( .A(n8336), .ZN(n7499) );
  NAND2_X2 U6171 ( .A1(n4080), .A2(n4417), .ZN(n5787) );
  NAND2_X2 U6172 ( .A1(n4746), .A2(memAddr[20]), .ZN(n5786) );
  NAND2_X2 U6173 ( .A1(n4748), .A2(regWrData[20]), .ZN(n5785) );
  INV_X4 U6174 ( .A(n8348), .ZN(n7498) );
  NAND2_X2 U6175 ( .A1(n4746), .A2(memAddr[19]), .ZN(n5789) );
  NAND2_X2 U6176 ( .A1(n4748), .A2(regWrData[19]), .ZN(n5788) );
  INV_X4 U6177 ( .A(n8349), .ZN(n7497) );
  NAND2_X2 U6178 ( .A1(n4746), .A2(memAddr[17]), .ZN(n5791) );
  NAND2_X2 U6179 ( .A1(n4748), .A2(regWrData[17]), .ZN(n5790) );
  INV_X4 U6180 ( .A(n7895), .ZN(n7496) );
  NAND2_X2 U6181 ( .A1(n4746), .A2(memAddr[18]), .ZN(n5793) );
  NAND2_X2 U6182 ( .A1(n4748), .A2(regWrData[18]), .ZN(n5792) );
  INV_X4 U6183 ( .A(n8448), .ZN(n7495) );
  NAND2_X2 U6184 ( .A1(n4746), .A2(memAddr[16]), .ZN(n5795) );
  NAND2_X2 U6185 ( .A1(n4748), .A2(regWrData[16]), .ZN(n5794) );
  INV_X4 U6186 ( .A(n8460), .ZN(n7494) );
  NAND4_X2 U6187 ( .A1(n7514), .A2(n7513), .A3(n4088), .A4(n7512), .ZN(n7724)
         );
  INV_X4 U6188 ( .A(n5796), .ZN(n5797) );
  NAND2_X2 U6189 ( .A1(n5797), .A2(n4791), .ZN(n7725) );
  NAND2_X2 U6190 ( .A1(n6072), .A2(n4824), .ZN(n7881) );
  INV_X4 U6191 ( .A(n7881), .ZN(n7493) );
  NAND2_X2 U6192 ( .A1(n7427), .A2(n4091), .ZN(n7293) );
  AOI22_X2 U6193 ( .A1(n6254), .A2(n5800), .B1(n8443), .B2(n4312), .ZN(n5804)
         );
  NAND2_X2 U6194 ( .A1(n5804), .A2(n5803), .ZN(n7898) );
  INV_X4 U6195 ( .A(n7412), .ZN(n7894) );
  INV_X4 U6196 ( .A(n5805), .ZN(n7518) );
  INV_X4 U6197 ( .A(n4738), .ZN(n6040) );
  INV_X4 U6198 ( .A(n8324), .ZN(n7491) );
  INV_X4 U6199 ( .A(n8323), .ZN(n7490) );
  NAND2_X2 U6200 ( .A1(n7219), .A2(n4091), .ZN(n8340) );
  INV_X4 U6201 ( .A(n8444), .ZN(n5807) );
  AOI22_X2 U6202 ( .A1(n4312), .A2(n5807), .B1(n6258), .B2(n5806), .ZN(n5810)
         );
  INV_X4 U6203 ( .A(n8416), .ZN(n5808) );
  AOI22_X2 U6204 ( .A1(n6254), .A2(n5808), .B1(n8443), .B2(n4735), .ZN(n5809)
         );
  NAND2_X2 U6205 ( .A1(n5810), .A2(n5809), .ZN(n7900) );
  AOI221_X2 U6206 ( .B1(n6040), .B2(n5812), .C1(n7209), .C2(n7695), .A(n5811), 
        .ZN(n7904) );
  INV_X4 U6207 ( .A(n5813), .ZN(n5814) );
  NAND2_X2 U6208 ( .A1(n5814), .A2(n7906), .ZN(n5816) );
  NAND2_X2 U6209 ( .A1(n7907), .A2(n7628), .ZN(n5815) );
  NAND2_X2 U6210 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  AOI21_X2 U6211 ( .B1(n7219), .B2(n7687), .A(n5817), .ZN(n7905) );
  NAND2_X2 U6212 ( .A1(n7657), .A2(n8502), .ZN(n5818) );
  INV_X4 U6213 ( .A(n7722), .ZN(n7501) );
  NAND3_X2 U6214 ( .A1(n8500), .A2(n5818), .A3(n4504), .ZN(n7383) );
  NAND2_X2 U6215 ( .A1(n4735), .A2(n7383), .ZN(n5824) );
  INV_X4 U6216 ( .A(n7720), .ZN(n6942) );
  NAND2_X2 U6217 ( .A1(n7661), .A2(n8502), .ZN(n5819) );
  OAI211_X2 U6218 ( .C1(n8486), .C2(n6942), .A(n5819), .B(n8487), .ZN(n7391)
         );
  NAND2_X2 U6219 ( .A1(n6254), .A2(n7391), .ZN(n5823) );
  NAND3_X2 U6220 ( .A1(n5824), .A2(n5823), .A3(n5822), .ZN(n7921) );
  NAND2_X2 U6221 ( .A1(n6258), .A2(n5825), .ZN(n5828) );
  NAND2_X2 U6222 ( .A1(n4312), .A2(n5930), .ZN(n5827) );
  OAI211_X2 U6223 ( .C1(n8440), .C2(n7525), .A(n8509), .B(n8510), .ZN(n6250)
         );
  AOI22_X2 U6224 ( .A1(n6254), .A2(n6250), .B1(n4735), .B2(n6257), .ZN(n5826)
         );
  NAND3_X2 U6225 ( .A1(n5828), .A2(n5827), .A3(n5826), .ZN(n7971) );
  OAI221_X2 U6226 ( .B1(n8341), .B2(n7393), .C1(n8393), .C2(n4317), .A(n5830), 
        .ZN(n5953) );
  AOI22_X2 U6227 ( .A1(n5831), .A2(n7918), .B1(n6040), .B2(n5953), .ZN(n5835)
         );
  NAND2_X2 U6228 ( .A1(n5935), .A2(n7546), .ZN(n5929) );
  OAI211_X2 U6229 ( .C1(n8402), .C2(n4317), .A(n5929), .B(n4127), .ZN(n7291)
         );
  NAND2_X2 U6230 ( .A1(n7427), .A2(n7291), .ZN(n5834) );
  NAND2_X2 U6231 ( .A1(n7919), .A2(n7661), .ZN(n5833) );
  AOI22_X2 U6232 ( .A1(n7209), .A2(n7971), .B1(n7219), .B2(n7921), .ZN(n5832)
         );
  NAND4_X2 U6233 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n7464)
         );
  MUX2_X2 U6234 ( .A(n7570), .B(n7058), .S(n4078), .Z(n7462) );
  AOI211_X2 U6235 ( .C1(n7507), .C2(n7464), .A(n5837), .B(n5836), .ZN(n7916)
         );
  NAND2_X2 U6236 ( .A1(n8903), .A2(n7123), .ZN(n6331) );
  NAND2_X2 U6237 ( .A1(n7123), .A2(n4090), .ZN(n6332) );
  NAND2_X2 U6238 ( .A1(n4745), .A2(n4486), .ZN(n5839) );
  NAND2_X2 U6239 ( .A1(n4744), .A2(n4510), .ZN(n5838) );
  OAI211_X2 U6240 ( .C1(n8192), .C2(n4755), .A(n5839), .B(n5838), .ZN(iAddr[3]) );
  NAND2_X2 U6241 ( .A1(n4745), .A2(n4489), .ZN(n5841) );
  NAND2_X2 U6242 ( .A1(n4744), .A2(n4556), .ZN(n5840) );
  OAI211_X2 U6243 ( .C1(n8204), .C2(n4755), .A(n5841), .B(n5840), .ZN(iAddr[2]) );
  NAND2_X2 U6244 ( .A1(n4745), .A2(n4485), .ZN(n5843) );
  NAND2_X2 U6245 ( .A1(n4744), .A2(n4511), .ZN(n5842) );
  OAI211_X2 U6246 ( .C1(n8189), .C2(n6331), .A(n5843), .B(n5842), .ZN(iAddr[4]) );
  NAND2_X2 U6247 ( .A1(n4745), .A2(n4484), .ZN(n5845) );
  NAND2_X2 U6248 ( .A1(n4744), .A2(n4512), .ZN(n5844) );
  OAI211_X2 U6249 ( .C1(n8186), .C2(n6331), .A(n5845), .B(n5844), .ZN(iAddr[5]) );
  NAND2_X2 U6250 ( .A1(n4745), .A2(n4488), .ZN(n5847) );
  NAND2_X2 U6251 ( .A1(n4744), .A2(n4513), .ZN(n5846) );
  OAI211_X2 U6252 ( .C1(n8183), .C2(n6331), .A(n5847), .B(n5846), .ZN(iAddr[6]) );
  NAND2_X2 U6253 ( .A1(iAddr[3]), .A2(iAddr[2]), .ZN(n6048) );
  INV_X4 U6254 ( .A(n6048), .ZN(n6050) );
  NAND2_X2 U6255 ( .A1(n6050), .A2(iAddr[4]), .ZN(n6049) );
  INV_X4 U6256 ( .A(n6049), .ZN(n6051) );
  NAND2_X2 U6257 ( .A1(n6051), .A2(iAddr[5]), .ZN(n6052) );
  INV_X4 U6258 ( .A(n6052), .ZN(n5848) );
  NAND2_X2 U6259 ( .A1(n5848), .A2(iAddr[6]), .ZN(n8040) );
  NAND2_X2 U6260 ( .A1(n4745), .A2(n4483), .ZN(n5850) );
  NAND2_X2 U6261 ( .A1(n4744), .A2(n4514), .ZN(n5849) );
  OAI211_X2 U6262 ( .C1(n8180), .C2(n6331), .A(n5850), .B(n5849), .ZN(iAddr[7]) );
  NAND2_X2 U6263 ( .A1(n4745), .A2(n4490), .ZN(n5852) );
  NAND2_X2 U6264 ( .A1(n4744), .A2(n4515), .ZN(n5851) );
  OAI211_X2 U6265 ( .C1(n8177), .C2(n6331), .A(n5852), .B(n5851), .ZN(iAddr[8]) );
  INV_X4 U6266 ( .A(n8040), .ZN(n6054) );
  NAND2_X2 U6267 ( .A1(iAddr[7]), .A2(n6054), .ZN(n6055) );
  INV_X4 U6268 ( .A(n6055), .ZN(n5853) );
  NAND2_X2 U6269 ( .A1(n5853), .A2(iAddr[8]), .ZN(n8052) );
  NAND2_X2 U6270 ( .A1(n4745), .A2(n4482), .ZN(n5855) );
  NAND2_X2 U6271 ( .A1(n4744), .A2(n4516), .ZN(n5854) );
  OAI211_X2 U6272 ( .C1(n8174), .C2(n4755), .A(n5855), .B(n5854), .ZN(iAddr[9]) );
  NAND2_X2 U6273 ( .A1(n4745), .A2(n4492), .ZN(n5857) );
  NAND2_X2 U6274 ( .A1(n4744), .A2(n4517), .ZN(n5856) );
  OAI211_X2 U6275 ( .C1(n8265), .C2(n4755), .A(n5857), .B(n5856), .ZN(
        iAddr[10]) );
  INV_X4 U6276 ( .A(n8052), .ZN(n6057) );
  NAND2_X2 U6277 ( .A1(iAddr[9]), .A2(n6057), .ZN(n6058) );
  INV_X4 U6278 ( .A(n6058), .ZN(n5858) );
  NAND2_X2 U6279 ( .A1(n5858), .A2(iAddr[10]), .ZN(n8064) );
  NAND2_X2 U6280 ( .A1(n4745), .A2(n4481), .ZN(n5860) );
  NAND2_X2 U6281 ( .A1(n4744), .A2(n4518), .ZN(n5859) );
  OAI211_X2 U6282 ( .C1(n8262), .C2(n4755), .A(n5860), .B(n5859), .ZN(
        iAddr[11]) );
  NAND2_X2 U6283 ( .A1(n4745), .A2(n4491), .ZN(n5862) );
  NAND2_X2 U6284 ( .A1(n4744), .A2(n4519), .ZN(n5861) );
  OAI211_X2 U6285 ( .C1(n8259), .C2(n4755), .A(n5862), .B(n5861), .ZN(
        iAddr[12]) );
  INV_X4 U6286 ( .A(n8064), .ZN(n6060) );
  NAND2_X2 U6287 ( .A1(iAddr[11]), .A2(n6060), .ZN(n6061) );
  INV_X4 U6288 ( .A(n6061), .ZN(n5863) );
  NAND2_X2 U6289 ( .A1(n5863), .A2(iAddr[12]), .ZN(n8076) );
  NAND2_X2 U6290 ( .A1(n4745), .A2(n4480), .ZN(n5865) );
  NAND2_X2 U6291 ( .A1(n4744), .A2(n4520), .ZN(n5864) );
  OAI211_X2 U6292 ( .C1(n8256), .C2(n4755), .A(n5865), .B(n5864), .ZN(
        iAddr[13]) );
  NAND2_X2 U6293 ( .A1(n4745), .A2(n4487), .ZN(n5867) );
  NAND2_X2 U6294 ( .A1(n4744), .A2(n4521), .ZN(n5866) );
  OAI211_X2 U6295 ( .C1(n8253), .C2(n4755), .A(n5867), .B(n5866), .ZN(
        iAddr[14]) );
  INV_X4 U6296 ( .A(n8076), .ZN(n6063) );
  NAND2_X2 U6297 ( .A1(iAddr[13]), .A2(n6063), .ZN(n6064) );
  INV_X4 U6298 ( .A(n6064), .ZN(n5868) );
  NAND2_X2 U6299 ( .A1(n5868), .A2(iAddr[14]), .ZN(n8000) );
  NAND2_X2 U6300 ( .A1(n4745), .A2(n4578), .ZN(n5870) );
  NAND2_X2 U6301 ( .A1(n4744), .A2(n4522), .ZN(n5869) );
  OAI211_X2 U6302 ( .C1(n8250), .C2(n4755), .A(n5870), .B(n5869), .ZN(
        iAddr[15]) );
  NAND2_X2 U6303 ( .A1(n4745), .A2(n4574), .ZN(n5872) );
  NAND2_X2 U6304 ( .A1(n4744), .A2(n4595), .ZN(n5871) );
  OAI211_X2 U6305 ( .C1(n8247), .C2(n4755), .A(n5872), .B(n5871), .ZN(
        iAddr[16]) );
  INV_X4 U6306 ( .A(n8000), .ZN(n6031) );
  NAND2_X2 U6307 ( .A1(iAddr[15]), .A2(n6031), .ZN(n6032) );
  INV_X4 U6308 ( .A(n6032), .ZN(n5873) );
  NAND2_X2 U6309 ( .A1(n5873), .A2(iAddr[16]), .ZN(n7998) );
  NAND2_X2 U6310 ( .A1(n4745), .A2(n4577), .ZN(n5875) );
  NAND2_X2 U6311 ( .A1(n4744), .A2(n4596), .ZN(n5874) );
  OAI211_X2 U6312 ( .C1(n8244), .C2(n4755), .A(n5875), .B(n5874), .ZN(
        iAddr[17]) );
  NAND2_X2 U6313 ( .A1(n4745), .A2(n4576), .ZN(n5877) );
  NAND2_X2 U6314 ( .A1(n4744), .A2(n4597), .ZN(n5876) );
  OAI211_X2 U6315 ( .C1(n8240), .C2(n4755), .A(n5877), .B(n5876), .ZN(
        iAddr[18]) );
  INV_X4 U6316 ( .A(n7998), .ZN(n6034) );
  NAND2_X2 U6317 ( .A1(iAddr[17]), .A2(n6034), .ZN(n6035) );
  INV_X4 U6318 ( .A(n6035), .ZN(n5878) );
  NAND2_X2 U6319 ( .A1(n5878), .A2(iAddr[18]), .ZN(n7925) );
  NAND2_X2 U6320 ( .A1(n4745), .A2(n4575), .ZN(n5880) );
  NAND2_X2 U6321 ( .A1(n4744), .A2(n4603), .ZN(n5879) );
  OAI211_X2 U6322 ( .C1(n8237), .C2(n4755), .A(n5880), .B(n5879), .ZN(
        iAddr[19]) );
  INV_X4 U6323 ( .A(n7925), .ZN(n5881) );
  NAND2_X2 U6324 ( .A1(iAddr[19]), .A2(n5881), .ZN(n5887) );
  INV_X4 U6325 ( .A(n5882), .ZN(n5883) );
  NAND2_X2 U6326 ( .A1(n4745), .A2(n4579), .ZN(n5886) );
  NAND2_X2 U6327 ( .A1(n4744), .A2(n4604), .ZN(n5885) );
  OAI211_X2 U6328 ( .C1(n8234), .C2(n4755), .A(n5886), .B(n5885), .ZN(
        iAddr[20]) );
  INV_X4 U6329 ( .A(n5887), .ZN(n5888) );
  NAND2_X2 U6330 ( .A1(n5888), .A2(iAddr[20]), .ZN(n5891) );
  NAND2_X2 U6331 ( .A1(n4745), .A2(n4358), .ZN(n5890) );
  NAND2_X2 U6332 ( .A1(n4744), .A2(n4605), .ZN(n5889) );
  OAI211_X2 U6333 ( .C1(n8231), .C2(n4755), .A(n5890), .B(n5889), .ZN(
        iAddr[21]) );
  INV_X4 U6334 ( .A(n5891), .ZN(n5892) );
  NAND2_X2 U6335 ( .A1(n5892), .A2(iAddr[21]), .ZN(n5897) );
  NAND2_X2 U6336 ( .A1(n4745), .A2(n4357), .ZN(n5894) );
  NAND2_X2 U6337 ( .A1(n4744), .A2(n4598), .ZN(n5893) );
  OAI211_X2 U6338 ( .C1(n8228), .C2(n4755), .A(n5894), .B(n5893), .ZN(
        iAddr[22]) );
  NAND2_X2 U6339 ( .A1(n4745), .A2(n4349), .ZN(n5896) );
  NAND2_X2 U6340 ( .A1(n4744), .A2(n4606), .ZN(n5895) );
  OAI211_X2 U6341 ( .C1(n8225), .C2(n4755), .A(n5896), .B(n5895), .ZN(
        iAddr[23]) );
  INV_X4 U6342 ( .A(n5897), .ZN(n6038) );
  NAND2_X2 U6343 ( .A1(n6038), .A2(iAddr[22]), .ZN(n6037) );
  INV_X4 U6344 ( .A(n6037), .ZN(n5898) );
  NAND2_X2 U6345 ( .A1(n5898), .A2(iAddr[23]), .ZN(n5901) );
  NAND2_X2 U6346 ( .A1(n4745), .A2(n4350), .ZN(n5900) );
  NAND2_X2 U6347 ( .A1(n4744), .A2(n4607), .ZN(n5899) );
  OAI211_X2 U6348 ( .C1(n8222), .C2(n4755), .A(n5900), .B(n5899), .ZN(
        iAddr[24]) );
  INV_X4 U6349 ( .A(n5901), .ZN(n5902) );
  NAND2_X2 U6350 ( .A1(n5902), .A2(iAddr[24]), .ZN(n5905) );
  NAND2_X2 U6351 ( .A1(n4745), .A2(n4355), .ZN(n5904) );
  NAND2_X2 U6352 ( .A1(n4744), .A2(n4608), .ZN(n5903) );
  OAI211_X2 U6353 ( .C1(n8219), .C2(n4755), .A(n5904), .B(n5903), .ZN(
        iAddr[25]) );
  INV_X4 U6354 ( .A(n5905), .ZN(n5906) );
  NAND2_X2 U6355 ( .A1(n5906), .A2(iAddr[25]), .ZN(n5909) );
  NAND2_X2 U6356 ( .A1(n4745), .A2(n4351), .ZN(n5908) );
  NAND2_X2 U6357 ( .A1(n4744), .A2(n4609), .ZN(n5907) );
  OAI211_X2 U6358 ( .C1(n8216), .C2(n4755), .A(n5908), .B(n5907), .ZN(
        iAddr[26]) );
  INV_X4 U6359 ( .A(n5909), .ZN(n5910) );
  NAND2_X2 U6360 ( .A1(n5910), .A2(iAddr[26]), .ZN(n5913) );
  NAND2_X2 U6361 ( .A1(n4745), .A2(n4354), .ZN(n5912) );
  NAND2_X2 U6362 ( .A1(n4744), .A2(n4599), .ZN(n5911) );
  OAI211_X2 U6363 ( .C1(n8213), .C2(n4755), .A(n5912), .B(n5911), .ZN(
        iAddr[27]) );
  INV_X4 U6364 ( .A(n5913), .ZN(n5914) );
  NAND2_X2 U6365 ( .A1(n5914), .A2(iAddr[27]), .ZN(n5917) );
  INV_X4 U6366 ( .A(n7666), .ZN(n7487) );
  NAND2_X2 U6367 ( .A1(n4745), .A2(n4352), .ZN(n5916) );
  NAND2_X2 U6368 ( .A1(n4744), .A2(n4600), .ZN(n5915) );
  OAI211_X2 U6369 ( .C1(n8210), .C2(n4755), .A(n5916), .B(n5915), .ZN(
        iAddr[28]) );
  INV_X4 U6370 ( .A(n5917), .ZN(n5918) );
  NAND2_X2 U6371 ( .A1(n5918), .A2(iAddr[28]), .ZN(n5921) );
  NAND2_X2 U6372 ( .A1(n4745), .A2(n4356), .ZN(n5920) );
  NAND2_X2 U6373 ( .A1(n4744), .A2(n4601), .ZN(n5919) );
  OAI211_X2 U6374 ( .C1(n8207), .C2(n4755), .A(n5920), .B(n5919), .ZN(
        iAddr[29]) );
  INV_X4 U6375 ( .A(n5921), .ZN(n5922) );
  NAND2_X2 U6376 ( .A1(n5922), .A2(iAddr[29]), .ZN(n6067) );
  NAND2_X2 U6377 ( .A1(n4745), .A2(n4353), .ZN(n5924) );
  NAND2_X2 U6378 ( .A1(n4744), .A2(n4602), .ZN(n5923) );
  OAI211_X2 U6379 ( .C1(n8201), .C2(n4755), .A(n5924), .B(n5923), .ZN(
        iAddr[30]) );
  NAND2_X2 U6380 ( .A1(n4387), .A2(n7212), .ZN(n5928) );
  NAND2_X2 U6381 ( .A1(n4381), .A2(n7479), .ZN(n5926) );
  INV_X4 U6382 ( .A(n7212), .ZN(n7470) );
  XNOR2_X2 U6383 ( .A(n7470), .B(n4387), .ZN(n6330) );
  NAND2_X2 U6384 ( .A1(n6329), .A2(n6330), .ZN(n5927) );
  NAND2_X2 U6385 ( .A1(n5928), .A2(n5927), .ZN(n8534) );
  MUX2_X2 U6386 ( .A(n8333), .B(n5941), .S(n6254), .Z(n7207) );
  INV_X4 U6387 ( .A(n7207), .ZN(n7713) );
  OAI221_X2 U6388 ( .B1(n7393), .B2(n6263), .C1(n8341), .C2(n4317), .A(n5929), 
        .ZN(n7962) );
  NAND2_X2 U6389 ( .A1(n8503), .A2(n6254), .ZN(n5933) );
  NAND2_X2 U6390 ( .A1(n6258), .A2(n5930), .ZN(n5932) );
  AOI22_X2 U6391 ( .A1(n4735), .A2(n6250), .B1(n4312), .B2(n6257), .ZN(n5931)
         );
  NAND3_X2 U6392 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(n7295) );
  AOI22_X2 U6393 ( .A1(n4735), .A2(n7391), .B1(n4312), .B2(n7383), .ZN(n5934)
         );
  OAI221_X2 U6394 ( .B1(n5945), .B2(n4128), .C1(n8495), .C2(n4317), .A(n5934), 
        .ZN(n7278) );
  AOI22_X2 U6395 ( .A1(n5936), .A2(n5935), .B1(n7219), .B2(n7278), .ZN(n5937)
         );
  MUX2_X2 U6396 ( .A(n7569), .B(n6934), .S(n4078), .Z(n7456) );
  AOI211_X2 U6397 ( .C1(n7507), .C2(n7458), .A(n5940), .B(n5939), .ZN(n7959)
         );
  INV_X4 U6398 ( .A(n5941), .ZN(n5942) );
  OAI221_X2 U6399 ( .B1(n8402), .B2(n7393), .C1(n8362), .C2(n4317), .A(n5943), 
        .ZN(n7972) );
  NAND2_X2 U6400 ( .A1(n6254), .A2(n7383), .ZN(n5950) );
  NAND3_X2 U6401 ( .A1(n4508), .A2(n5950), .A3(n5949), .ZN(n7980) );
  MUX2_X2 U6402 ( .A(n7568), .B(n5951), .S(n4078), .Z(n5952) );
  INV_X4 U6403 ( .A(n5952), .ZN(n7451) );
  INV_X4 U6404 ( .A(n5953), .ZN(n7488) );
  NAND2_X2 U6405 ( .A1(n4076), .A2(n7972), .ZN(n5958) );
  NAND2_X2 U6406 ( .A1(n7969), .A2(n7659), .ZN(n5957) );
  AOI22_X2 U6407 ( .A1(n7209), .A2(n7980), .B1(n7219), .B2(n7971), .ZN(n5956)
         );
  NAND4_X2 U6408 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n7452)
         );
  AOI221_X2 U6409 ( .B1(n7506), .B2(n7451), .C1(n7507), .C2(n7452), .A(n5960), 
        .ZN(n7966) );
  INV_X4 U6410 ( .A(n7972), .ZN(n8361) );
  NAND2_X2 U6411 ( .A1(n4076), .A2(n7670), .ZN(n5965) );
  NAND2_X2 U6412 ( .A1(n7978), .A2(n7657), .ZN(n5964) );
  AOI22_X2 U6413 ( .A1(n7209), .A2(n7675), .B1(n7219), .B2(n7980), .ZN(n5963)
         );
  OAI22_X2 U6414 ( .A1(n4126), .A2(n5967), .B1(n7656), .B2(n7982), .ZN(n5973)
         );
  NAND2_X2 U6415 ( .A1(n5969), .A2(n5968), .ZN(n5971) );
  NAND2_X2 U6416 ( .A1(n5971), .A2(n5970), .ZN(n7240) );
  MUX2_X2 U6417 ( .A(n7567), .B(n7240), .S(n4078), .Z(n7447) );
  INV_X4 U6418 ( .A(n7900), .ZN(n5974) );
  INV_X4 U6419 ( .A(n7898), .ZN(n5977) );
  OAI22_X2 U6420 ( .A1(n5978), .A2(n5977), .B1(n5976), .B2(n5975), .ZN(n5979)
         );
  INV_X4 U6421 ( .A(n7988), .ZN(n7541) );
  INV_X4 U6422 ( .A(n7641), .ZN(n7551) );
  AND2_X2 U6423 ( .A1(n7989), .A2(n7641), .ZN(n5982) );
  INV_X4 U6424 ( .A(n5987), .ZN(n6289) );
  INV_X4 U6425 ( .A(n5991), .ZN(n6293) );
  INV_X4 U6426 ( .A(n5995), .ZN(n6297) );
  INV_X4 U6427 ( .A(n5999), .ZN(n6301) );
  INV_X4 U6428 ( .A(n6003), .ZN(n6305) );
  OAI21_X4 U6429 ( .B1(n6006), .B2(n6005), .A(n6004), .ZN(n6007) );
  INV_X4 U6430 ( .A(n6007), .ZN(n6167) );
  INV_X4 U6431 ( .A(n6008), .ZN(n6011) );
  OAI21_X4 U6432 ( .B1(n6011), .B2(n6010), .A(n6009), .ZN(n6012) );
  INV_X4 U6433 ( .A(n6012), .ZN(n6085) );
  NAND2_X2 U6434 ( .A1(n4754), .A2(n7552), .ZN(n6015) );
  NAND2_X2 U6435 ( .A1(n4395), .A2(n7641), .ZN(n6083) );
  INV_X4 U6436 ( .A(n6084), .ZN(n6016) );
  XNOR2_X2 U6437 ( .A(n6085), .B(n6016), .ZN(n6017) );
  NAND2_X2 U6438 ( .A1(n4148), .A2(n6017), .ZN(n6165) );
  INV_X4 U6439 ( .A(n6166), .ZN(n6018) );
  XNOR2_X2 U6440 ( .A(n6167), .B(n6018), .ZN(n6019) );
  NAND2_X2 U6441 ( .A1(n4187), .A2(n6019), .ZN(n6303) );
  INV_X4 U6442 ( .A(n6304), .ZN(n6020) );
  XNOR2_X2 U6443 ( .A(n6305), .B(n6020), .ZN(n6021) );
  NAND2_X2 U6444 ( .A1(n4180), .A2(n6021), .ZN(n6299) );
  INV_X4 U6445 ( .A(n6300), .ZN(n6022) );
  XNOR2_X2 U6446 ( .A(n6301), .B(n6022), .ZN(n6023) );
  NAND2_X2 U6447 ( .A1(n4196), .A2(n6023), .ZN(n6295) );
  INV_X4 U6448 ( .A(n6296), .ZN(n6024) );
  XNOR2_X2 U6449 ( .A(n6297), .B(n6024), .ZN(n6025) );
  NAND2_X2 U6450 ( .A1(n4203), .A2(n6025), .ZN(n6291) );
  OAI21_X4 U6451 ( .B1(n4203), .B2(n6025), .A(n6291), .ZN(n6292) );
  INV_X4 U6452 ( .A(n6292), .ZN(n6026) );
  XNOR2_X2 U6453 ( .A(n6293), .B(n6026), .ZN(n6027) );
  NAND2_X2 U6454 ( .A1(n4215), .A2(n6027), .ZN(n6287) );
  INV_X4 U6455 ( .A(n6288), .ZN(n6028) );
  XNOR2_X2 U6456 ( .A(n6289), .B(n6028), .ZN(n7242) );
  MUX2_X2 U6457 ( .A(n4493), .B(n7242), .S(n4078), .Z(n6029) );
  NAND2_X2 U6458 ( .A1(n4166), .A2(n4493), .ZN(n6282) );
  INV_X4 U6459 ( .A(n6283), .ZN(n7486) );
  INV_X4 U6460 ( .A(iAddr[16]), .ZN(n6033) );
  NAND2_X2 U6461 ( .A1(n6033), .A2(n6032), .ZN(n7999) );
  INV_X4 U6462 ( .A(iAddr[18]), .ZN(n6036) );
  NAND2_X2 U6463 ( .A1(n6036), .A2(n6035), .ZN(n8007) );
  AOI22_X2 U6464 ( .A1(n6039), .A2(n8019), .B1(n7427), .B2(n7962), .ZN(n6044)
         );
  NAND2_X2 U6465 ( .A1(n7219), .A2(n7295), .ZN(n6043) );
  AOI22_X2 U6466 ( .A1(n8020), .A2(n7663), .B1(n6040), .B2(n7291), .ZN(n6042)
         );
  NAND2_X2 U6467 ( .A1(n7209), .A2(n7921), .ZN(n6041) );
  NAND4_X2 U6468 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n7441)
         );
  MUX2_X2 U6469 ( .A(n7566), .B(n6045), .S(n4078), .Z(n7442) );
  AOI211_X2 U6470 ( .C1(n7507), .C2(n7441), .A(n6047), .B(n4585), .ZN(n8017)
         );
  INV_X4 U6471 ( .A(n8477), .ZN(n7562) );
  INV_X4 U6472 ( .A(iAddr[6]), .ZN(n6053) );
  NAND2_X2 U6473 ( .A1(n6053), .A2(n6052), .ZN(n8041) );
  INV_X4 U6474 ( .A(iAddr[8]), .ZN(n6056) );
  NAND2_X2 U6475 ( .A1(n6056), .A2(n6055), .ZN(n8053) );
  INV_X4 U6476 ( .A(iAddr[10]), .ZN(n6059) );
  NAND2_X2 U6477 ( .A1(n6059), .A2(n6058), .ZN(n8065) );
  INV_X4 U6478 ( .A(iAddr[12]), .ZN(n6062) );
  NAND2_X2 U6479 ( .A1(n6062), .A2(n6061), .ZN(n8077) );
  INV_X4 U6480 ( .A(iAddr[14]), .ZN(n6065) );
  NAND2_X2 U6481 ( .A1(n6065), .A2(n6064), .ZN(n8088) );
  NAND2_X2 U6482 ( .A1(n4745), .A2(n4359), .ZN(n6066) );
  OAI221_X2 U6483 ( .B1(n8665), .B2(n7123), .C1(n8195), .C2(n4755), .A(n6066), 
        .ZN(iAddr[31]) );
  INV_X4 U6484 ( .A(iAddr[30]), .ZN(n6068) );
  XNOR2_X2 U6485 ( .A(n6069), .B(iAddr[31]), .ZN(n8120) );
  NAND2_X2 U6486 ( .A1(n4416), .A2(n4750), .ZN(n6075) );
  MUX2_X2 U6487 ( .A(n6075), .B(n6074), .S(n7547), .Z(n6076) );
  NAND2_X2 U6488 ( .A1(n6077), .A2(n6076), .ZN(n8300) );
  NAND2_X2 U6489 ( .A1(n4099), .A2(n8304), .ZN(n8303) );
  NAND2_X2 U6490 ( .A1(n4080), .A2(n4418), .ZN(n6082) );
  NAND2_X2 U6491 ( .A1(n4746), .A2(memAddr[15]), .ZN(n6081) );
  NAND2_X2 U6492 ( .A1(regWrData[15]), .A2(n4748), .ZN(n6080) );
  INV_X4 U6493 ( .A(n6169), .ZN(n6090) );
  NAND2_X2 U6494 ( .A1(n7726), .A2(n4753), .ZN(n6086) );
  INV_X4 U6495 ( .A(n6086), .ZN(n6087) );
  NAND2_X2 U6496 ( .A1(n4394), .A2(n7641), .ZN(n6089) );
  NAND2_X2 U6497 ( .A1(n6088), .A2(n6089), .ZN(n6168) );
  INV_X4 U6498 ( .A(n6091), .ZN(n6175) );
  INV_X4 U6499 ( .A(n7726), .ZN(n7485) );
  NAND2_X2 U6500 ( .A1(n4754), .A2(n7485), .ZN(n6094) );
  NAND2_X2 U6501 ( .A1(n4394), .A2(n8460), .ZN(n6095) );
  OAI21_X4 U6502 ( .B1(n6175), .B2(n6174), .A(n6095), .ZN(n6180) );
  INV_X4 U6503 ( .A(n6180), .ZN(n6100) );
  NAND2_X2 U6504 ( .A1(n7895), .A2(n4753), .ZN(n6096) );
  INV_X4 U6505 ( .A(n6096), .ZN(n6097) );
  NAND2_X2 U6506 ( .A1(n4396), .A2(n8460), .ZN(n6099) );
  NAND2_X2 U6507 ( .A1(n6098), .A2(n6099), .ZN(n6179) );
  INV_X4 U6508 ( .A(n6101), .ZN(n6185) );
  NAND2_X2 U6509 ( .A1(n4754), .A2(n7496), .ZN(n6104) );
  NAND2_X2 U6510 ( .A1(n4396), .A2(n8448), .ZN(n6105) );
  INV_X4 U6511 ( .A(n6191), .ZN(n6110) );
  NAND2_X2 U6512 ( .A1(n8349), .A2(n4753), .ZN(n6106) );
  INV_X4 U6513 ( .A(n6106), .ZN(n6107) );
  NAND2_X2 U6514 ( .A1(n4445), .A2(n8448), .ZN(n6109) );
  NAND2_X2 U6515 ( .A1(n6108), .A2(n6109), .ZN(n6190) );
  INV_X4 U6516 ( .A(n6111), .ZN(n6196) );
  NAND2_X2 U6517 ( .A1(n4754), .A2(n7497), .ZN(n6114) );
  NAND2_X2 U6518 ( .A1(n4445), .A2(n8348), .ZN(n6115) );
  INV_X4 U6519 ( .A(n6202), .ZN(n6119) );
  NAND2_X2 U6520 ( .A1(n8336), .A2(n4753), .ZN(n6116) );
  INV_X4 U6521 ( .A(n6116), .ZN(n6121) );
  NAND2_X2 U6522 ( .A1(n6118), .A2(n6117), .ZN(n6201) );
  INV_X4 U6523 ( .A(n6120), .ZN(n6207) );
  NAND2_X2 U6524 ( .A1(n4752), .A2(n7529), .ZN(n6124) );
  INV_X4 U6525 ( .A(n6213), .ZN(n6130) );
  NAND2_X2 U6526 ( .A1(n4750), .A2(n8364), .ZN(n6126) );
  NAND2_X2 U6527 ( .A1(n4753), .A2(n8326), .ZN(n6127) );
  NAND2_X2 U6528 ( .A1(n6126), .A2(n6127), .ZN(n6128) );
  INV_X4 U6529 ( .A(n6127), .ZN(n6132) );
  NAND2_X2 U6530 ( .A1(n6128), .A2(n6129), .ZN(n6212) );
  INV_X4 U6531 ( .A(n6131), .ZN(n6218) );
  NAND2_X2 U6532 ( .A1(n4754), .A2(n7527), .ZN(n6135) );
  OAI21_X4 U6533 ( .B1(n6218), .B2(n6217), .A(n6136), .ZN(n6224) );
  INV_X4 U6534 ( .A(n6224), .ZN(n6141) );
  NAND2_X2 U6535 ( .A1(n7723), .A2(n4107), .ZN(n6137) );
  NAND2_X2 U6536 ( .A1(n4753), .A2(n7722), .ZN(n6138) );
  NAND2_X2 U6537 ( .A1(n6137), .A2(n6138), .ZN(n6139) );
  INV_X4 U6538 ( .A(n6138), .ZN(n6143) );
  NAND2_X2 U6539 ( .A1(n6139), .A2(n6140), .ZN(n6223) );
  INV_X4 U6540 ( .A(n6142), .ZN(n6229) );
  NAND2_X2 U6541 ( .A1(n4754), .A2(n7501), .ZN(n6146) );
  INV_X4 U6542 ( .A(n6235), .ZN(n6153) );
  NAND2_X2 U6543 ( .A1(n7721), .A2(n4107), .ZN(n6148) );
  NAND2_X2 U6544 ( .A1(n4753), .A2(n7720), .ZN(n6149) );
  NAND2_X2 U6545 ( .A1(n6148), .A2(n6149), .ZN(n6151) );
  INV_X4 U6546 ( .A(n6149), .ZN(n6150) );
  NAND2_X2 U6547 ( .A1(n4446), .A2(n7721), .ZN(n6152) );
  NAND2_X2 U6548 ( .A1(n6151), .A2(n6152), .ZN(n6234) );
  INV_X4 U6549 ( .A(n6154), .ZN(n6240) );
  OAI22_X2 U6550 ( .A1(n4754), .A2(n7504), .B1(n6942), .B2(n4752), .ZN(n6155)
         );
  NAND2_X2 U6551 ( .A1(n4446), .A2(n8316), .ZN(n6156) );
  NAND2_X2 U6552 ( .A1(n6155), .A2(n6156), .ZN(n6239) );
  INV_X4 U6553 ( .A(n6246), .ZN(n6163) );
  NAND2_X2 U6554 ( .A1(n4752), .A2(n7503), .ZN(n6161) );
  NAND2_X2 U6555 ( .A1(n4178), .A2(n4416), .ZN(n8309) );
  NAND2_X2 U6556 ( .A1(n8316), .A2(n4099), .ZN(n8312) );
  INV_X4 U6557 ( .A(n8312), .ZN(n6164) );
  XNOR2_X2 U6558 ( .A(n8311), .B(n6164), .ZN(n7246) );
  INV_X4 U6559 ( .A(n6308), .ZN(n6172) );
  XNOR2_X2 U6560 ( .A(n6169), .B(n6168), .ZN(n6170) );
  NAND2_X2 U6561 ( .A1(n4149), .A2(n6170), .ZN(n6171) );
  INV_X4 U6562 ( .A(n6173), .ZN(n6367) );
  INV_X4 U6563 ( .A(n6174), .ZN(n6176) );
  XNOR2_X2 U6564 ( .A(n6176), .B(n6175), .ZN(n6177) );
  NAND2_X2 U6565 ( .A1(n4210), .A2(n6177), .ZN(n6178) );
  OAI21_X4 U6566 ( .B1(n6367), .B2(n6366), .A(n6178), .ZN(n6406) );
  INV_X4 U6567 ( .A(n6406), .ZN(n6183) );
  XNOR2_X2 U6568 ( .A(n6180), .B(n6179), .ZN(n6181) );
  NAND2_X2 U6569 ( .A1(n4211), .A2(n6181), .ZN(n6182) );
  OAI21_X4 U6570 ( .B1(n6183), .B2(n6405), .A(n6182), .ZN(n6432) );
  INV_X4 U6571 ( .A(n6432), .ZN(n6189) );
  INV_X4 U6572 ( .A(n6184), .ZN(n6186) );
  XNOR2_X2 U6573 ( .A(n6186), .B(n6185), .ZN(n6187) );
  NAND2_X2 U6574 ( .A1(n4110), .A2(n6187), .ZN(n6188) );
  INV_X4 U6575 ( .A(n6460), .ZN(n6194) );
  XNOR2_X2 U6576 ( .A(n6191), .B(n6190), .ZN(n6192) );
  NAND2_X2 U6577 ( .A1(n4111), .A2(n6192), .ZN(n6193) );
  OAI21_X4 U6578 ( .B1(n6194), .B2(n6459), .A(n6193), .ZN(n6485) );
  INV_X4 U6579 ( .A(n6485), .ZN(n6200) );
  INV_X4 U6580 ( .A(n6195), .ZN(n6197) );
  XNOR2_X2 U6581 ( .A(n6197), .B(n6196), .ZN(n6198) );
  NAND2_X2 U6582 ( .A1(n4112), .A2(n6198), .ZN(n6199) );
  OAI21_X4 U6583 ( .B1(n6200), .B2(n6484), .A(n6199), .ZN(n6515) );
  INV_X4 U6584 ( .A(n6515), .ZN(n6205) );
  XNOR2_X2 U6585 ( .A(n6202), .B(n6201), .ZN(n6203) );
  NAND2_X2 U6586 ( .A1(n4113), .A2(n6203), .ZN(n6204) );
  INV_X4 U6587 ( .A(n6740), .ZN(n6211) );
  INV_X4 U6588 ( .A(n6206), .ZN(n6208) );
  XNOR2_X2 U6589 ( .A(n6208), .B(n6207), .ZN(n6209) );
  NAND2_X2 U6590 ( .A1(n4114), .A2(n6209), .ZN(n6210) );
  OAI21_X4 U6591 ( .B1(n6211), .B2(n6739), .A(n6210), .ZN(n6765) );
  INV_X4 U6592 ( .A(n6765), .ZN(n6216) );
  XNOR2_X2 U6593 ( .A(n6213), .B(n6212), .ZN(n6214) );
  NAND2_X2 U6594 ( .A1(n4212), .A2(n6214), .ZN(n6215) );
  INV_X4 U6595 ( .A(n6786), .ZN(n6222) );
  INV_X4 U6596 ( .A(n6217), .ZN(n6219) );
  XNOR2_X2 U6597 ( .A(n6219), .B(n6218), .ZN(n6220) );
  NAND2_X2 U6598 ( .A1(n4183), .A2(n6220), .ZN(n6221) );
  OAI21_X4 U6599 ( .B1(n6222), .B2(n6785), .A(n6221), .ZN(n6818) );
  INV_X4 U6600 ( .A(n6818), .ZN(n6227) );
  XNOR2_X2 U6601 ( .A(n6224), .B(n6223), .ZN(n6225) );
  NAND2_X2 U6602 ( .A1(n4184), .A2(n6225), .ZN(n6226) );
  INV_X4 U6603 ( .A(n6829), .ZN(n6233) );
  INV_X4 U6604 ( .A(n6228), .ZN(n6230) );
  XNOR2_X2 U6605 ( .A(n6230), .B(n6229), .ZN(n6231) );
  NAND2_X2 U6606 ( .A1(n4115), .A2(n6231), .ZN(n6232) );
  OAI21_X4 U6607 ( .B1(n6233), .B2(n6828), .A(n6232), .ZN(n6871) );
  INV_X4 U6608 ( .A(n6871), .ZN(n6238) );
  XNOR2_X2 U6609 ( .A(n6235), .B(n6234), .ZN(n6236) );
  NAND2_X2 U6610 ( .A1(n4185), .A2(n6236), .ZN(n6237) );
  INV_X4 U6611 ( .A(n6996), .ZN(n6244) );
  INV_X4 U6612 ( .A(n6239), .ZN(n6241) );
  XNOR2_X2 U6613 ( .A(n6241), .B(n6240), .ZN(n6242) );
  NAND2_X2 U6614 ( .A1(n4213), .A2(n6242), .ZN(n6243) );
  OAI21_X4 U6615 ( .B1(n6244), .B2(n6995), .A(n6243), .ZN(n7035) );
  INV_X4 U6616 ( .A(n7035), .ZN(n6249) );
  XNOR2_X2 U6617 ( .A(n6246), .B(n6245), .ZN(n6247) );
  NAND2_X2 U6618 ( .A1(n4186), .A2(n6247), .ZN(n6248) );
  NAND2_X2 U6619 ( .A1(n7246), .A2(n7245), .ZN(n8313) );
  NAND2_X2 U6620 ( .A1(n4084), .A2(n8316), .ZN(n8314) );
  INV_X4 U6621 ( .A(n7723), .ZN(n7500) );
  NAND2_X2 U6622 ( .A1(n4312), .A2(n6250), .ZN(n6262) );
  OAI22_X2 U6623 ( .A1(n8407), .A2(n5182), .B1(n8486), .B2(n7528), .ZN(n6256)
         );
  NAND2_X2 U6624 ( .A1(n7212), .A2(n8502), .ZN(n6253) );
  NAND2_X2 U6625 ( .A1(n6251), .A2(n8019), .ZN(n6252) );
  INV_X4 U6626 ( .A(n4317), .ZN(n6254) );
  NAND2_X2 U6627 ( .A1(n6258), .A2(n6257), .ZN(n6260) );
  NAND2_X2 U6628 ( .A1(n8503), .A2(n4735), .ZN(n6259) );
  NAND4_X2 U6629 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .ZN(n7396)
         );
  INV_X4 U6630 ( .A(n7396), .ZN(n6264) );
  MUX2_X2 U6631 ( .A(n8333), .B(n6263), .S(n6254), .Z(n7429) );
  OAI22_X2 U6632 ( .A1(n8324), .A2(n6264), .B1(n8323), .B2(n7429), .ZN(n8322)
         );
  INV_X4 U6633 ( .A(n7278), .ZN(n6265) );
  OAI22_X2 U6634 ( .A1(n8323), .A2(n7207), .B1(n8324), .B2(n6265), .ZN(n8332)
         );
  INV_X4 U6635 ( .A(n6266), .ZN(n7544) );
  INV_X4 U6636 ( .A(n7291), .ZN(n8022) );
  INV_X4 U6637 ( .A(n6267), .ZN(n7535) );
  INV_X4 U6638 ( .A(n7971), .ZN(n7917) );
  INV_X4 U6639 ( .A(n6268), .ZN(n7543) );
  INV_X4 U6640 ( .A(n7980), .ZN(n7967) );
  INV_X4 U6641 ( .A(n6269), .ZN(n7517) );
  INV_X4 U6642 ( .A(n7675), .ZN(n7976) );
  INV_X4 U6643 ( .A(n6270), .ZN(n7522) );
  INV_X4 U6644 ( .A(n7676), .ZN(n8377) );
  INV_X4 U6645 ( .A(n7913), .ZN(n7669) );
  INV_X4 U6646 ( .A(n6271), .ZN(n7510) );
  INV_X4 U6647 ( .A(n6272), .ZN(n7511) );
  INV_X4 U6648 ( .A(n6273), .ZN(n7534) );
  INV_X4 U6649 ( .A(n7686), .ZN(n7705) );
  INV_X4 U6650 ( .A(n8420), .ZN(n8419) );
  INV_X4 U6651 ( .A(n6274), .ZN(n7542) );
  INV_X4 U6652 ( .A(n8408), .ZN(n8429) );
  INV_X4 U6653 ( .A(n6275), .ZN(n7533) );
  INV_X4 U6654 ( .A(n7695), .ZN(n8433) );
  INV_X4 U6655 ( .A(n8407), .ZN(n7560) );
  INV_X4 U6656 ( .A(n8447), .ZN(n7561) );
  INV_X4 U6657 ( .A(n6276), .ZN(n7519) );
  AOI22_X2 U6658 ( .A1(n8430), .A2(n4735), .B1(n8404), .B2(n6254), .ZN(n6280)
         );
  NAND2_X2 U6659 ( .A1(n6281), .A2(n6280), .ZN(n8462) );
  INV_X4 U6660 ( .A(n7991), .ZN(n6284) );
  INV_X4 U6661 ( .A(n6285), .ZN(n8463) );
  INV_X4 U6662 ( .A(n6286), .ZN(n7360) );
  INV_X4 U6663 ( .A(n6290), .ZN(n6363) );
  INV_X4 U6664 ( .A(n6294), .ZN(n6390) );
  INV_X4 U6665 ( .A(n6298), .ZN(n6384) );
  INV_X4 U6666 ( .A(n6302), .ZN(n6378) );
  INV_X4 U6667 ( .A(n6306), .ZN(n6372) );
  XNOR2_X2 U6668 ( .A(n6308), .B(n6307), .ZN(n6309) );
  NAND2_X2 U6669 ( .A1(n4233), .A2(n6309), .ZN(n6370) );
  INV_X4 U6670 ( .A(n6371), .ZN(n6310) );
  XNOR2_X2 U6671 ( .A(n6372), .B(n6310), .ZN(n6311) );
  NAND2_X2 U6672 ( .A1(n4188), .A2(n6311), .ZN(n6376) );
  INV_X4 U6673 ( .A(n6377), .ZN(n6312) );
  XNOR2_X2 U6674 ( .A(n6378), .B(n6312), .ZN(n6313) );
  NAND2_X2 U6675 ( .A1(n4181), .A2(n6313), .ZN(n6382) );
  INV_X4 U6676 ( .A(n6383), .ZN(n6314) );
  XNOR2_X2 U6677 ( .A(n6384), .B(n6314), .ZN(n6315) );
  NAND2_X2 U6678 ( .A1(n4204), .A2(n6315), .ZN(n6388) );
  INV_X4 U6679 ( .A(n6389), .ZN(n6316) );
  XNOR2_X2 U6680 ( .A(n6390), .B(n6316), .ZN(n6317) );
  NAND2_X2 U6681 ( .A1(n4229), .A2(n6317), .ZN(n6361) );
  INV_X4 U6682 ( .A(n6362), .ZN(n6318) );
  XNOR2_X2 U6683 ( .A(n6363), .B(n6318), .ZN(n7363) );
  MUX2_X2 U6684 ( .A(n4580), .B(n7363), .S(n4078), .Z(n6319) );
  NAND2_X2 U6685 ( .A1(n4162), .A2(n4580), .ZN(n6530) );
  INV_X4 U6686 ( .A(n7663), .ZN(n7516) );
  INV_X4 U6687 ( .A(n8486), .ZN(n7559) );
  INV_X4 U6688 ( .A(n8502), .ZN(n8485) );
  INV_X4 U6689 ( .A(n8458), .ZN(n7521) );
  INV_X4 U6690 ( .A(n7381), .ZN(n7509) );
  XNOR2_X2 U6691 ( .A(n7381), .B(n7379), .ZN(n8524) );
  INV_X4 U6692 ( .A(n8524), .ZN(n8317) );
  INV_X4 U6693 ( .A(n8018), .ZN(n7662) );
  XNOR2_X2 U6694 ( .A(n8536), .B(n6320), .ZN(n6325) );
  INV_X4 U6695 ( .A(n6325), .ZN(n6321) );
  XNOR2_X2 U6696 ( .A(n7192), .B(n6321), .ZN(n6327) );
  INV_X4 U6697 ( .A(n6327), .ZN(n8595) );
  INV_X4 U6698 ( .A(n6322), .ZN(n6323) );
  XNOR2_X2 U6699 ( .A(n8605), .B(n6323), .ZN(n6324) );
  XNOR2_X2 U6700 ( .A(n6324), .B(n4737), .ZN(n7484) );
  NAND2_X2 U6701 ( .A1(n8544), .A2(n7484), .ZN(n8545) );
  INV_X4 U6702 ( .A(n8594), .ZN(n6328) );
  NAND2_X2 U6703 ( .A1(n6325), .A2(n6365), .ZN(n6326) );
  INV_X4 U6704 ( .A(n8643), .ZN(n7555) );
  INV_X4 U6705 ( .A(n7658), .ZN(n7557) );
  INV_X4 U6706 ( .A(n7616), .ZN(n7556) );
  XNOR2_X2 U6707 ( .A(n8604), .B(n8317), .ZN(n7399) );
  INV_X4 U6708 ( .A(n7399), .ZN(n8318) );
  INV_X4 U6709 ( .A(n7721), .ZN(n7502) );
  INV_X4 U6710 ( .A(n8335), .ZN(n7545) );
  INV_X4 U6711 ( .A(iAddr[2]), .ZN(n6694) );
  MUX2_X2 U6712 ( .A(n4556), .B(n6694), .S(n4793), .Z(n3524) );
  OAI22_X2 U6713 ( .A1(n8761), .A2(n6332), .B1(n7882), .B2(n6331), .ZN(n7112)
         );
  OAI22_X2 U6714 ( .A1(n7666), .A2(n7113), .B1(n8871), .B2(n4124), .ZN(n9196)
         );
  OAI22_X2 U6715 ( .A1(n8816), .A2(n6332), .B1(n7862), .B2(n6331), .ZN(n7121)
         );
  OAI22_X2 U6716 ( .A1(n7666), .A2(n7122), .B1(n8902), .B2(n4124), .ZN(n9195)
         );
  NAND2_X2 U6717 ( .A1(n6333), .A2(n6338), .ZN(n6337) );
  NAND2_X2 U6718 ( .A1(not_trap_2), .A2(n4792), .ZN(n6334) );
  OAI211_X2 U6719 ( .C1(n4772), .C2(n4716), .A(n6337), .B(n6334), .ZN(n3667)
         );
  NAND2_X2 U6720 ( .A1(n4791), .A2(n4726), .ZN(n6335) );
  OAI211_X2 U6721 ( .C1(n7589), .C2(n4772), .A(n6337), .B(n6335), .ZN(n3686)
         );
  NAND2_X2 U6722 ( .A1(n4791), .A2(n4725), .ZN(n6336) );
  OAI211_X2 U6723 ( .C1(n7591), .C2(n4772), .A(n6337), .B(n6336), .ZN(n3690)
         );
  OAI221_X2 U6724 ( .B1(n7593), .B2(n4772), .C1(n7594), .C2(n4787), .A(n6337), 
        .ZN(n3694) );
  MUX2_X2 U6725 ( .A(n4106), .B(n4627), .S(n4796), .Z(n3762) );
  NAND2_X2 U6726 ( .A1(instruction[4]), .A2(n4806), .ZN(n6340) );
  NAND2_X2 U6727 ( .A1(n4129), .A2(n4811), .ZN(n6339) );
  NAND2_X2 U6728 ( .A1(instruction[2]), .A2(n4806), .ZN(n6342) );
  NAND2_X2 U6729 ( .A1(n4539), .A2(n4811), .ZN(n6341) );
  NAND2_X2 U6730 ( .A1(n4321), .A2(n4811), .ZN(n6344) );
  NAND2_X2 U6731 ( .A1(instruction[0]), .A2(n4806), .ZN(n6343) );
  NAND2_X2 U6732 ( .A1(n4762), .A2(regWrData[15]), .ZN(n6348) );
  NAND2_X2 U6733 ( .A1(n4759), .A2(memAddr[15]), .ZN(n6347) );
  NAND2_X2 U6734 ( .A1(n4781), .A2(n4683), .ZN(n6346) );
  NAND2_X2 U6735 ( .A1(n8173), .A2(n4792), .ZN(n7164) );
  NAND2_X2 U6736 ( .A1(n4757), .A2(n4652), .ZN(n6345) );
  NAND4_X2 U6737 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n3372)
         );
  NAND2_X2 U6738 ( .A1(n4762), .A2(regWrData[10]), .ZN(n6352) );
  NAND2_X2 U6739 ( .A1(n4759), .A2(memAddr[10]), .ZN(n6351) );
  NAND2_X2 U6740 ( .A1(n4779), .A2(n4684), .ZN(n6350) );
  NAND2_X2 U6741 ( .A1(n4757), .A2(n4704), .ZN(n6349) );
  NAND4_X2 U6742 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n3373)
         );
  NAND2_X2 U6743 ( .A1(n4762), .A2(regWrData[20]), .ZN(n6356) );
  NAND2_X2 U6744 ( .A1(n4759), .A2(memAddr[20]), .ZN(n6355) );
  NAND2_X2 U6745 ( .A1(n4779), .A2(n4685), .ZN(n6354) );
  NAND2_X2 U6746 ( .A1(n4757), .A2(n4653), .ZN(n6353) );
  NAND4_X2 U6747 ( .A1(n6356), .A2(n6355), .A3(n6354), .A4(n6353), .ZN(n3374)
         );
  OAI22_X2 U6748 ( .A1(n8916), .A2(n4789), .B1(n8650), .B2(n4772), .ZN(n3375)
         );
  OAI22_X2 U6749 ( .A1(n8651), .A2(n4789), .B1(n8849), .B2(n4783), .ZN(n3376)
         );
  OAI22_X2 U6750 ( .A1(n8652), .A2(n4789), .B1(n8848), .B2(n4783), .ZN(n3378)
         );
  NAND2_X2 U6751 ( .A1(n4762), .A2(regWrData[21]), .ZN(n6360) );
  NAND2_X2 U6752 ( .A1(memAddr[21]), .A2(n4758), .ZN(n6359) );
  NAND2_X2 U6753 ( .A1(n4779), .A2(n4686), .ZN(n6358) );
  NAND2_X2 U6754 ( .A1(n4757), .A2(n4705), .ZN(n6357) );
  NAND4_X2 U6755 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(n3381)
         );
  INV_X4 U6756 ( .A(n6364), .ZN(n6532) );
  INV_X4 U6757 ( .A(n6366), .ZN(n6368) );
  XNOR2_X2 U6758 ( .A(n6368), .B(n6367), .ZN(n6369) );
  NAND2_X2 U6759 ( .A1(n4235), .A2(n6369), .ZN(n6402) );
  INV_X4 U6760 ( .A(n6403), .ZN(n6374) );
  OAI21_X4 U6761 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6373) );
  INV_X4 U6762 ( .A(n6373), .ZN(n6404) );
  XNOR2_X2 U6763 ( .A(n6374), .B(n6404), .ZN(n6375) );
  NAND2_X2 U6764 ( .A1(n4234), .A2(n6375), .ZN(n6399) );
  INV_X4 U6765 ( .A(n6400), .ZN(n6380) );
  INV_X4 U6766 ( .A(n6379), .ZN(n6401) );
  XNOR2_X2 U6767 ( .A(n6380), .B(n6401), .ZN(n6381) );
  NAND2_X2 U6768 ( .A1(n4189), .A2(n6381), .ZN(n6396) );
  INV_X4 U6769 ( .A(n6397), .ZN(n6386) );
  OAI21_X4 U6770 ( .B1(n6384), .B2(n6383), .A(n6382), .ZN(n6385) );
  INV_X4 U6771 ( .A(n6385), .ZN(n6398) );
  XNOR2_X2 U6772 ( .A(n6386), .B(n6398), .ZN(n6387) );
  NAND2_X2 U6773 ( .A1(n4182), .A2(n6387), .ZN(n6411) );
  INV_X4 U6774 ( .A(n6412), .ZN(n6392) );
  OAI21_X4 U6775 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6391) );
  INV_X4 U6776 ( .A(n6391), .ZN(n6413) );
  XNOR2_X2 U6777 ( .A(n6392), .B(n6413), .ZN(n6393) );
  NAND2_X2 U6778 ( .A1(n4262), .A2(n6393), .ZN(n6394) );
  INV_X4 U6779 ( .A(n6395), .ZN(n6541) );
  XNOR2_X2 U6780 ( .A(n6406), .B(n6405), .ZN(n6407) );
  NAND2_X2 U6781 ( .A1(n4230), .A2(n6407), .ZN(n6428) );
  XNOR2_X2 U6782 ( .A(n6427), .B(n6429), .ZN(n6408) );
  NAND2_X2 U6783 ( .A1(n4236), .A2(n6408), .ZN(n6424) );
  XNOR2_X2 U6784 ( .A(n6423), .B(n6425), .ZN(n6409) );
  NAND2_X2 U6785 ( .A1(n4218), .A2(n6409), .ZN(n6420) );
  XNOR2_X2 U6786 ( .A(n6419), .B(n6421), .ZN(n6410) );
  NAND2_X2 U6787 ( .A1(n4190), .A2(n6410), .ZN(n6437) );
  INV_X4 U6788 ( .A(n6438), .ZN(n6415) );
  OAI21_X4 U6789 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(n6414) );
  INV_X4 U6790 ( .A(n6414), .ZN(n6439) );
  XNOR2_X2 U6791 ( .A(n6415), .B(n6439), .ZN(n6416) );
  NAND2_X2 U6792 ( .A1(n4281), .A2(n6416), .ZN(n6417) );
  INV_X4 U6793 ( .A(n6418), .ZN(n6550) );
  INV_X4 U6794 ( .A(n6419), .ZN(n6422) );
  OAI21_X4 U6795 ( .B1(n6422), .B2(n6421), .A(n6420), .ZN(n6447) );
  INV_X4 U6796 ( .A(n6423), .ZN(n6426) );
  OAI21_X4 U6797 ( .B1(n6426), .B2(n6425), .A(n6424), .ZN(n6451) );
  INV_X4 U6798 ( .A(n6427), .ZN(n6430) );
  OAI21_X4 U6799 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6455) );
  XNOR2_X2 U6800 ( .A(n6432), .B(n6431), .ZN(n6433) );
  NAND2_X2 U6801 ( .A1(n4237), .A2(n6433), .ZN(n6456) );
  XNOR2_X2 U6802 ( .A(n6455), .B(n6457), .ZN(n6434) );
  NAND2_X2 U6803 ( .A1(n4231), .A2(n6434), .ZN(n6452) );
  XNOR2_X2 U6804 ( .A(n6451), .B(n6453), .ZN(n6435) );
  NAND2_X2 U6805 ( .A1(n4219), .A2(n6435), .ZN(n6448) );
  XNOR2_X2 U6806 ( .A(n6447), .B(n6449), .ZN(n6436) );
  NAND2_X2 U6807 ( .A1(n4225), .A2(n6436), .ZN(n6444) );
  INV_X4 U6808 ( .A(n6445), .ZN(n6441) );
  INV_X4 U6809 ( .A(n6440), .ZN(n6446) );
  XNOR2_X2 U6810 ( .A(n6441), .B(n6446), .ZN(n6442) );
  NAND2_X2 U6811 ( .A1(n4282), .A2(n6442), .ZN(n6443) );
  INV_X4 U6812 ( .A(n6559), .ZN(n6467) );
  INV_X4 U6813 ( .A(n6447), .ZN(n6450) );
  INV_X4 U6814 ( .A(n6451), .ZN(n6454) );
  INV_X4 U6815 ( .A(n6455), .ZN(n6458) );
  XNOR2_X2 U6816 ( .A(n6460), .B(n6459), .ZN(n6461) );
  NAND2_X2 U6817 ( .A1(n4239), .A2(n6461), .ZN(n6481) );
  XNOR2_X2 U6818 ( .A(n6480), .B(n6482), .ZN(n6462) );
  NAND2_X2 U6819 ( .A1(n4238), .A2(n6462), .ZN(n6477) );
  XNOR2_X2 U6820 ( .A(n6476), .B(n6478), .ZN(n6463) );
  NAND2_X2 U6821 ( .A1(n4220), .A2(n6463), .ZN(n6473) );
  XNOR2_X2 U6822 ( .A(n6472), .B(n6474), .ZN(n6464) );
  NAND2_X2 U6823 ( .A1(n4226), .A2(n6464), .ZN(n6469) );
  XNOR2_X2 U6824 ( .A(n6468), .B(n6470), .ZN(n6465) );
  NAND2_X2 U6825 ( .A1(n4298), .A2(n6465), .ZN(n6466) );
  INV_X4 U6826 ( .A(n6567), .ZN(n6492) );
  INV_X4 U6827 ( .A(n6468), .ZN(n6471) );
  OAI21_X4 U6828 ( .B1(n6471), .B2(n6470), .A(n6469), .ZN(n6494) );
  INV_X4 U6829 ( .A(n6472), .ZN(n6475) );
  OAI21_X4 U6830 ( .B1(n6475), .B2(n6474), .A(n6473), .ZN(n6499) );
  INV_X4 U6831 ( .A(n6476), .ZN(n6479) );
  OAI21_X4 U6832 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6504) );
  INV_X4 U6833 ( .A(n6480), .ZN(n6483) );
  OAI21_X4 U6834 ( .B1(n6483), .B2(n6482), .A(n6481), .ZN(n6509) );
  XNOR2_X2 U6835 ( .A(n6485), .B(n6484), .ZN(n6486) );
  NAND2_X2 U6836 ( .A1(n4252), .A2(n6486), .ZN(n6510) );
  XNOR2_X2 U6837 ( .A(n6509), .B(n6511), .ZN(n6487) );
  NAND2_X2 U6838 ( .A1(n4240), .A2(n6487), .ZN(n6505) );
  XNOR2_X2 U6839 ( .A(n6504), .B(n6506), .ZN(n6488) );
  NAND2_X2 U6840 ( .A1(n4221), .A2(n6488), .ZN(n6500) );
  XNOR2_X2 U6841 ( .A(n6499), .B(n6501), .ZN(n6489) );
  NAND2_X2 U6842 ( .A1(n4227), .A2(n6489), .ZN(n6495) );
  XNOR2_X2 U6843 ( .A(n6494), .B(n6496), .ZN(n6490) );
  NAND2_X2 U6844 ( .A1(n4299), .A2(n6490), .ZN(n6491) );
  INV_X4 U6845 ( .A(n6493), .ZN(n6726) );
  INV_X4 U6846 ( .A(n6494), .ZN(n6497) );
  INV_X4 U6847 ( .A(n6498), .ZN(n6729) );
  INV_X4 U6848 ( .A(n6499), .ZN(n6502) );
  INV_X4 U6849 ( .A(n6503), .ZN(n6732) );
  INV_X4 U6850 ( .A(n6504), .ZN(n6507) );
  INV_X4 U6851 ( .A(n6508), .ZN(n6735) );
  INV_X4 U6852 ( .A(n6509), .ZN(n6512) );
  INV_X4 U6853 ( .A(n6513), .ZN(n6738) );
  XNOR2_X2 U6854 ( .A(n6515), .B(n6514), .ZN(n6516) );
  NAND2_X2 U6855 ( .A1(n4243), .A2(n6516), .ZN(n6736) );
  INV_X4 U6856 ( .A(n6737), .ZN(n6517) );
  XNOR2_X2 U6857 ( .A(n6738), .B(n6517), .ZN(n6518) );
  NAND2_X2 U6858 ( .A1(n4253), .A2(n6518), .ZN(n6733) );
  INV_X4 U6859 ( .A(n6734), .ZN(n6519) );
  XNOR2_X2 U6860 ( .A(n6735), .B(n6519), .ZN(n6520) );
  NAND2_X2 U6861 ( .A1(n4222), .A2(n6520), .ZN(n6730) );
  INV_X4 U6862 ( .A(n6731), .ZN(n6521) );
  XNOR2_X2 U6863 ( .A(n6732), .B(n6521), .ZN(n6522) );
  NAND2_X2 U6864 ( .A1(n4289), .A2(n6522), .ZN(n6727) );
  INV_X4 U6865 ( .A(n6728), .ZN(n6523) );
  XNOR2_X2 U6866 ( .A(n6729), .B(n6523), .ZN(n6524) );
  NAND2_X2 U6867 ( .A1(n4296), .A2(n6524), .ZN(n6724) );
  INV_X4 U6868 ( .A(n6725), .ZN(n6525) );
  XNOR2_X2 U6869 ( .A(n6726), .B(n6525), .ZN(n7044) );
  MUX2_X2 U6870 ( .A(n4581), .B(n7044), .S(n4078), .Z(n6529) );
  INV_X4 U6871 ( .A(n7045), .ZN(n6527) );
  NAND2_X2 U6872 ( .A1(n7243), .A2(n7046), .ZN(n6526) );
  NAND2_X2 U6873 ( .A1(n6528), .A2(n4581), .ZN(n6900) );
  INV_X4 U6874 ( .A(n7227), .ZN(n6539) );
  INV_X4 U6875 ( .A(n6531), .ZN(n6533) );
  XNOR2_X2 U6876 ( .A(n6533), .B(n6532), .ZN(n6894) );
  INV_X4 U6877 ( .A(n6894), .ZN(n6536) );
  INV_X4 U6878 ( .A(n6892), .ZN(n6534) );
  NAND2_X2 U6879 ( .A1(n7273), .A2(n6534), .ZN(n6535) );
  OAI221_X2 U6880 ( .B1(n6897), .B2(n7362), .C1(n6536), .C2(n4784), .A(n6535), 
        .ZN(n6537) );
  OAI21_X4 U6881 ( .B1(n6539), .B2(n7226), .A(n6538), .ZN(n7080) );
  INV_X4 U6882 ( .A(n7080), .ZN(n6548) );
  INV_X4 U6883 ( .A(n6540), .ZN(n6542) );
  XNOR2_X2 U6884 ( .A(n6542), .B(n6541), .ZN(n6925) );
  INV_X4 U6885 ( .A(n6925), .ZN(n6545) );
  NAND2_X2 U6886 ( .A1(n7243), .A2(n4205), .ZN(n6544) );
  NAND2_X2 U6887 ( .A1(n7273), .A2(n6924), .ZN(n6543) );
  OAI211_X2 U6888 ( .C1(n6545), .C2(n4784), .A(n6544), .B(n6543), .ZN(n6546)
         );
  NAND3_X2 U6889 ( .A1(n6546), .A2(n4784), .A3(n4570), .ZN(n6547) );
  OAI21_X4 U6890 ( .B1(n6548), .B2(n7079), .A(n6547), .ZN(n6955) );
  INV_X4 U6891 ( .A(n6955), .ZN(n6557) );
  INV_X4 U6892 ( .A(n6549), .ZN(n6551) );
  INV_X4 U6893 ( .A(n6934), .ZN(n6552) );
  NAND2_X2 U6894 ( .A1(n6552), .A2(n7243), .ZN(n6553) );
  OAI221_X2 U6895 ( .B1(n6554), .B2(n4169), .C1(n4389), .C2(n4784), .A(n6553), 
        .ZN(n6555) );
  NAND2_X2 U6896 ( .A1(n4306), .A2(n6555), .ZN(n6556) );
  OAI21_X4 U6897 ( .B1(n6557), .B2(n6954), .A(n6556), .ZN(n6709) );
  INV_X4 U6898 ( .A(n6709), .ZN(n6565) );
  XNOR2_X2 U6899 ( .A(n6559), .B(n6558), .ZN(n6882) );
  MUX2_X2 U6900 ( .A(n4582), .B(n6882), .S(n4078), .Z(n6563) );
  INV_X4 U6901 ( .A(n6883), .ZN(n6561) );
  NAND2_X2 U6902 ( .A1(n7243), .A2(n6884), .ZN(n6560) );
  NAND2_X2 U6903 ( .A1(n6562), .A2(n4582), .ZN(n6564) );
  INV_X4 U6904 ( .A(n7199), .ZN(n6574) );
  XNOR2_X2 U6905 ( .A(n6567), .B(n6566), .ZN(n7060) );
  INV_X4 U6906 ( .A(n7060), .ZN(n6570) );
  INV_X4 U6907 ( .A(n7058), .ZN(n6568) );
  NAND2_X2 U6908 ( .A1(n6568), .A2(n7243), .ZN(n6569) );
  OAI221_X2 U6909 ( .B1(n6571), .B2(n4169), .C1(n6570), .C2(n4784), .A(n6569), 
        .ZN(n6572) );
  NAND2_X2 U6910 ( .A1(n4307), .A2(n6572), .ZN(n6573) );
  OAI21_X4 U6911 ( .B1(n6574), .B2(n7198), .A(n6573), .ZN(n6899) );
  XNOR2_X2 U6912 ( .A(n6901), .B(n6899), .ZN(n6577) );
  NAND2_X2 U6913 ( .A1(n7499), .A2(n7412), .ZN(n6575) );
  NAND4_X2 U6914 ( .A1(n8398), .A2(n8397), .A3(n8399), .A4(n6578), .ZN(
        aluRes_2[21]) );
  NAND2_X2 U6915 ( .A1(memAddr[21]), .A2(n4781), .ZN(n6580) );
  NAND2_X2 U6916 ( .A1(aluRes_2[21]), .A2(n4792), .ZN(n6579) );
  NAND2_X2 U6917 ( .A1(n6580), .A2(n6579), .ZN(n9160) );
  NAND2_X2 U6918 ( .A1(n4762), .A2(regWrData[22]), .ZN(n6584) );
  NAND2_X2 U6919 ( .A1(memAddr[22]), .A2(n4759), .ZN(n6583) );
  NAND2_X2 U6920 ( .A1(n4779), .A2(n4687), .ZN(n6582) );
  NAND2_X2 U6921 ( .A1(n4757), .A2(n4706), .ZN(n6581) );
  NAND4_X2 U6922 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n3384)
         );
  AOI22_X2 U6923 ( .A1(n4761), .A2(regWrData[17]), .B1(memAddr[17]), .B2(n4759), .ZN(n6586) );
  AOI22_X2 U6924 ( .A1(n4778), .A2(n4675), .B1(n4757), .B2(n4343), .ZN(n6585)
         );
  NAND2_X2 U6925 ( .A1(n6586), .A2(n6585), .ZN(n3385) );
  NAND2_X2 U6926 ( .A1(n4762), .A2(regWrData[12]), .ZN(n6590) );
  NAND2_X2 U6927 ( .A1(n4759), .A2(memAddr[12]), .ZN(n6589) );
  NAND2_X2 U6928 ( .A1(n4779), .A2(n4688), .ZN(n6588) );
  NAND2_X2 U6929 ( .A1(n4757), .A2(n4707), .ZN(n6587) );
  NAND4_X2 U6930 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n3386)
         );
  NAND2_X2 U6931 ( .A1(n4762), .A2(regWrData[29]), .ZN(n6594) );
  NAND2_X2 U6932 ( .A1(n4759), .A2(memAddr[29]), .ZN(n6593) );
  NAND2_X2 U6933 ( .A1(n4779), .A2(n4689), .ZN(n6592) );
  NAND2_X2 U6934 ( .A1(n4757), .A2(n4654), .ZN(n6591) );
  NAND4_X2 U6935 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n3387)
         );
  AOI22_X2 U6936 ( .A1(n4762), .A2(regWrData[8]), .B1(n4758), .B2(memAddr[8]), 
        .ZN(n6596) );
  AOI22_X2 U6937 ( .A1(n4778), .A2(n4676), .B1(n4757), .B2(n4346), .ZN(n6595)
         );
  NAND2_X2 U6938 ( .A1(n6596), .A2(n6595), .ZN(n3388) );
  AOI22_X2 U6939 ( .A1(n4762), .A2(regWrData[25]), .B1(memAddr[25]), .B2(n4759), .ZN(n6598) );
  AOI22_X2 U6940 ( .A1(n4778), .A2(n4677), .B1(n4757), .B2(n4341), .ZN(n6597)
         );
  NAND2_X2 U6941 ( .A1(n6598), .A2(n6597), .ZN(n3389) );
  NAND2_X2 U6942 ( .A1(n4762), .A2(regWrData[18]), .ZN(n6602) );
  NAND2_X2 U6943 ( .A1(n4759), .A2(memAddr[18]), .ZN(n6601) );
  NAND2_X2 U6944 ( .A1(n4779), .A2(n4690), .ZN(n6600) );
  NAND2_X2 U6945 ( .A1(n4757), .A2(n4708), .ZN(n6599) );
  NAND4_X2 U6946 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n3390)
         );
  NAND2_X2 U6947 ( .A1(n4762), .A2(regWrData[27]), .ZN(n6606) );
  NAND2_X2 U6948 ( .A1(memAddr[27]), .A2(n4759), .ZN(n6605) );
  NAND2_X2 U6949 ( .A1(n4779), .A2(n4691), .ZN(n6604) );
  NAND2_X2 U6950 ( .A1(n4757), .A2(n4709), .ZN(n6603) );
  NAND4_X2 U6951 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n3391)
         );
  NAND2_X2 U6952 ( .A1(n7163), .A2(regWrData[19]), .ZN(n6610) );
  NAND2_X2 U6953 ( .A1(memAddr[19]), .A2(n4758), .ZN(n6609) );
  NAND2_X2 U6954 ( .A1(n4779), .A2(n4692), .ZN(n6608) );
  NAND2_X2 U6955 ( .A1(n4757), .A2(n4710), .ZN(n6607) );
  NAND4_X2 U6956 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n3392)
         );
  OAI22_X2 U6957 ( .A1(n8663), .A2(n4789), .B1(n8851), .B2(n4777), .ZN(n3394)
         );
  NAND2_X2 U6958 ( .A1(n7163), .A2(regWrData[6]), .ZN(n6614) );
  NAND2_X2 U6959 ( .A1(n4759), .A2(memAddr[6]), .ZN(n6613) );
  NAND2_X2 U6960 ( .A1(n4779), .A2(n4693), .ZN(n6612) );
  NAND2_X2 U6961 ( .A1(n4757), .A2(n4655), .ZN(n6611) );
  NAND4_X2 U6962 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n3398)
         );
  NAND2_X2 U6963 ( .A1(n4762), .A2(regWrData[14]), .ZN(n6618) );
  NAND2_X2 U6964 ( .A1(n4759), .A2(memAddr[14]), .ZN(n6617) );
  NAND2_X2 U6965 ( .A1(n4780), .A2(n4694), .ZN(n6616) );
  NAND2_X2 U6966 ( .A1(n4757), .A2(n4671), .ZN(n6615) );
  NAND4_X2 U6967 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n3399)
         );
  INV_X4 U6968 ( .A(n6619), .ZN(n6620) );
  NAND2_X2 U6969 ( .A1(n6620), .A2(n4792), .ZN(n6621) );
  NAND2_X2 U6970 ( .A1(n4764), .A2(regWrData[23]), .ZN(n6629) );
  INV_X4 U6971 ( .A(n6622), .ZN(n6623) );
  NAND2_X2 U6972 ( .A1(n6623), .A2(n4792), .ZN(n6624) );
  INV_X4 U6973 ( .A(n6624), .ZN(n7186) );
  NAND2_X2 U6974 ( .A1(n4767), .A2(memAddr[23]), .ZN(n6628) );
  NAND2_X2 U6975 ( .A1(n4780), .A2(n4349), .ZN(n6627) );
  NAND2_X2 U6976 ( .A1(n8116), .A2(n4792), .ZN(n6625) );
  NAND2_X2 U6977 ( .A1(n4768), .A2(n4656), .ZN(n6626) );
  NAND4_X2 U6978 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n3401)
         );
  NAND2_X2 U6979 ( .A1(n4765), .A2(regWrData[24]), .ZN(n6633) );
  NAND2_X2 U6980 ( .A1(memAddr[24]), .A2(n7186), .ZN(n6632) );
  NAND2_X2 U6981 ( .A1(n4779), .A2(n4350), .ZN(n6631) );
  NAND2_X2 U6982 ( .A1(n4769), .A2(n4657), .ZN(n6630) );
  NAND4_X2 U6983 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n3403)
         );
  NAND2_X2 U6984 ( .A1(n4764), .A2(regWrData[26]), .ZN(n6637) );
  NAND2_X2 U6985 ( .A1(n4766), .A2(memAddr[26]), .ZN(n6636) );
  NAND2_X2 U6986 ( .A1(n4779), .A2(n4351), .ZN(n6635) );
  NAND2_X2 U6987 ( .A1(n4769), .A2(n4475), .ZN(n6634) );
  NAND4_X2 U6988 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n3406)
         );
  NAND2_X2 U6989 ( .A1(n7163), .A2(regWrData[3]), .ZN(n6641) );
  NAND2_X2 U6990 ( .A1(n7162), .A2(memAddr[3]), .ZN(n6640) );
  NAND2_X2 U6991 ( .A1(n4779), .A2(n4695), .ZN(n6639) );
  NAND2_X2 U6992 ( .A1(n4757), .A2(n4658), .ZN(n6638) );
  NAND4_X2 U6993 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n3409)
         );
  NAND2_X2 U6994 ( .A1(n4765), .A2(regWrData[16]), .ZN(n6645) );
  NAND2_X2 U6995 ( .A1(n4766), .A2(memAddr[16]), .ZN(n6644) );
  NAND2_X2 U6996 ( .A1(n4779), .A2(n4574), .ZN(n6643) );
  NAND2_X2 U6997 ( .A1(n4768), .A2(n4659), .ZN(n6642) );
  NAND4_X2 U6998 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n3412)
         );
  OAI22_X2 U6999 ( .A1(n8669), .A2(n4789), .B1(n8881), .B2(n4777), .ZN(n3419)
         );
  NAND2_X2 U7000 ( .A1(n4765), .A2(regWrData[13]), .ZN(n6649) );
  NAND2_X2 U7001 ( .A1(n4766), .A2(memAddr[13]), .ZN(n6648) );
  NAND2_X2 U7002 ( .A1(n4779), .A2(n4480), .ZN(n6647) );
  NAND2_X2 U7003 ( .A1(n4768), .A2(n4208), .ZN(n6646) );
  NAND4_X2 U7004 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n3423)
         );
  OAI22_X2 U7005 ( .A1(n8672), .A2(n4788), .B1(n8882), .B2(n4777), .ZN(n3425)
         );
  OAI22_X2 U7006 ( .A1(n8675), .A2(n4788), .B1(n8885), .B2(n4777), .ZN(n3430)
         );
  NAND2_X2 U7007 ( .A1(n4764), .A2(regWrData[11]), .ZN(n6653) );
  NAND2_X2 U7008 ( .A1(n4766), .A2(memAddr[11]), .ZN(n6652) );
  NAND2_X2 U7009 ( .A1(n4779), .A2(n4481), .ZN(n6651) );
  NAND2_X2 U7010 ( .A1(n4769), .A2(n4207), .ZN(n6650) );
  NAND4_X2 U7011 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n3434)
         );
  OAI22_X2 U7012 ( .A1(n8678), .A2(n4788), .B1(n8886), .B2(n4777), .ZN(n3436)
         );
  OAI22_X2 U7013 ( .A1(n8681), .A2(n4788), .B1(n8889), .B2(n4777), .ZN(n3441)
         );
  NAND2_X2 U7014 ( .A1(n4764), .A2(regWrData[9]), .ZN(n6657) );
  NAND2_X2 U7015 ( .A1(n4766), .A2(memAddr[9]), .ZN(n6656) );
  NAND2_X2 U7016 ( .A1(n4779), .A2(n4482), .ZN(n6655) );
  NAND2_X2 U7017 ( .A1(n4768), .A2(n4559), .ZN(n6654) );
  NAND4_X2 U7018 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n3445)
         );
  OAI22_X2 U7019 ( .A1(n8684), .A2(n4788), .B1(n8890), .B2(n4777), .ZN(n3447)
         );
  OAI22_X2 U7020 ( .A1(n8687), .A2(n4788), .B1(n8892), .B2(n4777), .ZN(n3452)
         );
  NAND2_X2 U7021 ( .A1(n4765), .A2(regWrData[7]), .ZN(n6661) );
  NAND2_X2 U7022 ( .A1(n4766), .A2(memAddr[7]), .ZN(n6660) );
  NAND2_X2 U7023 ( .A1(n4779), .A2(n4483), .ZN(n6659) );
  NAND2_X2 U7024 ( .A1(n4769), .A2(n4206), .ZN(n6658) );
  NAND4_X2 U7025 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n3456)
         );
  OAI22_X2 U7026 ( .A1(n8690), .A2(n4788), .B1(n8893), .B2(n4777), .ZN(n3458)
         );
  OAI22_X2 U7027 ( .A1(n8693), .A2(n4788), .B1(n8895), .B2(n4777), .ZN(n3463)
         );
  NAND2_X2 U7028 ( .A1(n4764), .A2(regWrData[5]), .ZN(n6665) );
  NAND2_X2 U7029 ( .A1(n4766), .A2(memAddr[5]), .ZN(n6664) );
  NAND2_X2 U7030 ( .A1(n4779), .A2(n4484), .ZN(n6663) );
  NAND2_X2 U7031 ( .A1(n4768), .A2(n4337), .ZN(n6662) );
  NAND4_X2 U7032 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n3467)
         );
  OAI22_X2 U7033 ( .A1(n8696), .A2(n4788), .B1(n8896), .B2(n4777), .ZN(n3469)
         );
  NAND2_X2 U7034 ( .A1(n4765), .A2(regWrData[4]), .ZN(n6669) );
  NAND2_X2 U7035 ( .A1(n4766), .A2(memAddr[4]), .ZN(n6668) );
  NAND2_X2 U7036 ( .A1(n4780), .A2(n4485), .ZN(n6667) );
  NAND2_X2 U7037 ( .A1(n4769), .A2(n4335), .ZN(n6666) );
  NAND4_X2 U7038 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n3473)
         );
  OAI22_X2 U7039 ( .A1(n8699), .A2(n4788), .B1(n8898), .B2(n4777), .ZN(n3475)
         );
  OAI22_X2 U7040 ( .A1(n8702), .A2(n4788), .B1(n8847), .B2(n4777), .ZN(n3480)
         );
  NAND2_X2 U7041 ( .A1(n4765), .A2(regWrData[3]), .ZN(n6673) );
  NAND2_X2 U7042 ( .A1(n4766), .A2(memAddr[3]), .ZN(n6672) );
  NAND2_X2 U7043 ( .A1(n4780), .A2(n4486), .ZN(n6671) );
  NAND2_X2 U7044 ( .A1(n4769), .A2(n4340), .ZN(n6670) );
  NAND4_X2 U7045 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n3484)
         );
  NAND2_X2 U7046 ( .A1(n4765), .A2(regWrData[28]), .ZN(n6677) );
  NAND2_X2 U7047 ( .A1(n4766), .A2(memAddr[28]), .ZN(n6676) );
  NAND2_X2 U7048 ( .A1(n4780), .A2(n4352), .ZN(n6675) );
  NAND2_X2 U7049 ( .A1(n4769), .A2(n4711), .ZN(n6674) );
  NAND4_X2 U7050 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n3487)
         );
  OAI22_X2 U7051 ( .A1(n8705), .A2(n4788), .B1(n8867), .B2(n4777), .ZN(n3490)
         );
  OAI22_X2 U7052 ( .A1(n8708), .A2(n4788), .B1(n8874), .B2(n4777), .ZN(n3494)
         );
  OAI22_X2 U7053 ( .A1(n8711), .A2(n4788), .B1(n8875), .B2(n4777), .ZN(n3498)
         );
  OAI22_X2 U7054 ( .A1(n8714), .A2(n4788), .B1(n8877), .B2(n4777), .ZN(n3502)
         );
  OAI22_X2 U7055 ( .A1(n8717), .A2(n4788), .B1(n8878), .B2(n4777), .ZN(n3506)
         );
  NAND2_X2 U7056 ( .A1(n4765), .A2(regWrData[14]), .ZN(n6681) );
  NAND2_X2 U7057 ( .A1(n4767), .A2(memAddr[14]), .ZN(n6680) );
  NAND2_X2 U7058 ( .A1(n4780), .A2(n4487), .ZN(n6679) );
  NAND2_X2 U7059 ( .A1(n4769), .A2(n4339), .ZN(n6678) );
  NAND4_X2 U7060 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n3510)
         );
  NAND2_X2 U7061 ( .A1(n4765), .A2(regWrData[6]), .ZN(n6685) );
  NAND2_X2 U7062 ( .A1(n4767), .A2(memAddr[6]), .ZN(n6684) );
  NAND2_X2 U7063 ( .A1(n4780), .A2(n4488), .ZN(n6683) );
  NAND2_X2 U7064 ( .A1(n4769), .A2(n4338), .ZN(n6682) );
  NAND4_X2 U7065 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n3513)
         );
  NAND2_X2 U7066 ( .A1(n4762), .A2(regWrData[5]), .ZN(n6689) );
  NAND2_X2 U7067 ( .A1(n7162), .A2(memAddr[5]), .ZN(n6688) );
  NAND2_X2 U7068 ( .A1(n4780), .A2(n4696), .ZN(n6687) );
  NAND2_X2 U7069 ( .A1(n4757), .A2(n4660), .ZN(n6686) );
  NAND4_X2 U7070 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n3516)
         );
  NAND2_X2 U7071 ( .A1(n4761), .A2(regWrData[2]), .ZN(n6693) );
  NAND2_X2 U7072 ( .A1(n4759), .A2(memAddr[2]), .ZN(n6692) );
  NAND2_X2 U7073 ( .A1(n4780), .A2(n4697), .ZN(n6691) );
  NAND2_X2 U7074 ( .A1(n4757), .A2(n4661), .ZN(n6690) );
  NAND4_X2 U7075 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n3519)
         );
  OAI22_X2 U7076 ( .A1(n8722), .A2(n4788), .B1(n8900), .B2(n4776), .ZN(n3521)
         );
  NAND2_X2 U7077 ( .A1(n4806), .A2(n6694), .ZN(n6695) );
  NAND2_X2 U7078 ( .A1(n4765), .A2(regWrData[2]), .ZN(n6699) );
  NAND2_X2 U7079 ( .A1(n4767), .A2(memAddr[2]), .ZN(n6698) );
  NAND2_X2 U7080 ( .A1(n4780), .A2(n4489), .ZN(n6697) );
  NAND2_X2 U7081 ( .A1(n4769), .A2(n4336), .ZN(n6696) );
  NAND4_X2 U7082 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n3525)
         );
  NAND2_X2 U7083 ( .A1(n4765), .A2(regWrData[30]), .ZN(n6703) );
  NAND2_X2 U7084 ( .A1(n4767), .A2(memAddr[30]), .ZN(n6702) );
  NAND2_X2 U7085 ( .A1(n4780), .A2(n4353), .ZN(n6701) );
  NAND2_X2 U7086 ( .A1(n4769), .A2(n4712), .ZN(n6700) );
  NAND4_X2 U7087 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n3528)
         );
  OAI22_X2 U7088 ( .A1(n8724), .A2(n4788), .B1(n8852), .B2(n4776), .ZN(n3530)
         );
  OAI22_X2 U7089 ( .A1(n8727), .A2(n4787), .B1(n8854), .B2(n4776), .ZN(n3534)
         );
  OAI22_X2 U7090 ( .A1(n8730), .A2(n4787), .B1(n8856), .B2(n4776), .ZN(n3538)
         );
  OAI22_X2 U7091 ( .A1(n8733), .A2(n4787), .B1(n8857), .B2(n4776), .ZN(n3542)
         );
  OAI22_X2 U7092 ( .A1(n8736), .A2(n4787), .B1(n8859), .B2(n4776), .ZN(n3546)
         );
  OAI22_X2 U7093 ( .A1(n8739), .A2(n4787), .B1(n8860), .B2(n4776), .ZN(n3550)
         );
  OAI22_X2 U7094 ( .A1(n8742), .A2(n4787), .B1(n8863), .B2(n4776), .ZN(n3554)
         );
  OAI22_X2 U7095 ( .A1(n8745), .A2(n4787), .B1(n8864), .B2(n4776), .ZN(n3558)
         );
  OAI22_X2 U7096 ( .A1(n8748), .A2(n4787), .B1(n8868), .B2(n4776), .ZN(n3562)
         );
  OAI22_X2 U7097 ( .A1(n8751), .A2(n4787), .B1(n8870), .B2(n4776), .ZN(n3566)
         );
  OAI22_X2 U7098 ( .A1(n8754), .A2(n4787), .B1(n8872), .B2(n4776), .ZN(n3570)
         );
  NAND2_X2 U7099 ( .A1(n4765), .A2(regWrData[19]), .ZN(n6707) );
  NAND2_X2 U7100 ( .A1(memAddr[19]), .A2(n7186), .ZN(n6706) );
  NAND2_X2 U7101 ( .A1(n4780), .A2(n4575), .ZN(n6705) );
  NAND2_X2 U7102 ( .A1(n4769), .A2(n4662), .ZN(n6704) );
  NAND4_X2 U7103 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n3574)
         );
  XNOR2_X2 U7104 ( .A(n6709), .B(n6708), .ZN(n6712) );
  NAND2_X2 U7105 ( .A1(n7497), .A2(n7412), .ZN(n6710) );
  NAND4_X2 U7106 ( .A1(n8424), .A2(n8423), .A3(n8425), .A4(n6713), .ZN(
        aluRes_2[19]) );
  NAND2_X2 U7107 ( .A1(memAddr[19]), .A2(n4781), .ZN(n6715) );
  NAND2_X2 U7108 ( .A1(aluRes_2[19]), .A2(n4792), .ZN(n6714) );
  NAND2_X2 U7109 ( .A1(n6715), .A2(n6714), .ZN(n9158) );
  NAND2_X2 U7110 ( .A1(n4762), .A2(regWrData[4]), .ZN(n6719) );
  NAND2_X2 U7111 ( .A1(n4758), .A2(memAddr[4]), .ZN(n6718) );
  NAND2_X2 U7112 ( .A1(n4781), .A2(n4698), .ZN(n6717) );
  NAND2_X2 U7113 ( .A1(n4757), .A2(n4713), .ZN(n6716) );
  NAND4_X2 U7114 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n3577)
         );
  NAND2_X2 U7115 ( .A1(n4765), .A2(regWrData[27]), .ZN(n6723) );
  NAND2_X2 U7116 ( .A1(memAddr[27]), .A2(n7186), .ZN(n6722) );
  NAND2_X2 U7117 ( .A1(n4781), .A2(n4354), .ZN(n6721) );
  NAND2_X2 U7118 ( .A1(n4769), .A2(n4663), .ZN(n6720) );
  NAND4_X2 U7119 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n3580)
         );
  INV_X4 U7120 ( .A(n6904), .ZN(n6747) );
  XNOR2_X2 U7121 ( .A(n6740), .B(n6739), .ZN(n6741) );
  NAND2_X2 U7122 ( .A1(n4249), .A2(n6741), .ZN(n6761) );
  XNOR2_X2 U7123 ( .A(n6760), .B(n6762), .ZN(n6742) );
  NAND2_X2 U7124 ( .A1(n4244), .A2(n6742), .ZN(n6757) );
  XNOR2_X2 U7125 ( .A(n6756), .B(n6758), .ZN(n6743) );
  NAND2_X2 U7126 ( .A1(n4223), .A2(n6743), .ZN(n6753) );
  XNOR2_X2 U7127 ( .A(n6752), .B(n6754), .ZN(n6744) );
  NAND2_X2 U7128 ( .A1(n4290), .A2(n6744), .ZN(n6749) );
  XNOR2_X2 U7129 ( .A(n6748), .B(n6750), .ZN(n6745) );
  NAND2_X2 U7130 ( .A1(n4300), .A2(n6745), .ZN(n6746) );
  INV_X4 U7131 ( .A(n6912), .ZN(n6772) );
  INV_X4 U7132 ( .A(n6748), .ZN(n6751) );
  OAI21_X4 U7133 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6773) );
  INV_X4 U7134 ( .A(n6752), .ZN(n6755) );
  OAI21_X4 U7135 ( .B1(n6755), .B2(n6754), .A(n6753), .ZN(n6777) );
  INV_X4 U7136 ( .A(n6756), .ZN(n6759) );
  INV_X4 U7137 ( .A(n6760), .ZN(n6763) );
  OAI21_X4 U7138 ( .B1(n6763), .B2(n6762), .A(n6761), .ZN(n6788) );
  XNOR2_X2 U7139 ( .A(n6765), .B(n6764), .ZN(n6766) );
  NAND2_X2 U7140 ( .A1(n4241), .A2(n6766), .ZN(n6789) );
  XNOR2_X2 U7141 ( .A(n6788), .B(n6790), .ZN(n6767) );
  NAND2_X2 U7142 ( .A1(n4250), .A2(n6767), .ZN(n6782) );
  XNOR2_X2 U7143 ( .A(n6781), .B(n6783), .ZN(n6768) );
  NAND2_X2 U7144 ( .A1(n4224), .A2(n6768), .ZN(n6778) );
  XNOR2_X2 U7145 ( .A(n6777), .B(n6779), .ZN(n6769) );
  NAND2_X2 U7146 ( .A1(n4291), .A2(n6769), .ZN(n6774) );
  XNOR2_X2 U7147 ( .A(n6773), .B(n6775), .ZN(n6770) );
  NAND2_X2 U7148 ( .A1(n4301), .A2(n6770), .ZN(n6771) );
  INV_X4 U7149 ( .A(n6773), .ZN(n6776) );
  INV_X4 U7150 ( .A(n6777), .ZN(n6780) );
  INV_X4 U7151 ( .A(n6781), .ZN(n6784) );
  OAI21_X4 U7152 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(n6807) );
  XNOR2_X2 U7153 ( .A(n6786), .B(n6785), .ZN(n6787) );
  NAND2_X2 U7154 ( .A1(n4255), .A2(n6787), .ZN(n6813) );
  INV_X4 U7155 ( .A(n6788), .ZN(n6791) );
  XNOR2_X2 U7156 ( .A(n6814), .B(n6812), .ZN(n6792) );
  NAND2_X2 U7157 ( .A1(n4242), .A2(n6792), .ZN(n6808) );
  XNOR2_X2 U7158 ( .A(n6807), .B(n6809), .ZN(n6793) );
  NAND2_X2 U7159 ( .A1(n4116), .A2(n6793), .ZN(n6803) );
  XNOR2_X2 U7160 ( .A(n6802), .B(n6804), .ZN(n6794) );
  NAND2_X2 U7161 ( .A1(n4292), .A2(n6794), .ZN(n6799) );
  XNOR2_X2 U7162 ( .A(n6798), .B(n6800), .ZN(n6796) );
  NAND2_X2 U7163 ( .A1(n7895), .A2(n4770), .ZN(n6795) );
  XNOR2_X2 U7164 ( .A(n6796), .B(n6795), .ZN(n6891) );
  INV_X4 U7165 ( .A(n6795), .ZN(n6797) );
  AOI22_X2 U7166 ( .A1(n6890), .A2(n6891), .B1(n6797), .B2(n6796), .ZN(n6923)
         );
  INV_X4 U7167 ( .A(n6798), .ZN(n6801) );
  OAI21_X4 U7168 ( .B1(n6801), .B2(n6800), .A(n6799), .ZN(n6843) );
  INV_X4 U7169 ( .A(n6802), .ZN(n6805) );
  OAI21_X4 U7170 ( .B1(n6805), .B2(n6804), .A(n6803), .ZN(n6806) );
  INV_X4 U7171 ( .A(n6806), .ZN(n6841) );
  INV_X4 U7172 ( .A(n6807), .ZN(n6810) );
  INV_X4 U7173 ( .A(n6811), .ZN(n6837) );
  INV_X4 U7174 ( .A(n6812), .ZN(n6815) );
  OAI21_X4 U7175 ( .B1(n6815), .B2(n6814), .A(n6813), .ZN(n6816) );
  INV_X4 U7176 ( .A(n6816), .ZN(n6833) );
  XNOR2_X2 U7177 ( .A(n6818), .B(n6817), .ZN(n6819) );
  NAND2_X2 U7178 ( .A1(n4256), .A2(n6819), .ZN(n6831) );
  INV_X4 U7179 ( .A(n6832), .ZN(n6820) );
  XNOR2_X2 U7180 ( .A(n6833), .B(n6820), .ZN(n6821) );
  NAND2_X2 U7181 ( .A1(n4251), .A2(n6821), .ZN(n6835) );
  INV_X4 U7182 ( .A(n6836), .ZN(n6822) );
  XNOR2_X2 U7183 ( .A(n6837), .B(n6822), .ZN(n6823) );
  NAND2_X2 U7184 ( .A1(n4117), .A2(n6823), .ZN(n6839) );
  INV_X4 U7185 ( .A(n6840), .ZN(n6824) );
  XNOR2_X2 U7186 ( .A(n6841), .B(n6824), .ZN(n6825) );
  NAND2_X2 U7187 ( .A1(n4293), .A2(n6825), .ZN(n6844) );
  XNOR2_X2 U7188 ( .A(n6843), .B(n6845), .ZN(n6826) );
  NAND2_X2 U7189 ( .A1(n4303), .A2(n6826), .ZN(n6827) );
  XNOR2_X2 U7190 ( .A(n6829), .B(n6828), .ZN(n6830) );
  NAND2_X2 U7191 ( .A1(n4263), .A2(n6830), .ZN(n6866) );
  OAI21_X4 U7192 ( .B1(n6833), .B2(n6832), .A(n6831), .ZN(n6865) );
  XNOR2_X2 U7193 ( .A(n6867), .B(n6865), .ZN(n6834) );
  NAND2_X2 U7194 ( .A1(n4257), .A2(n6834), .ZN(n6861) );
  XNOR2_X2 U7195 ( .A(n6862), .B(n6860), .ZN(n6838) );
  NAND2_X2 U7196 ( .A1(n4123), .A2(n6838), .ZN(n6856) );
  XNOR2_X2 U7197 ( .A(n6857), .B(n6855), .ZN(n6842) );
  NAND2_X2 U7198 ( .A1(n4125), .A2(n6842), .ZN(n6851) );
  INV_X4 U7199 ( .A(n6843), .ZN(n6846) );
  XNOR2_X2 U7200 ( .A(n6852), .B(n6850), .ZN(n6848) );
  NAND2_X2 U7201 ( .A1(n8349), .A2(n4770), .ZN(n6847) );
  XNOR2_X2 U7202 ( .A(n6848), .B(n6847), .ZN(n6933) );
  INV_X4 U7203 ( .A(n6847), .ZN(n6849) );
  AOI22_X2 U7204 ( .A1(n6932), .A2(n6933), .B1(n6849), .B2(n6848), .ZN(n6994)
         );
  INV_X4 U7205 ( .A(n6850), .ZN(n6853) );
  OAI21_X4 U7206 ( .B1(n6853), .B2(n6852), .A(n6851), .ZN(n6854) );
  INV_X4 U7207 ( .A(n6854), .ZN(n7012) );
  INV_X4 U7208 ( .A(n6855), .ZN(n6858) );
  OAI21_X4 U7209 ( .B1(n6858), .B2(n6857), .A(n6856), .ZN(n6859) );
  INV_X4 U7210 ( .A(n6859), .ZN(n7008) );
  INV_X4 U7211 ( .A(n6860), .ZN(n6863) );
  INV_X4 U7212 ( .A(n6864), .ZN(n7004) );
  INV_X4 U7213 ( .A(n6865), .ZN(n6868) );
  INV_X4 U7214 ( .A(n6869), .ZN(n7000) );
  XNOR2_X2 U7215 ( .A(n6871), .B(n6870), .ZN(n6872) );
  NAND2_X2 U7216 ( .A1(n4232), .A2(n6872), .ZN(n6998) );
  INV_X4 U7217 ( .A(n6999), .ZN(n6873) );
  XNOR2_X2 U7218 ( .A(n7000), .B(n6873), .ZN(n6874) );
  NAND2_X2 U7219 ( .A1(n4264), .A2(n6874), .ZN(n7002) );
  INV_X4 U7220 ( .A(n7003), .ZN(n6875) );
  XNOR2_X2 U7221 ( .A(n7004), .B(n6875), .ZN(n6876) );
  NAND2_X2 U7222 ( .A1(n4283), .A2(n6876), .ZN(n7006) );
  INV_X4 U7223 ( .A(n7007), .ZN(n6877) );
  XNOR2_X2 U7224 ( .A(n7008), .B(n6877), .ZN(n6878) );
  NAND2_X2 U7225 ( .A1(n4294), .A2(n6878), .ZN(n7010) );
  OAI21_X4 U7226 ( .B1(n4294), .B2(n6878), .A(n7010), .ZN(n7011) );
  INV_X4 U7227 ( .A(n7011), .ZN(n6879) );
  XNOR2_X2 U7228 ( .A(n7012), .B(n6879), .ZN(n6880) );
  NAND2_X2 U7229 ( .A1(n4302), .A2(n6880), .ZN(n6992) );
  XOR2_X2 U7230 ( .A(n6994), .B(n6993), .Z(n6881) );
  MUX2_X2 U7231 ( .A(n4583), .B(n6881), .S(n4078), .Z(n6889) );
  INV_X4 U7232 ( .A(n6882), .ZN(n6887) );
  NAND2_X2 U7233 ( .A1(n7243), .A2(n6883), .ZN(n6886) );
  NAND2_X2 U7234 ( .A1(n7361), .A2(n6884), .ZN(n6885) );
  OAI211_X2 U7235 ( .C1(n6887), .C2(n4169), .A(n6886), .B(n6885), .ZN(n6888)
         );
  NAND2_X2 U7236 ( .A1(n6888), .A2(n4583), .ZN(n7053) );
  XNOR2_X2 U7237 ( .A(n6891), .B(n6890), .ZN(n6896) );
  OAI221_X2 U7238 ( .B1(n6897), .B2(n7241), .C1(n6896), .C2(n4784), .A(n6895), 
        .ZN(n6898) );
  INV_X4 U7239 ( .A(n6898), .ZN(n6921) );
  NAND2_X2 U7240 ( .A1(ex_multing_set_product_in_sig_z1[24]), .A2(n4784), .ZN(
        n6920) );
  XNOR2_X2 U7241 ( .A(n6898), .B(n6920), .ZN(n7410) );
  INV_X4 U7242 ( .A(n6899), .ZN(n6902) );
  OAI21_X4 U7243 ( .B1(n6902), .B2(n6901), .A(n6900), .ZN(n7100) );
  INV_X4 U7244 ( .A(n7100), .ZN(n6910) );
  INV_X4 U7245 ( .A(n7242), .ZN(n6907) );
  XNOR2_X2 U7246 ( .A(n6904), .B(n6903), .ZN(n7272) );
  INV_X4 U7247 ( .A(n7272), .ZN(n6906) );
  NAND2_X2 U7248 ( .A1(n7244), .A2(n7243), .ZN(n6905) );
  OAI221_X2 U7249 ( .B1(n6907), .B2(n4169), .C1(n6906), .C2(n4784), .A(n6905), 
        .ZN(n6908) );
  NAND2_X2 U7250 ( .A1(n4308), .A2(n6908), .ZN(n6909) );
  INV_X4 U7251 ( .A(n7313), .ZN(n6918) );
  XNOR2_X2 U7252 ( .A(n6912), .B(n6911), .ZN(n7364) );
  INV_X4 U7253 ( .A(n7364), .ZN(n6915) );
  NAND2_X2 U7254 ( .A1(n7273), .A2(n7363), .ZN(n6914) );
  NAND2_X2 U7255 ( .A1(n7243), .A2(n7360), .ZN(n6913) );
  OAI211_X2 U7256 ( .C1(n6915), .C2(n4784), .A(n6914), .B(n6913), .ZN(n6916)
         );
  NAND3_X2 U7257 ( .A1(n6916), .A2(n4784), .A3(n4571), .ZN(n6917) );
  NAND2_X2 U7258 ( .A1(n7410), .A2(n7409), .ZN(n6919) );
  OAI21_X4 U7259 ( .B1(n6921), .B2(n6920), .A(n6919), .ZN(n6969) );
  INV_X4 U7260 ( .A(n6969), .ZN(n6931) );
  XNOR2_X2 U7261 ( .A(n6923), .B(n6922), .ZN(n6928) );
  AOI22_X2 U7262 ( .A1(n7361), .A2(n4205), .B1(n7243), .B2(n6924), .ZN(n6927)
         );
  NAND2_X2 U7263 ( .A1(n7273), .A2(n6925), .ZN(n6926) );
  OAI211_X2 U7264 ( .C1(n4784), .C2(n6928), .A(n6927), .B(n6926), .ZN(n6929)
         );
  NAND3_X2 U7265 ( .A1(n6929), .A2(n4784), .A3(n4572), .ZN(n6930) );
  INV_X4 U7266 ( .A(n7303), .ZN(n6941) );
  XNOR2_X2 U7267 ( .A(n6933), .B(n6932), .ZN(n6938) );
  OAI221_X2 U7268 ( .B1(n4389), .B2(n4169), .C1(n6938), .C2(n4784), .A(n6937), 
        .ZN(n6939) );
  NAND2_X2 U7269 ( .A1(n4309), .A2(n6939), .ZN(n6940) );
  OAI21_X4 U7270 ( .B1(n6941), .B2(n7302), .A(n6940), .ZN(n7052) );
  XNOR2_X2 U7271 ( .A(n7054), .B(n7052), .ZN(n6945) );
  NAND2_X2 U7272 ( .A1(n6942), .A2(n7412), .ZN(n6943) );
  NAND4_X2 U7273 ( .A1(n8345), .A2(n8344), .A3(n8346), .A4(n6946), .ZN(
        aluRes_2[27]) );
  NAND2_X2 U7274 ( .A1(n4781), .A2(memAddr[27]), .ZN(n6948) );
  NAND2_X2 U7275 ( .A1(aluRes_2[27]), .A2(n4792), .ZN(n6947) );
  NAND2_X2 U7276 ( .A1(n6948), .A2(n6947), .ZN(n9166) );
  NAND2_X2 U7277 ( .A1(n4765), .A2(regWrData[18]), .ZN(n6952) );
  NAND2_X2 U7278 ( .A1(n4767), .A2(memAddr[18]), .ZN(n6951) );
  NAND2_X2 U7279 ( .A1(n4781), .A2(n4576), .ZN(n6950) );
  NAND2_X2 U7280 ( .A1(n4769), .A2(n4568), .ZN(n6949) );
  NAND4_X2 U7281 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n3583)
         );
  INV_X4 U7282 ( .A(n8436), .ZN(n6953) );
  XNOR2_X2 U7283 ( .A(n6955), .B(n6954), .ZN(n6958) );
  NAND2_X2 U7284 ( .A1(n7495), .A2(n7412), .ZN(n6956) );
  NAND3_X2 U7285 ( .A1(n8437), .A2(n6960), .A3(n6959), .ZN(aluRes_2[18]) );
  NAND2_X2 U7286 ( .A1(n4781), .A2(memAddr[18]), .ZN(n6962) );
  NAND2_X2 U7287 ( .A1(aluRes_2[18]), .A2(n4792), .ZN(n6961) );
  NAND2_X2 U7288 ( .A1(n6962), .A2(n6961), .ZN(n9157) );
  NAND2_X2 U7289 ( .A1(n4765), .A2(regWrData[25]), .ZN(n6966) );
  NAND2_X2 U7290 ( .A1(memAddr[25]), .A2(n7186), .ZN(n6965) );
  NAND2_X2 U7291 ( .A1(n4780), .A2(n4355), .ZN(n6964) );
  NAND2_X2 U7292 ( .A1(n4769), .A2(n4664), .ZN(n6963) );
  NAND4_X2 U7293 ( .A1(n6966), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n3586)
         );
  INV_X4 U7294 ( .A(n8357), .ZN(n6967) );
  XNOR2_X2 U7295 ( .A(n6969), .B(n6968), .ZN(n6972) );
  NAND2_X2 U7296 ( .A1(n7501), .A2(n7412), .ZN(n6970) );
  NAND3_X2 U7297 ( .A1(n8358), .A2(n6974), .A3(n6973), .ZN(aluRes_2[25]) );
  NAND2_X2 U7298 ( .A1(n4780), .A2(memAddr[25]), .ZN(n6976) );
  NAND2_X2 U7299 ( .A1(aluRes_2[25]), .A2(n4792), .ZN(n6975) );
  NAND2_X2 U7300 ( .A1(n6976), .A2(n6975), .ZN(n9164) );
  NAND2_X2 U7301 ( .A1(n4765), .A2(regWrData[8]), .ZN(n6980) );
  NAND2_X2 U7302 ( .A1(n4767), .A2(memAddr[8]), .ZN(n6979) );
  NAND2_X2 U7303 ( .A1(n4780), .A2(n4490), .ZN(n6978) );
  NAND2_X2 U7304 ( .A1(n4769), .A2(n4560), .ZN(n6977) );
  NAND4_X2 U7305 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n3589)
         );
  AOI22_X2 U7306 ( .A1(n4132), .A2(n4560), .B1(n4096), .B2(regWrData[8]), .ZN(
        n6986) );
  INV_X4 U7307 ( .A(n7914), .ZN(n6981) );
  NAND2_X2 U7308 ( .A1(n6981), .A2(n7565), .ZN(n6985) );
  NAND2_X2 U7309 ( .A1(n7677), .A2(memAddr[8]), .ZN(n6984) );
  AOI22_X2 U7310 ( .A1(n7506), .A2(n7508), .B1(n7507), .B2(n6982), .ZN(n6983)
         );
  NAND4_X2 U7311 ( .A1(n6986), .A2(n6985), .A3(n6984), .A4(n6983), .ZN(n3591)
         );
  NAND2_X2 U7312 ( .A1(n4764), .A2(regWrData[29]), .ZN(n6990) );
  NAND2_X2 U7313 ( .A1(n4767), .A2(memAddr[29]), .ZN(n6989) );
  NAND2_X2 U7314 ( .A1(n4780), .A2(n4356), .ZN(n6988) );
  NAND2_X2 U7315 ( .A1(n4768), .A2(n4714), .ZN(n6987) );
  NAND4_X2 U7316 ( .A1(n6990), .A2(n6989), .A3(n6988), .A4(n6987), .ZN(n3592)
         );
  NAND2_X2 U7317 ( .A1(n6991), .A2(n8335), .ZN(n7069) );
  XNOR2_X2 U7318 ( .A(n6996), .B(n6995), .ZN(n6997) );
  NAND2_X2 U7319 ( .A1(n4266), .A2(n6997), .ZN(n7031) );
  XNOR2_X2 U7320 ( .A(n7032), .B(n7030), .ZN(n7001) );
  NAND2_X2 U7321 ( .A1(n4297), .A2(n7001), .ZN(n7026) );
  OAI21_X4 U7322 ( .B1(n7004), .B2(n7003), .A(n7002), .ZN(n7025) );
  XNOR2_X2 U7323 ( .A(n7027), .B(n7025), .ZN(n7005) );
  NAND2_X2 U7324 ( .A1(n4284), .A2(n7005), .ZN(n7022) );
  OAI21_X4 U7325 ( .B1(n7008), .B2(n7007), .A(n7006), .ZN(n7021) );
  XNOR2_X2 U7326 ( .A(n7023), .B(n7021), .ZN(n7009) );
  NAND2_X2 U7327 ( .A1(n4285), .A2(n7009), .ZN(n7017) );
  OAI21_X4 U7328 ( .B1(n7012), .B2(n7011), .A(n7010), .ZN(n7016) );
  XNOR2_X2 U7329 ( .A(n7018), .B(n7016), .ZN(n7014) );
  NAND2_X2 U7330 ( .A1(n8336), .A2(n7266), .ZN(n7013) );
  XNOR2_X2 U7331 ( .A(n7014), .B(n7013), .ZN(n7057) );
  INV_X4 U7332 ( .A(n7013), .ZN(n7015) );
  AOI22_X2 U7333 ( .A1(n7056), .A2(n7057), .B1(n7015), .B2(n7014), .ZN(n7270)
         );
  INV_X4 U7334 ( .A(n7016), .ZN(n7019) );
  INV_X4 U7335 ( .A(n7020), .ZN(n7265) );
  INV_X4 U7336 ( .A(n7021), .ZN(n7024) );
  INV_X4 U7337 ( .A(n7025), .ZN(n7028) );
  INV_X4 U7338 ( .A(n7029), .ZN(n7254) );
  INV_X4 U7339 ( .A(n7030), .ZN(n7033) );
  OAI21_X4 U7340 ( .B1(n7033), .B2(n7032), .A(n7031), .ZN(n7248) );
  XNOR2_X2 U7341 ( .A(n7035), .B(n7034), .ZN(n7036) );
  NAND2_X2 U7342 ( .A1(n4248), .A2(n7036), .ZN(n7249) );
  XNOR2_X2 U7343 ( .A(n7248), .B(n7250), .ZN(n7037) );
  NAND2_X2 U7344 ( .A1(n4311), .A2(n7037), .ZN(n7252) );
  INV_X4 U7345 ( .A(n7253), .ZN(n7038) );
  XNOR2_X2 U7346 ( .A(n7254), .B(n7038), .ZN(n7039) );
  NAND2_X2 U7347 ( .A1(n4288), .A2(n7039), .ZN(n7260) );
  XNOR2_X2 U7348 ( .A(n7259), .B(n7261), .ZN(n7040) );
  NAND2_X2 U7349 ( .A1(n4286), .A2(n7040), .ZN(n7263) );
  INV_X4 U7350 ( .A(n7264), .ZN(n7041) );
  XNOR2_X2 U7351 ( .A(n7265), .B(n7041), .ZN(n7042) );
  NAND2_X2 U7352 ( .A1(n4304), .A2(n7042), .ZN(n7268) );
  XOR2_X2 U7353 ( .A(n7270), .B(n7269), .Z(n7043) );
  MUX2_X2 U7354 ( .A(n4584), .B(n7043), .S(n4078), .Z(n7051) );
  INV_X4 U7355 ( .A(n7044), .ZN(n7049) );
  NAND2_X2 U7356 ( .A1(n7243), .A2(n7045), .ZN(n7048) );
  NAND2_X2 U7357 ( .A1(n7361), .A2(n7046), .ZN(n7047) );
  OAI211_X2 U7358 ( .C1(n7049), .C2(n4169), .A(n7048), .B(n7047), .ZN(n7050)
         );
  NAND2_X2 U7359 ( .A1(n7050), .A2(n4584), .ZN(n7236) );
  INV_X4 U7360 ( .A(n7052), .ZN(n7055) );
  INV_X4 U7361 ( .A(n7287), .ZN(n7066) );
  XNOR2_X2 U7362 ( .A(n7057), .B(n7056), .ZN(n7063) );
  AOI22_X2 U7363 ( .A1(n6568), .A2(n7361), .B1(n7243), .B2(n7059), .ZN(n7062)
         );
  NAND2_X2 U7364 ( .A1(n7273), .A2(n7060), .ZN(n7061) );
  OAI211_X2 U7365 ( .C1(n4784), .C2(n7063), .A(n7062), .B(n7061), .ZN(n7064)
         );
  NAND2_X2 U7366 ( .A1(n4310), .A2(n7064), .ZN(n7065) );
  XNOR2_X2 U7367 ( .A(n7237), .B(n7235), .ZN(n7067) );
  AOI21_X2 U7368 ( .B1(n7067), .B2(n4794), .A(n4509), .ZN(n7068) );
  NAND4_X2 U7369 ( .A1(n8330), .A2(n8329), .A3(n7069), .A4(n7068), .ZN(
        aluRes_2[29]) );
  NAND2_X2 U7370 ( .A1(aluRes_2[29]), .A2(n4792), .ZN(n7070) );
  NAND2_X2 U7371 ( .A1(n4764), .A2(regWrData[12]), .ZN(n7074) );
  NAND2_X2 U7372 ( .A1(n4767), .A2(memAddr[12]), .ZN(n7073) );
  NAND2_X2 U7373 ( .A1(n4780), .A2(n4491), .ZN(n7072) );
  NAND2_X2 U7374 ( .A1(n4768), .A2(n4334), .ZN(n7071) );
  NAND4_X2 U7375 ( .A1(n7074), .A2(n7073), .A3(n7072), .A4(n7071), .ZN(n3595)
         );
  NAND2_X2 U7376 ( .A1(n4764), .A2(regWrData[17]), .ZN(n7078) );
  NAND2_X2 U7377 ( .A1(memAddr[17]), .A2(n7186), .ZN(n7077) );
  NAND2_X2 U7378 ( .A1(n4780), .A2(n4577), .ZN(n7076) );
  NAND2_X2 U7379 ( .A1(n4768), .A2(n4665), .ZN(n7075) );
  NAND4_X2 U7380 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n3598)
         );
  XNOR2_X2 U7381 ( .A(n7080), .B(n7079), .ZN(n7083) );
  NAND2_X2 U7382 ( .A1(n7496), .A2(n7412), .ZN(n7081) );
  NAND4_X2 U7383 ( .A1(n7892), .A2(n7891), .A3(n7893), .A4(n7084), .ZN(n9183)
         );
  NAND2_X2 U7384 ( .A1(n4780), .A2(memAddr[17]), .ZN(n7086) );
  NAND2_X2 U7385 ( .A1(n9183), .A2(n4791), .ZN(n7085) );
  NAND2_X2 U7386 ( .A1(n7086), .A2(n7085), .ZN(n3600) );
  AOI22_X2 U7387 ( .A1(n4761), .A2(regWrData[9]), .B1(n4758), .B2(memAddr[9]), 
        .ZN(n7088) );
  AOI22_X2 U7388 ( .A1(n4779), .A2(n4678), .B1(n4757), .B2(n4345), .ZN(n7087)
         );
  NAND2_X2 U7389 ( .A1(n7088), .A2(n7087), .ZN(n3601) );
  NAND2_X2 U7390 ( .A1(n7652), .A2(n7565), .ZN(n7093) );
  AOI22_X2 U7391 ( .A1(n4132), .A2(n4559), .B1(n4096), .B2(regWrData[9]), .ZN(
        n7092) );
  NAND2_X2 U7392 ( .A1(n7677), .A2(memAddr[9]), .ZN(n7091) );
  AOI22_X2 U7393 ( .A1(n7651), .A2(n7506), .B1(n7507), .B2(n7089), .ZN(n7090)
         );
  NAND4_X2 U7394 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n3603)
         );
  NAND2_X2 U7395 ( .A1(n4764), .A2(regWrData[22]), .ZN(n7097) );
  NAND2_X2 U7396 ( .A1(memAddr[22]), .A2(n7186), .ZN(n7096) );
  NAND2_X2 U7397 ( .A1(n4781), .A2(n4357), .ZN(n7095) );
  NAND2_X2 U7398 ( .A1(n4768), .A2(n4666), .ZN(n7094) );
  NAND4_X2 U7399 ( .A1(n7097), .A2(n7096), .A3(n7095), .A4(n7094), .ZN(n3604)
         );
  INV_X4 U7400 ( .A(n8385), .ZN(n7098) );
  XNOR2_X2 U7401 ( .A(n7100), .B(n7099), .ZN(n7103) );
  NAND2_X2 U7402 ( .A1(n7529), .A2(n7412), .ZN(n7101) );
  NAND3_X2 U7403 ( .A1(n8386), .A2(n7105), .A3(n7104), .ZN(aluRes_2[22]) );
  NAND2_X2 U7404 ( .A1(memAddr[22]), .A2(n4782), .ZN(n7107) );
  NAND2_X2 U7405 ( .A1(aluRes_2[22]), .A2(n4791), .ZN(n7106) );
  NAND2_X2 U7406 ( .A1(n7107), .A2(n7106), .ZN(n9161) );
  NAND2_X2 U7407 ( .A1(n4764), .A2(regWrData[21]), .ZN(n7111) );
  NAND2_X2 U7408 ( .A1(memAddr[21]), .A2(n7186), .ZN(n7110) );
  NAND2_X2 U7409 ( .A1(n4781), .A2(n4358), .ZN(n7109) );
  NAND2_X2 U7410 ( .A1(n4768), .A2(n4667), .ZN(n7108) );
  NAND4_X2 U7411 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n3607)
         );
  OAI22_X2 U7412 ( .A1(n8759), .A2(n4787), .B1(n4368), .B2(n4776), .ZN(n3609)
         );
  INV_X4 U7413 ( .A(n7112), .ZN(n7113) );
  NAND2_X2 U7414 ( .A1(iAddr[1]), .A2(n4806), .ZN(n7114) );
  NAND2_X2 U7415 ( .A1(n4764), .A2(regWrData[1]), .ZN(n7118) );
  NAND2_X2 U7416 ( .A1(n4767), .A2(memAddr[1]), .ZN(n7117) );
  NAND2_X2 U7417 ( .A1(n4781), .A2(n4672), .ZN(n7116) );
  NAND2_X2 U7418 ( .A1(n4768), .A2(n4371), .ZN(n7115) );
  NAND4_X2 U7419 ( .A1(n7118), .A2(n7117), .A3(n7116), .A4(n7115), .ZN(n3613)
         );
  AOI22_X2 U7420 ( .A1(n4761), .A2(regWrData[0]), .B1(n4758), .B2(memAddr[0]), 
        .ZN(n7120) );
  AOI22_X2 U7421 ( .A1(n4778), .A2(n4679), .B1(n4757), .B2(n4348), .ZN(n7119)
         );
  NAND2_X2 U7422 ( .A1(n7120), .A2(n7119), .ZN(n3615) );
  OAI22_X2 U7423 ( .A1(n4361), .A2(n4787), .B1(n4612), .B2(n4776), .ZN(n3619)
         );
  OAI22_X2 U7424 ( .A1(n8927), .A2(n4787), .B1(n8763), .B2(n4776), .ZN(n3621)
         );
  OAI22_X2 U7425 ( .A1(n8910), .A2(n4787), .B1(n8764), .B2(n4776), .ZN(n3623)
         );
  OAI22_X2 U7426 ( .A1(n8766), .A2(n4787), .B1(n8765), .B2(n4776), .ZN(n3625)
         );
  OAI22_X2 U7427 ( .A1(n8768), .A2(n4787), .B1(n8767), .B2(n4776), .ZN(n3627)
         );
  OAI22_X2 U7428 ( .A1(n8770), .A2(n4787), .B1(n8769), .B2(n4775), .ZN(n3629)
         );
  OAI22_X2 U7429 ( .A1(n8772), .A2(n4787), .B1(n8771), .B2(n4775), .ZN(n3631)
         );
  OAI22_X2 U7430 ( .A1(n8914), .A2(n4788), .B1(n8773), .B2(n4775), .ZN(n3633)
         );
  OAI22_X2 U7431 ( .A1(n8913), .A2(n4788), .B1(n8774), .B2(n4775), .ZN(n3635)
         );
  OAI22_X2 U7432 ( .A1(n8912), .A2(n4788), .B1(n8775), .B2(n4775), .ZN(n3637)
         );
  OAI22_X2 U7433 ( .A1(n8911), .A2(n4788), .B1(n8776), .B2(n4775), .ZN(n3639)
         );
  OAI22_X2 U7434 ( .A1(n8909), .A2(n4788), .B1(n8777), .B2(n4775), .ZN(n3641)
         );
  OAI22_X2 U7435 ( .A1(n8925), .A2(n4788), .B1(n8778), .B2(n4775), .ZN(n3643)
         );
  OAI22_X2 U7436 ( .A1(n8923), .A2(n4788), .B1(n8779), .B2(n4775), .ZN(n3645)
         );
  OAI22_X2 U7437 ( .A1(n8924), .A2(n4788), .B1(n8780), .B2(n4775), .ZN(n3647)
         );
  OAI22_X2 U7438 ( .A1(n8922), .A2(n4788), .B1(n8781), .B2(n4775), .ZN(n3649)
         );
  OAI22_X2 U7439 ( .A1(n8921), .A2(n4788), .B1(n8782), .B2(n4775), .ZN(n3651)
         );
  OAI22_X2 U7440 ( .A1(n8920), .A2(n4788), .B1(n8783), .B2(n4775), .ZN(n3653)
         );
  OAI22_X2 U7441 ( .A1(n8919), .A2(n4788), .B1(n8784), .B2(n4775), .ZN(n3655)
         );
  OAI22_X2 U7442 ( .A1(n8786), .A2(n4788), .B1(n8785), .B2(n4775), .ZN(n3657)
         );
  OAI22_X2 U7443 ( .A1(n8931), .A2(n4788), .B1(n8787), .B2(n4775), .ZN(n3659)
         );
  OAI22_X2 U7444 ( .A1(n8788), .A2(n4788), .B1(n4532), .B2(n4775), .ZN(n3663)
         );
  INV_X4 U7445 ( .A(n7121), .ZN(n7122) );
  NAND2_X2 U7446 ( .A1(n4806), .A2(iAddr[0]), .ZN(n7124) );
  INV_X4 U7447 ( .A(n7125), .ZN(n7127) );
  OAI22_X2 U7448 ( .A1(n4610), .A2(n4788), .B1(n4360), .B2(n4775), .ZN(n3670)
         );
  OAI22_X2 U7449 ( .A1(n8791), .A2(n4788), .B1(n8790), .B2(n4774), .ZN(n3672)
         );
  OAI22_X2 U7450 ( .A1(n8917), .A2(n4786), .B1(n8792), .B2(n4774), .ZN(n3674)
         );
  OAI22_X2 U7451 ( .A1(n8918), .A2(n4786), .B1(n8793), .B2(n4774), .ZN(n3676)
         );
  OAI22_X2 U7452 ( .A1(n8928), .A2(n4786), .B1(n8794), .B2(n4774), .ZN(n3678)
         );
  OAI22_X2 U7453 ( .A1(n8930), .A2(n4786), .B1(n8795), .B2(n4774), .ZN(n3680)
         );
  OAI22_X2 U7454 ( .A1(n8929), .A2(n4786), .B1(n8796), .B2(n4774), .ZN(n3682)
         );
  OAI22_X2 U7455 ( .A1(n8926), .A2(n4786), .B1(n8797), .B2(n4774), .ZN(n3684)
         );
  OAI22_X2 U7456 ( .A1(n8915), .A2(n4786), .B1(n8798), .B2(n4774), .ZN(n3688)
         );
  OAI22_X2 U7457 ( .A1(n8800), .A2(n4786), .B1(n8799), .B2(n4774), .ZN(n3692)
         );
  AOI22_X2 U7458 ( .A1(n4761), .A2(regWrData[1]), .B1(n4758), .B2(memAddr[1]), 
        .ZN(n7129) );
  AOI22_X2 U7459 ( .A1(n4778), .A2(n4680), .B1(n4757), .B2(n4347), .ZN(n7128)
         );
  NAND2_X2 U7460 ( .A1(n7129), .A2(n7128), .ZN(n3696) );
  NAND2_X2 U7461 ( .A1(n4761), .A2(regWrData[7]), .ZN(n7133) );
  NAND2_X2 U7462 ( .A1(n7162), .A2(memAddr[7]), .ZN(n7132) );
  NAND2_X2 U7463 ( .A1(n4780), .A2(n4699), .ZN(n7131) );
  NAND2_X2 U7464 ( .A1(n4757), .A2(n4668), .ZN(n7130) );
  NAND4_X2 U7465 ( .A1(n7133), .A2(n7132), .A3(n7131), .A4(n7130), .ZN(n3697)
         );
  NAND2_X2 U7466 ( .A1(n4761), .A2(regWrData[11]), .ZN(n7137) );
  NAND2_X2 U7467 ( .A1(n4759), .A2(memAddr[11]), .ZN(n7136) );
  NAND2_X2 U7468 ( .A1(n4781), .A2(n4700), .ZN(n7135) );
  NAND2_X2 U7469 ( .A1(n4757), .A2(n4715), .ZN(n7134) );
  NAND4_X2 U7470 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(n3698)
         );
  NAND2_X2 U7471 ( .A1(n4762), .A2(regWrData[13]), .ZN(n7141) );
  NAND2_X2 U7472 ( .A1(n4759), .A2(memAddr[13]), .ZN(n7140) );
  NAND2_X2 U7473 ( .A1(n4781), .A2(n4701), .ZN(n7139) );
  NAND2_X2 U7474 ( .A1(n4757), .A2(n4669), .ZN(n7138) );
  NAND4_X2 U7475 ( .A1(n7141), .A2(n7140), .A3(n7139), .A4(n7138), .ZN(n3699)
         );
  AOI22_X2 U7476 ( .A1(n4761), .A2(regWrData[16]), .B1(n4758), .B2(memAddr[16]), .ZN(n7143) );
  AOI22_X2 U7477 ( .A1(n4778), .A2(n4681), .B1(n4757), .B2(n4344), .ZN(n7142)
         );
  NAND2_X2 U7478 ( .A1(n7143), .A2(n7142), .ZN(n3700) );
  AOI22_X2 U7479 ( .A1(n4761), .A2(regWrData[23]), .B1(n4758), .B2(memAddr[23]), .ZN(n7147) );
  NAND2_X2 U7480 ( .A1(n7147), .A2(n7146), .ZN(n3701) );
  AOI22_X2 U7481 ( .A1(n4761), .A2(regWrData[24]), .B1(memAddr[24]), .B2(n4758), .ZN(n7149) );
  AOI22_X2 U7482 ( .A1(n4778), .A2(n4682), .B1(n4757), .B2(n4342), .ZN(n7148)
         );
  NAND2_X2 U7483 ( .A1(n7149), .A2(n7148), .ZN(n3702) );
  AOI22_X2 U7484 ( .A1(n4761), .A2(regWrData[26]), .B1(n4758), .B2(memAddr[26]), .ZN(n7153) );
  NAND2_X2 U7485 ( .A1(n7153), .A2(n7152), .ZN(n3703) );
  AOI22_X2 U7486 ( .A1(n4761), .A2(regWrData[28]), .B1(n4758), .B2(memAddr[28]), .ZN(n7157) );
  NAND2_X2 U7487 ( .A1(n7157), .A2(n7156), .ZN(n3704) );
  AOI22_X2 U7488 ( .A1(n4761), .A2(regWrData[30]), .B1(n4758), .B2(memAddr[30]), .ZN(n7161) );
  NAND2_X2 U7489 ( .A1(n7161), .A2(n7160), .ZN(n3705) );
  AOI22_X2 U7490 ( .A1(n4761), .A2(regWrData[31]), .B1(n4758), .B2(memAddr[31]), .ZN(n7168) );
  NAND2_X2 U7491 ( .A1(n7168), .A2(n7167), .ZN(n3706) );
  OAI22_X2 U7492 ( .A1(n8839), .A2(n4786), .B1(n8901), .B2(n4774), .ZN(n3707)
         );
  OAI22_X2 U7493 ( .A1(n8818), .A2(n4786), .B1(n8812), .B2(n4774), .ZN(n3708)
         );
  OAI22_X2 U7494 ( .A1(n8840), .A2(n4786), .B1(n8899), .B2(n4774), .ZN(n3709)
         );
  OAI22_X2 U7495 ( .A1(n8819), .A2(n4786), .B1(n8813), .B2(n4774), .ZN(n3710)
         );
  OAI22_X2 U7496 ( .A1(n8964), .A2(n4786), .B1(n8965), .B2(n4774), .ZN(n9174)
         );
  OAI22_X2 U7497 ( .A1(n8820), .A2(n4786), .B1(n8897), .B2(n4774), .ZN(n3712)
         );
  OAI22_X2 U7498 ( .A1(n8962), .A2(n4786), .B1(n8963), .B2(n4774), .ZN(n9175)
         );
  OAI22_X2 U7499 ( .A1(n8821), .A2(n4786), .B1(n8894), .B2(n4773), .ZN(n3714)
         );
  OAI22_X2 U7500 ( .A1(n8960), .A2(n4786), .B1(n8961), .B2(n4774), .ZN(n9176)
         );
  OAI22_X2 U7501 ( .A1(n8822), .A2(n4786), .B1(n8891), .B2(n4773), .ZN(n3716)
         );
  OAI22_X2 U7502 ( .A1(n8823), .A2(n4785), .B1(n8888), .B2(n4773), .ZN(n3717)
         );
  OAI22_X2 U7503 ( .A1(n8825), .A2(n4785), .B1(n8887), .B2(n4773), .ZN(n3718)
         );
  OAI22_X2 U7504 ( .A1(n8828), .A2(n4785), .B1(n8884), .B2(n4773), .ZN(n3719)
         );
  OAI22_X2 U7505 ( .A1(n8830), .A2(n4785), .B1(n8883), .B2(n4773), .ZN(n3720)
         );
  OAI22_X2 U7506 ( .A1(n8833), .A2(n4788), .B1(n8880), .B2(n4773), .ZN(n3721)
         );
  OAI22_X2 U7507 ( .A1(n8837), .A2(n4785), .B1(n8879), .B2(n4773), .ZN(n3722)
         );
  OAI22_X2 U7508 ( .A1(n8974), .A2(n4785), .B1(n8975), .B2(n4773), .ZN(n9169)
         );
  OAI22_X2 U7509 ( .A1(n8943), .A2(n4785), .B1(n8876), .B2(n4773), .ZN(n3724)
         );
  OAI22_X2 U7510 ( .A1(n8972), .A2(n4785), .B1(n8973), .B2(n4773), .ZN(n9170)
         );
  OAI22_X2 U7511 ( .A1(n8942), .A2(n4785), .B1(n8873), .B2(n4773), .ZN(n3726)
         );
  OAI22_X2 U7512 ( .A1(n8970), .A2(n4785), .B1(n8971), .B2(n4773), .ZN(n9171)
         );
  OAI22_X2 U7513 ( .A1(n8941), .A2(n4785), .B1(n8869), .B2(n4773), .ZN(n3728)
         );
  OAI22_X2 U7514 ( .A1(n8939), .A2(n4785), .B1(n8866), .B2(n4773), .ZN(n3729)
         );
  OAI22_X2 U7515 ( .A1(n8937), .A2(n4785), .B1(n8865), .B2(n4773), .ZN(n3730)
         );
  OAI22_X2 U7516 ( .A1(n8935), .A2(n4785), .B1(n8862), .B2(n4772), .ZN(n3731)
         );
  OAI22_X2 U7517 ( .A1(n8933), .A2(n4785), .B1(n8861), .B2(n4772), .ZN(n3732)
         );
  OAI22_X2 U7518 ( .A1(n8968), .A2(n4785), .B1(n8969), .B2(n4772), .ZN(n9172)
         );
  OAI22_X2 U7519 ( .A1(n8826), .A2(n4785), .B1(n8858), .B2(n4773), .ZN(n3734)
         );
  OAI22_X2 U7520 ( .A1(n8966), .A2(n4785), .B1(n8967), .B2(n4772), .ZN(n9173)
         );
  OAI22_X2 U7521 ( .A1(n8831), .A2(n4788), .B1(n8855), .B2(n4772), .ZN(n3736)
         );
  OAI22_X2 U7522 ( .A1(n8834), .A2(n4788), .B1(n8853), .B2(n4772), .ZN(n3737)
         );
  OAI22_X2 U7523 ( .A1(n8836), .A2(n4787), .B1(n8850), .B2(n4772), .ZN(n3738)
         );
  OAI22_X2 U7524 ( .A1(n8845), .A2(n4788), .B1(n8814), .B2(n4773), .ZN(n3740)
         );
  OAI22_X2 U7525 ( .A1(n8844), .A2(n4788), .B1(n8986), .B2(n4772), .ZN(n3742)
         );
  OAI22_X2 U7526 ( .A1(n8843), .A2(n4787), .B1(n8903), .B2(n4772), .ZN(n3743)
         );
  OAI22_X2 U7527 ( .A1(n8932), .A2(n4788), .B1(n8815), .B2(n4772), .ZN(n3745)
         );
  NAND2_X2 U7528 ( .A1(op0_2), .A2(n4791), .ZN(n7169) );
  OAI22_X2 U7529 ( .A1(n4324), .A2(n4788), .B1(n4092), .B2(n4772), .ZN(n3748)
         );
  OAI22_X2 U7530 ( .A1(n4533), .A2(n4788), .B1(n4320), .B2(n4772), .ZN(n3750)
         );
  NAND2_X2 U7531 ( .A1(n4764), .A2(regWrData[0]), .ZN(n7173) );
  NAND2_X2 U7532 ( .A1(n4766), .A2(memAddr[0]), .ZN(n7172) );
  NAND2_X2 U7533 ( .A1(n4781), .A2(n4673), .ZN(n7171) );
  NAND2_X2 U7534 ( .A1(n4768), .A2(n4372), .ZN(n7170) );
  NAND4_X2 U7535 ( .A1(n7173), .A2(n7172), .A3(n7171), .A4(n7170), .ZN(n3751)
         );
  NAND2_X2 U7536 ( .A1(n4764), .A2(regWrData[10]), .ZN(n7177) );
  NAND2_X2 U7537 ( .A1(n4767), .A2(memAddr[10]), .ZN(n7176) );
  NAND2_X2 U7538 ( .A1(n4781), .A2(n4492), .ZN(n7175) );
  NAND2_X2 U7539 ( .A1(n4768), .A2(n4209), .ZN(n7174) );
  NAND4_X2 U7540 ( .A1(n7177), .A2(n7176), .A3(n7175), .A4(n7174), .ZN(n3752)
         );
  NAND2_X2 U7541 ( .A1(n4764), .A2(regWrData[15]), .ZN(n7181) );
  NAND2_X2 U7542 ( .A1(n7186), .A2(memAddr[15]), .ZN(n7180) );
  NAND2_X2 U7543 ( .A1(n4779), .A2(n4578), .ZN(n7179) );
  NAND2_X2 U7544 ( .A1(n4768), .A2(n4418), .ZN(n7178) );
  NAND4_X2 U7545 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n3753)
         );
  NAND2_X2 U7546 ( .A1(n4764), .A2(regWrData[20]), .ZN(n7185) );
  NAND2_X2 U7547 ( .A1(n4767), .A2(memAddr[20]), .ZN(n7184) );
  NAND2_X2 U7548 ( .A1(n4781), .A2(n4579), .ZN(n7183) );
  NAND2_X2 U7549 ( .A1(n4768), .A2(n4417), .ZN(n7182) );
  NAND4_X2 U7550 ( .A1(n7185), .A2(n7184), .A3(n7183), .A4(n7182), .ZN(n3754)
         );
  NAND2_X2 U7551 ( .A1(n4764), .A2(regWrData[31]), .ZN(n7190) );
  NAND2_X2 U7552 ( .A1(n4766), .A2(memAddr[31]), .ZN(n7189) );
  NAND2_X2 U7553 ( .A1(n4781), .A2(n4359), .ZN(n7188) );
  NAND2_X2 U7554 ( .A1(n4768), .A2(n4474), .ZN(n7187) );
  NAND4_X2 U7555 ( .A1(n7190), .A2(n7189), .A3(n7188), .A4(n7187), .ZN(n3755)
         );
  OAI22_X2 U7556 ( .A1(n4095), .A2(n4788), .B1(n4081), .B2(n4772), .ZN(n3757)
         );
  OAI22_X2 U7557 ( .A1(n4322), .A2(n4787), .B1(n4093), .B2(n4772), .ZN(n3759)
         );
  OAI22_X2 U7558 ( .A1(n4094), .A2(n4787), .B1(n4319), .B2(n4772), .ZN(n3761)
         );
  NAND4_X2 U7559 ( .A1(n7193), .A2(n5700), .A3(n7470), .A4(n7192), .ZN(n7196)
         );
  NAND4_X2 U7560 ( .A1(n7715), .A2(n7714), .A3(n7549), .A4(n7194), .ZN(n7195)
         );
  OAI22_X2 U7561 ( .A1(n7196), .A2(n7195), .B1(n8846), .B2(n4772), .ZN(n3963)
         );
  INV_X4 U7562 ( .A(n8412), .ZN(n7197) );
  XNOR2_X2 U7563 ( .A(n7199), .B(n7198), .ZN(n7202) );
  NAND2_X2 U7564 ( .A1(n7498), .A2(n7412), .ZN(n7200) );
  NAND3_X2 U7565 ( .A1(n8413), .A2(n7204), .A3(n7203), .ZN(aluRes_2[20]) );
  NAND2_X2 U7566 ( .A1(n4781), .A2(memAddr[20]), .ZN(n7206) );
  NAND2_X2 U7567 ( .A1(aluRes_2[20]), .A2(n4791), .ZN(n7205) );
  NAND2_X2 U7568 ( .A1(n7206), .A2(n7205), .ZN(n9159) );
  AOI22_X2 U7569 ( .A1(n4096), .A2(regWrData[1]), .B1(n4132), .B2(n4371), .ZN(
        n7225) );
  NAND2_X2 U7570 ( .A1(n7677), .A2(memAddr[1]), .ZN(n7224) );
  AOI21_X2 U7571 ( .B1(n7209), .B2(n7278), .A(n7208), .ZN(n7222) );
  NAND2_X2 U7572 ( .A1(n4498), .A2(n7562), .ZN(n7221) );
  MUX2_X2 U7573 ( .A(n4731), .B(n4077), .S(n7470), .Z(n7210) );
  NAND2_X2 U7574 ( .A1(n7213), .A2(n7212), .ZN(n7214) );
  NAND2_X2 U7575 ( .A1(n7215), .A2(n7214), .ZN(n7218) );
  AOI211_X2 U7576 ( .C1(n7219), .C2(n7396), .A(n7218), .B(n7217), .ZN(n7220)
         );
  NAND3_X2 U7577 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(n7468) );
  MUX2_X2 U7578 ( .A(n4589), .B(n4205), .S(n4078), .Z(n7471) );
  AOI22_X2 U7579 ( .A1(n7507), .A2(n7468), .B1(n7506), .B2(n7471), .ZN(n7223)
         );
  XNOR2_X2 U7580 ( .A(n7227), .B(n7226), .ZN(n7230) );
  INV_X4 U7581 ( .A(n8455), .ZN(n7229) );
  NAND2_X2 U7582 ( .A1(n8453), .A2(n8454), .ZN(n7228) );
  INV_X4 U7583 ( .A(n7231), .ZN(aluRes_2[16]) );
  NAND2_X2 U7584 ( .A1(memAddr[16]), .A2(n4782), .ZN(n7233) );
  NAND2_X2 U7585 ( .A1(aluRes_2[16]), .A2(n4791), .ZN(n7232) );
  NAND2_X2 U7586 ( .A1(n7233), .A2(n7232), .ZN(n9156) );
  INV_X4 U7587 ( .A(aluRes_2[15]), .ZN(n7234) );
  OAI22_X2 U7588 ( .A1(n4788), .A2(n7234), .B1(n9013), .B2(n4772), .ZN(n9155)
         );
  INV_X4 U7589 ( .A(n7235), .ZN(n7238) );
  INV_X4 U7590 ( .A(n7239), .ZN(n7372) );
  INV_X4 U7591 ( .A(n7240), .ZN(n7244) );
  AOI22_X2 U7592 ( .A1(n7244), .A2(n7361), .B1(n7243), .B2(n7242), .ZN(n7276)
         );
  NAND2_X2 U7593 ( .A1(n4084), .A2(n7720), .ZN(n7247) );
  XNOR2_X2 U7594 ( .A(n7247), .B(n7337), .ZN(n7335) );
  INV_X4 U7595 ( .A(n7248), .ZN(n7251) );
  XNOR2_X2 U7596 ( .A(n7335), .B(n7333), .ZN(n7353) );
  NAND2_X2 U7597 ( .A1(n7721), .A2(n4085), .ZN(n7349) );
  XNOR2_X2 U7598 ( .A(n7353), .B(n7349), .ZN(n7351) );
  XNOR2_X2 U7599 ( .A(n7351), .B(n7350), .ZN(n7257) );
  INV_X4 U7600 ( .A(n7257), .ZN(n7255) );
  NAND2_X2 U7601 ( .A1(n4100), .A2(n7722), .ZN(n7256) );
  NAND2_X2 U7602 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  NAND2_X2 U7603 ( .A1(n7327), .A2(n7258), .ZN(n7329) );
  INV_X4 U7604 ( .A(n7259), .ZN(n7262) );
  OAI21_X4 U7605 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n7326) );
  XNOR2_X2 U7606 ( .A(n7329), .B(n7326), .ZN(n7347) );
  NAND2_X2 U7607 ( .A1(n7723), .A2(n4108), .ZN(n7346) );
  XNOR2_X2 U7608 ( .A(n7347), .B(n7346), .ZN(n7343) );
  XNOR2_X2 U7609 ( .A(n7343), .B(n7342), .ZN(n7321) );
  NAND2_X2 U7610 ( .A1(n7266), .A2(n8326), .ZN(n7267) );
  NAND2_X2 U7611 ( .A1(n4168), .A2(n7271), .ZN(n7322) );
  OAI211_X2 U7612 ( .C1(n4168), .C2(n7271), .A(n7322), .B(n4078), .ZN(n7275)
         );
  NAND2_X2 U7613 ( .A1(n7273), .A2(n7272), .ZN(n7274) );
  NAND3_X2 U7614 ( .A1(n7277), .A2(n4784), .A3(n4573), .ZN(n7370) );
  XNOR2_X2 U7615 ( .A(n7372), .B(n7371), .ZN(n7283) );
  NAND2_X2 U7616 ( .A1(n7492), .A2(n7278), .ZN(n7282) );
  NAND2_X2 U7617 ( .A1(n7279), .A2(n8325), .ZN(n7280) );
  AND3_X2 U7618 ( .A1(n8320), .A2(n8319), .A3(n7280), .ZN(n7281) );
  OAI211_X2 U7619 ( .C1(n7615), .C2(n7283), .A(n7282), .B(n7281), .ZN(
        aluRes_2[30]) );
  NAND2_X2 U7620 ( .A1(n4781), .A2(memAddr[30]), .ZN(n7285) );
  NAND2_X2 U7621 ( .A1(aluRes_2[30]), .A2(n4791), .ZN(n7284) );
  NAND2_X2 U7622 ( .A1(n7285), .A2(n7284), .ZN(n9168) );
  XNOR2_X2 U7623 ( .A(n7287), .B(n7286), .ZN(n7290) );
  NAND2_X2 U7624 ( .A1(n7504), .A2(n7412), .ZN(n7288) );
  AOI21_X2 U7625 ( .B1(n7290), .B2(n4794), .A(n7289), .ZN(n7298) );
  INV_X4 U7626 ( .A(n7921), .ZN(n7294) );
  NAND2_X2 U7627 ( .A1(n7291), .A2(n7489), .ZN(n7292) );
  NAND4_X2 U7628 ( .A1(n8339), .A2(n8338), .A3(n7298), .A4(n7297), .ZN(
        aluRes_2[28]) );
  INV_X4 U7629 ( .A(aluRes_2[28]), .ZN(n7300) );
  OAI22_X2 U7630 ( .A1(n4788), .A2(n7300), .B1(n9043), .B2(n4774), .ZN(n3971)
         );
  INV_X4 U7631 ( .A(n8352), .ZN(n7301) );
  XNOR2_X2 U7632 ( .A(n7303), .B(n7302), .ZN(n7306) );
  NAND2_X2 U7633 ( .A1(n7502), .A2(n7412), .ZN(n7304) );
  AOI21_X2 U7634 ( .B1(n7306), .B2(n4794), .A(n7305), .ZN(n7307) );
  NAND3_X2 U7635 ( .A1(n8353), .A2(n7308), .A3(n7307), .ZN(aluRes_2[26]) );
  NAND2_X2 U7636 ( .A1(n4781), .A2(memAddr[26]), .ZN(n7310) );
  NAND2_X2 U7637 ( .A1(aluRes_2[26]), .A2(n4791), .ZN(n7309) );
  NAND2_X2 U7638 ( .A1(n7310), .A2(n7309), .ZN(n9165) );
  INV_X4 U7639 ( .A(n8373), .ZN(n7311) );
  XNOR2_X2 U7640 ( .A(n7313), .B(n7312), .ZN(n7316) );
  NAND2_X2 U7641 ( .A1(n7527), .A2(n7412), .ZN(n7314) );
  NAND3_X2 U7642 ( .A1(n8374), .A2(n7318), .A3(n7317), .ZN(aluRes_2[23]) );
  NAND2_X2 U7643 ( .A1(memAddr[23]), .A2(n4782), .ZN(n7320) );
  NAND2_X2 U7644 ( .A1(aluRes_2[23]), .A2(n4791), .ZN(n7319) );
  NAND2_X2 U7645 ( .A1(n7320), .A2(n7319), .ZN(n9162) );
  INV_X4 U7646 ( .A(n7321), .ZN(n7324) );
  INV_X4 U7647 ( .A(n7322), .ZN(n7323) );
  INV_X4 U7648 ( .A(n7326), .ZN(n7328) );
  XNOR2_X2 U7649 ( .A(n7331), .B(n7330), .ZN(n7332) );
  XNOR2_X2 U7650 ( .A(n7332), .B(n4374), .ZN(n7341) );
  NAND2_X2 U7651 ( .A1(n7721), .A2(n4100), .ZN(n7339) );
  NAND2_X2 U7652 ( .A1(n7720), .A2(n4084), .ZN(n7336) );
  INV_X4 U7653 ( .A(n7333), .ZN(n7334) );
  OAI22_X2 U7654 ( .A1(n7337), .A2(n7336), .B1(n7335), .B2(n7334), .ZN(n7338)
         );
  XNOR2_X2 U7655 ( .A(n7339), .B(n7338), .ZN(n7340) );
  XNOR2_X2 U7656 ( .A(n7341), .B(n7340), .ZN(n7359) );
  NAND2_X2 U7657 ( .A1(n4108), .A2(n7722), .ZN(n7345) );
  NAND2_X2 U7658 ( .A1(n7343), .A2(n7342), .ZN(n7344) );
  XOR2_X2 U7659 ( .A(n7345), .B(n7344), .Z(n7357) );
  INV_X4 U7660 ( .A(n7346), .ZN(n7348) );
  NAND2_X2 U7661 ( .A1(n7348), .A2(n7347), .ZN(n7356) );
  INV_X4 U7662 ( .A(n7349), .ZN(n7352) );
  AOI22_X2 U7663 ( .A1(n7353), .A2(n7352), .B1(n7351), .B2(n7350), .ZN(n7354)
         );
  XNOR2_X2 U7664 ( .A(n7354), .B(n4507), .ZN(n7355) );
  FA_X1 U7665 ( .A(n7357), .B(n7356), .CI(n7355), .S(n7358) );
  XNOR2_X2 U7666 ( .A(n7359), .B(n7358), .ZN(n7369) );
  NAND2_X2 U7667 ( .A1(n7361), .A2(n7360), .ZN(n7367) );
  NAND2_X2 U7668 ( .A1(n7363), .A2(n7243), .ZN(n7366) );
  NAND2_X2 U7669 ( .A1(n7273), .A2(n7364), .ZN(n7365) );
  AOI21_X4 U7670 ( .B1(n4078), .B2(n7369), .A(n7368), .ZN(n7376) );
  NAND2_X2 U7671 ( .A1(n4784), .A2(n4588), .ZN(n7374) );
  XNOR2_X2 U7672 ( .A(n7374), .B(n7373), .ZN(n7375) );
  XNOR2_X2 U7673 ( .A(n7376), .B(n7375), .ZN(n7377) );
  NAND2_X2 U7674 ( .A1(n7377), .A2(n4794), .ZN(n7405) );
  INV_X4 U7675 ( .A(n7429), .ZN(n7378) );
  NAND2_X2 U7676 ( .A1(n7378), .A2(n7489), .ZN(n7404) );
  INV_X4 U7677 ( .A(n7383), .ZN(n7394) );
  AOI211_X2 U7678 ( .C1(n7385), .C2(n8019), .A(n7384), .B(n8488), .ZN(n7389)
         );
  INV_X4 U7679 ( .A(n8378), .ZN(n7387) );
  AOI21_X2 U7680 ( .B1(n7389), .B2(n7388), .A(n4317), .ZN(n7390) );
  AOI21_X2 U7681 ( .B1(n4312), .B2(n7391), .A(n7390), .ZN(n7392) );
  OAI221_X2 U7682 ( .B1(n7394), .B2(n4128), .C1(n8495), .C2(n4736), .A(n7392), 
        .ZN(n7395) );
  MUX2_X2 U7683 ( .A(n7396), .B(n7395), .S(n7430), .Z(n7426) );
  NAND2_X2 U7684 ( .A1(n7426), .A2(n4083), .ZN(n7397) );
  MUX2_X2 U7685 ( .A(n7547), .B(n7397), .S(n4091), .Z(n7398) );
  INV_X4 U7686 ( .A(n7398), .ZN(n7401) );
  OAI22_X2 U7687 ( .A1(n4728), .A2(n7399), .B1(n7894), .B2(n8524), .ZN(n7400)
         );
  NAND4_X2 U7688 ( .A1(n7405), .A2(n7404), .A3(n7403), .A4(n7402), .ZN(
        aluRes_2[31]) );
  NAND2_X2 U7689 ( .A1(n4781), .A2(memAddr[31]), .ZN(n7407) );
  NAND2_X2 U7690 ( .A1(aluRes_2[31]), .A2(n4791), .ZN(n7406) );
  NAND2_X2 U7691 ( .A1(n7407), .A2(n7406), .ZN(n3976) );
  INV_X4 U7692 ( .A(n8366), .ZN(n7408) );
  INV_X4 U7693 ( .A(n7409), .ZN(n7411) );
  XNOR2_X2 U7694 ( .A(n7411), .B(n7410), .ZN(n7415) );
  NAND2_X2 U7695 ( .A1(n7500), .A2(n7412), .ZN(n7413) );
  NAND3_X2 U7696 ( .A1(n8367), .A2(n7417), .A3(n7416), .ZN(aluRes_2[24]) );
  NAND2_X2 U7697 ( .A1(n4780), .A2(memAddr[24]), .ZN(n7419) );
  NAND2_X2 U7698 ( .A1(aluRes_2[24]), .A2(n4792), .ZN(n7418) );
  NAND2_X2 U7699 ( .A1(n7419), .A2(n7418), .ZN(n9163) );
  AOI22_X2 U7700 ( .A1(n4096), .A2(regWrData[0]), .B1(n4132), .B2(n4372), .ZN(
        n7440) );
  NAND2_X2 U7701 ( .A1(n7677), .A2(memAddr[0]), .ZN(n7439) );
  XNOR2_X2 U7702 ( .A(n7430), .B(n7479), .ZN(n7420) );
  MUX2_X2 U7703 ( .A(n8513), .B(n7420), .S(n9050), .Z(n7421) );
  NAND2_X2 U7704 ( .A1(n8482), .A2(n7421), .ZN(n7436) );
  NAND2_X2 U7705 ( .A1(n7422), .A2(n4731), .ZN(n7424) );
  AOI21_X2 U7706 ( .B1(n8475), .B2(n7426), .A(n7425), .ZN(n7435) );
  NAND2_X2 U7707 ( .A1(n7427), .A2(n7546), .ZN(n7428) );
  NAND4_X2 U7708 ( .A1(n8484), .A2(n7436), .A3(n7435), .A4(n7434), .ZN(n7478)
         );
  MUX2_X2 U7709 ( .A(n4590), .B(n7437), .S(n4078), .Z(n7481) );
  AOI22_X2 U7710 ( .A1(n7507), .A2(n7478), .B1(n7506), .B2(n7481), .ZN(n7438)
         );
  MUX2_X2 U7711 ( .A(n7663), .B(n7441), .S(n4091), .Z(n7444) );
  NAND2_X2 U7712 ( .A1(n7554), .A2(n8018), .ZN(n7445) );
  NAND2_X2 U7713 ( .A1(n7446), .A2(n7445), .ZN(n9193) );
  INV_X4 U7714 ( .A(n7447), .ZN(n7448) );
  NAND2_X2 U7715 ( .A1(n7448), .A2(n4794), .ZN(n7450) );
  MUX2_X2 U7716 ( .A(n7513), .B(n4126), .S(n4091), .Z(n7449) );
  NAND3_X2 U7717 ( .A1(n7450), .A2(n7449), .A3(n4506), .ZN(n9190) );
  NAND2_X2 U7718 ( .A1(n7451), .A2(n4794), .ZN(n7455) );
  INV_X4 U7719 ( .A(n7452), .ZN(n7453) );
  MUX2_X2 U7720 ( .A(n7514), .B(n7453), .S(n4091), .Z(n7454) );
  NAND3_X2 U7721 ( .A1(n7455), .A2(n7454), .A3(n4500), .ZN(n9191) );
  INV_X4 U7722 ( .A(n7456), .ZN(n7457) );
  NAND2_X2 U7723 ( .A1(n7457), .A2(n4794), .ZN(n7461) );
  INV_X4 U7724 ( .A(n7458), .ZN(n7459) );
  MUX2_X2 U7725 ( .A(n7520), .B(n7459), .S(n4091), .Z(n7460) );
  NAND3_X2 U7726 ( .A1(n7461), .A2(n7460), .A3(n4594), .ZN(n9194) );
  INV_X4 U7727 ( .A(n7462), .ZN(n7463) );
  NAND2_X2 U7728 ( .A1(n7463), .A2(n4794), .ZN(n7467) );
  INV_X4 U7729 ( .A(n7464), .ZN(n7465) );
  MUX2_X2 U7730 ( .A(n7515), .B(n7465), .S(n4091), .Z(n7466) );
  NAND3_X2 U7731 ( .A1(n7467), .A2(n7466), .A3(n4586), .ZN(n9192) );
  INV_X4 U7732 ( .A(n7468), .ZN(n7469) );
  MUX2_X2 U7733 ( .A(n7470), .B(n7469), .S(n4091), .Z(n7473) );
  NAND2_X2 U7734 ( .A1(n7471), .A2(n4794), .ZN(n7472) );
  NAND2_X2 U7735 ( .A1(n7473), .A2(n7472), .ZN(n9186) );
  MUX2_X2 U7736 ( .A(n7617), .B(n7474), .S(n4091), .Z(n7477) );
  OAI22_X2 U7737 ( .A1(n7615), .A2(n7475), .B1(n7616), .B2(n4728), .ZN(n7476)
         );
  MUX2_X2 U7738 ( .A(n7479), .B(n7478), .S(n4091), .Z(n7480) );
  INV_X4 U7739 ( .A(n7480), .ZN(n7483) );
  NAND2_X2 U7740 ( .A1(n7481), .A2(n4794), .ZN(n7482) );
  NAND2_X2 U7741 ( .A1(n7483), .A2(n7482), .ZN(aluRes_2[0]) );
  MUX2_X1 U7742 ( .A(wb_dsize_reg_z2[9]), .B(memRdData[9]), .S(n4802), .Z(
        n9059) );
  MUX2_X1 U7743 ( .A(wb_dsize_reg_z2[8]), .B(memRdData[8]), .S(n4795), .Z(
        n9060) );
  MUX2_X1 U7744 ( .A(wb_dsize_reg_z2[7]), .B(memRdData[7]), .S(n4802), .Z(
        n9061) );
  MUX2_X1 U7745 ( .A(wb_dsize_reg_z2[6]), .B(memRdData[6]), .S(n4795), .Z(
        n9062) );
  MUX2_X1 U7746 ( .A(wb_dsize_reg_z2[5]), .B(memRdData[5]), .S(n4802), .Z(
        n9063) );
  MUX2_X1 U7747 ( .A(wb_dsize_reg_z2[4]), .B(memRdData[4]), .S(n4795), .Z(
        n9064) );
  MUX2_X1 U7748 ( .A(wb_dsize_reg_z2[3]), .B(memRdData[3]), .S(n4802), .Z(
        n9065) );
  MUX2_X1 U7749 ( .A(wb_dsize_reg_z2[31]), .B(memRdData[31]), .S(n4795), .Z(
        n9066) );
  MUX2_X1 U7750 ( .A(wb_dsize_reg_z2[30]), .B(memRdData[30]), .S(n4802), .Z(
        n9067) );
  MUX2_X1 U7751 ( .A(wb_dsize_reg_z2[2]), .B(memRdData[2]), .S(n4795), .Z(
        n9068) );
  MUX2_X1 U7752 ( .A(wb_dsize_reg_z2[29]), .B(memRdData[29]), .S(n4802), .Z(
        n9069) );
  MUX2_X1 U7753 ( .A(wb_dsize_reg_z2[28]), .B(memRdData[28]), .S(n4795), .Z(
        n9070) );
  MUX2_X1 U7754 ( .A(wb_dsize_reg_z2[27]), .B(memRdData[27]), .S(n4795), .Z(
        n9071) );
  MUX2_X1 U7755 ( .A(wb_dsize_reg_z2[26]), .B(memRdData[26]), .S(n4795), .Z(
        n9072) );
  MUX2_X1 U7756 ( .A(wb_dsize_reg_z2[25]), .B(memRdData[25]), .S(n4795), .Z(
        n9073) );
  MUX2_X1 U7757 ( .A(wb_dsize_reg_z2[24]), .B(memRdData[24]), .S(n4795), .Z(
        n9074) );
  MUX2_X1 U7758 ( .A(wb_dsize_reg_z2[23]), .B(memRdData[23]), .S(n4795), .Z(
        n9075) );
  MUX2_X1 U7759 ( .A(wb_dsize_reg_z2[22]), .B(memRdData[22]), .S(n4795), .Z(
        n9076) );
  MUX2_X1 U7760 ( .A(wb_dsize_reg_z2[21]), .B(memRdData[21]), .S(n4795), .Z(
        n9077) );
  MUX2_X1 U7761 ( .A(wb_dsize_reg_z2[20]), .B(memRdData[20]), .S(n4795), .Z(
        n9078) );
  MUX2_X1 U7762 ( .A(wb_dsize_reg_z2[1]), .B(memRdData[1]), .S(n4795), .Z(
        n9079) );
  MUX2_X1 U7763 ( .A(wb_dsize_reg_z2[19]), .B(memRdData[19]), .S(n4795), .Z(
        n9080) );
  MUX2_X1 U7764 ( .A(wb_dsize_reg_z2[18]), .B(memRdData[18]), .S(n4796), .Z(
        n9081) );
  MUX2_X1 U7765 ( .A(wb_dsize_reg_z2[17]), .B(memRdData[17]), .S(n4796), .Z(
        n9082) );
  MUX2_X1 U7766 ( .A(wb_dsize_reg_z2[16]), .B(memRdData[16]), .S(n4796), .Z(
        n9083) );
  MUX2_X1 U7767 ( .A(wb_dsize_reg_z2[15]), .B(memRdData[15]), .S(n4796), .Z(
        n9084) );
  MUX2_X1 U7768 ( .A(wb_dsize_reg_z2[14]), .B(memRdData[14]), .S(n4796), .Z(
        n9085) );
  MUX2_X1 U7769 ( .A(wb_dsize_reg_z2[13]), .B(memRdData[13]), .S(n4796), .Z(
        n9086) );
  MUX2_X1 U7770 ( .A(wb_dsize_reg_z2[12]), .B(memRdData[12]), .S(n4796), .Z(
        n9087) );
  MUX2_X1 U7771 ( .A(wb_dsize_reg_z2[11]), .B(memRdData[11]), .S(n4796), .Z(
        n9088) );
  MUX2_X1 U7772 ( .A(wb_dsize_reg_z2[10]), .B(memRdData[10]), .S(n4796), .Z(
        n9089) );
  MUX2_X1 U7773 ( .A(wb_dsize_reg_z2[0]), .B(memRdData[0]), .S(n4796), .Z(
        n9090) );
  MUX2_X1 U7774 ( .A(busA[31]), .B(n4474), .S(n4814), .Z(n9091) );
  MUX2_X1 U7775 ( .A(busA[30]), .B(n4712), .S(n4812), .Z(n9092) );
  MUX2_X1 U7776 ( .A(busA[29]), .B(n4714), .S(n4820), .Z(n9093) );
  MUX2_X1 U7777 ( .A(busA[28]), .B(n4711), .S(n4820), .Z(n9094) );
  MUX2_X1 U7778 ( .A(busA[27]), .B(n4663), .S(n4817), .Z(n9095) );
  MUX2_X1 U7779 ( .A(busA[26]), .B(n4475), .S(n4817), .Z(n9096) );
  MUX2_X1 U7780 ( .A(busA[25]), .B(n4664), .S(n4817), .Z(n9097) );
  MUX2_X1 U7781 ( .A(busA[24]), .B(n4657), .S(n4817), .Z(n9098) );
  MUX2_X1 U7782 ( .A(busA[23]), .B(n4656), .S(n4817), .Z(n9099) );
  MUX2_X1 U7783 ( .A(busA[22]), .B(n4666), .S(n4817), .Z(n9100) );
  MUX2_X1 U7784 ( .A(busA[21]), .B(n4667), .S(n4817), .Z(n9101) );
  MUX2_X1 U7785 ( .A(busA[20]), .B(n4417), .S(n4817), .Z(n9102) );
  MUX2_X1 U7786 ( .A(busA[19]), .B(n4662), .S(n4816), .Z(n9103) );
  MUX2_X1 U7787 ( .A(busA[18]), .B(n4568), .S(n4816), .Z(n9104) );
  MUX2_X1 U7788 ( .A(busA[17]), .B(n4665), .S(n4816), .Z(n9105) );
  MUX2_X1 U7789 ( .A(busA[16]), .B(n4659), .S(n4816), .Z(n9106) );
  MUX2_X1 U7790 ( .A(busA[15]), .B(n4418), .S(n4816), .Z(n9107) );
  MUX2_X1 U7791 ( .A(busA[14]), .B(n4339), .S(n4816), .Z(n9108) );
  MUX2_X1 U7792 ( .A(busA[13]), .B(n4208), .S(n4816), .Z(n9109) );
  MUX2_X1 U7793 ( .A(busA[12]), .B(n4334), .S(n4816), .Z(n9110) );
  MUX2_X1 U7794 ( .A(busA[11]), .B(n4207), .S(n4816), .Z(n9111) );
  MUX2_X1 U7795 ( .A(busA[10]), .B(n4209), .S(n4816), .Z(n9112) );
  MUX2_X1 U7796 ( .A(busA[9]), .B(n4559), .S(n4816), .Z(n9113) );
  MUX2_X1 U7797 ( .A(busA[8]), .B(n4560), .S(n4815), .Z(n9114) );
  MUX2_X1 U7798 ( .A(busA[7]), .B(n4206), .S(n4816), .Z(n9115) );
  MUX2_X1 U7799 ( .A(busA[6]), .B(n4338), .S(n4816), .Z(n9116) );
  MUX2_X1 U7800 ( .A(busA[5]), .B(n4337), .S(n4815), .Z(n9117) );
  MUX2_X1 U7801 ( .A(busA[4]), .B(n4335), .S(n4816), .Z(n9118) );
  MUX2_X1 U7802 ( .A(busA[3]), .B(n4340), .S(n4815), .Z(n9119) );
  MUX2_X1 U7803 ( .A(busA[2]), .B(n4336), .S(n4816), .Z(n9120) );
  MUX2_X1 U7804 ( .A(busA[1]), .B(n4371), .S(n4815), .Z(n9121) );
  MUX2_X1 U7805 ( .A(busA[0]), .B(n4372), .S(n4816), .Z(n9122) );
  MUX2_X1 U7806 ( .A(busB[31]), .B(n4550), .S(n4815), .Z(n9123) );
  MUX2_X1 U7807 ( .A(busB[30]), .B(n4551), .S(n4815), .Z(n9124) );
  MUX2_X1 U7808 ( .A(busB[29]), .B(n4654), .S(n4815), .Z(n9125) );
  MUX2_X1 U7809 ( .A(busB[28]), .B(n4552), .S(n4815), .Z(n9126) );
  MUX2_X1 U7810 ( .A(busB[27]), .B(n4709), .S(n4815), .Z(n9127) );
  MUX2_X1 U7811 ( .A(busB[26]), .B(n4553), .S(n4815), .Z(n9128) );
  MUX2_X1 U7812 ( .A(busB[25]), .B(n4341), .S(n4815), .Z(n9129) );
  MUX2_X1 U7813 ( .A(busB[24]), .B(n4342), .S(n4815), .Z(n9130) );
  MUX2_X1 U7814 ( .A(busB[23]), .B(n4333), .S(n4814), .Z(n9131) );
  MUX2_X1 U7815 ( .A(busB[22]), .B(n4706), .S(n4814), .Z(n9132) );
  MUX2_X1 U7816 ( .A(busB[21]), .B(n4705), .S(n4814), .Z(n9133) );
  MUX2_X1 U7817 ( .A(busB[20]), .B(n4653), .S(n4814), .Z(n9134) );
  MUX2_X1 U7818 ( .A(busB[19]), .B(n4710), .S(n4814), .Z(n9135) );
  MUX2_X1 U7819 ( .A(busB[18]), .B(n4708), .S(n4814), .Z(n9136) );
  MUX2_X1 U7820 ( .A(busB[17]), .B(n4343), .S(n4814), .Z(n9137) );
  MUX2_X1 U7821 ( .A(busB[16]), .B(n4344), .S(n4814), .Z(n9138) );
  MUX2_X1 U7822 ( .A(busB[15]), .B(n4652), .S(n4815), .Z(n9139) );
  MUX2_X1 U7823 ( .A(busB[14]), .B(n4671), .S(n4812), .Z(n9140) );
  MUX2_X1 U7824 ( .A(busB[13]), .B(n4669), .S(n4812), .Z(n9141) );
  MUX2_X1 U7825 ( .A(busB[12]), .B(n4707), .S(n4812), .Z(n9142) );
  MUX2_X1 U7826 ( .A(busB[11]), .B(n4715), .S(n4812), .Z(n9143) );
  MUX2_X1 U7827 ( .A(busB[10]), .B(n4704), .S(n4812), .Z(n9144) );
  MUX2_X1 U7828 ( .A(busB[9]), .B(n4345), .S(n4812), .Z(n9145) );
  MUX2_X1 U7829 ( .A(busB[8]), .B(n4346), .S(n4812), .Z(n9146) );
  MUX2_X1 U7830 ( .A(busB[7]), .B(n4668), .S(n4812), .Z(n9147) );
  MUX2_X1 U7831 ( .A(busB[6]), .B(n4655), .S(n4812), .Z(n9148) );
  MUX2_X1 U7832 ( .A(busB[5]), .B(n4660), .S(n4812), .Z(n9149) );
  MUX2_X1 U7833 ( .A(busB[4]), .B(n4713), .S(n4813), .Z(n9150) );
  MUX2_X1 U7834 ( .A(busB[3]), .B(n4658), .S(n4813), .Z(n9151) );
  MUX2_X1 U7835 ( .A(busB[2]), .B(n4661), .S(n4813), .Z(n9152) );
  MUX2_X1 U7836 ( .A(busB[1]), .B(n4347), .S(n4813), .Z(n9153) );
  MUX2_X1 U7837 ( .A(busB[0]), .B(n4348), .S(n4813), .Z(n9154) );
  MUX2_X1 U7838 ( .A(op0_1), .B(op0_2), .S(n4813), .Z(n9178) );
  MUX2_X1 U7839 ( .A(n7614), .B(n4628), .S(n4813), .Z(n9179) );
  INV_X1 U7840 ( .A(n7618), .ZN(n9180) );
  AOI221_X1 U7841 ( .B1(n4794), .B2(n7619), .C1(n7620), .C2(n4729), .A(n7621), 
        .ZN(n7618) );
  MUX2_X1 U7842 ( .A(n7622), .B(n7623), .S(n4130), .Z(n7621) );
  INV_X1 U7843 ( .A(n7624), .ZN(n9181) );
  AOI221_X1 U7844 ( .B1(n7625), .B2(n4794), .C1(n4729), .C2(n7626), .A(n7627), 
        .ZN(n7624) );
  MUX2_X1 U7845 ( .A(n7628), .B(n7629), .S(n4091), .Z(n7627) );
  OAI221_X1 U7846 ( .B1(n7615), .B2(n7630), .C1(n7631), .C2(n4728), .A(n7632), 
        .ZN(n9182) );
  INV_X1 U7847 ( .A(n7633), .ZN(n7632) );
  MUX2_X1 U7848 ( .A(n7634), .B(n7635), .S(n4091), .Z(n7633) );
  INV_X1 U7849 ( .A(n7636), .ZN(n7630) );
  OAI221_X1 U7850 ( .B1(n7615), .B2(n7637), .C1(n4728), .C2(n7638), .A(n7639), 
        .ZN(n9184) );
  INV_X1 U7851 ( .A(n7640), .ZN(n7639) );
  MUX2_X1 U7852 ( .A(n7641), .B(n7642), .S(n4091), .Z(n7640) );
  INV_X1 U7853 ( .A(n7643), .ZN(n9185) );
  AOI221_X1 U7854 ( .B1(n7644), .B2(n4794), .C1(n4729), .C2(n7645), .A(n7646), 
        .ZN(n7643) );
  MUX2_X1 U7855 ( .A(n7647), .B(n7648), .S(n4130), .Z(n7646) );
  AOI21_X1 U7856 ( .B1(n7572), .B2(n7649), .A(n4537), .ZN(n9187) );
  INV_X1 U7857 ( .A(n7650), .ZN(n9188) );
  AOI221_X1 U7858 ( .B1(n7651), .B2(n4794), .C1(n7652), .C2(n4729), .A(n7653), 
        .ZN(n7650) );
  INV_X1 U7859 ( .A(n7654), .ZN(n9189) );
  AOI221_X1 U7860 ( .B1(n4794), .B2(n7508), .C1(n7554), .C2(n6981), .A(n7655), 
        .ZN(n7654) );
  NAND2_X1 U7861 ( .A1(n7667), .A2(n7668), .ZN(n3975) );
  NAND2_X1 U7862 ( .A1(n7673), .A2(n4804), .ZN(n7672) );
  MUX2_X1 U7863 ( .A(n7674), .B(n4805), .S(n7538), .Z(n7673) );
  AOI222_X1 U7864 ( .A1(n7677), .A2(memAddr[7]), .B1(n4132), .B2(n4206), .C1(
        n4096), .C2(regWrData[7]), .ZN(n7667) );
  NAND2_X1 U7865 ( .A1(n7678), .A2(n7679), .ZN(n3972) );
  AOI222_X1 U7866 ( .A1(n7565), .A2(n7620), .B1(n7506), .B2(n7619), .C1(n7507), 
        .C2(n7622), .ZN(n7679) );
  NAND2_X1 U7867 ( .A1(n7680), .A2(n7681), .ZN(n7622) );
  NAND2_X1 U7868 ( .A1(n7684), .A2(n4804), .ZN(n7683) );
  MUX2_X1 U7869 ( .A(n7674), .B(n4805), .S(n7536), .Z(n7684) );
  XOR2_X1 U7870 ( .A(n7688), .B(n7689), .Z(n7619) );
  AOI222_X1 U7871 ( .A1(n7677), .A2(memAddr[11]), .B1(n4132), .B2(n4207), .C1(
        n4096), .C2(regWrData[11]), .ZN(n7678) );
  NAND2_X1 U7872 ( .A1(n7690), .A2(n7691), .ZN(n3970) );
  AOI222_X1 U7873 ( .A1(n7565), .A2(n7692), .B1(n7506), .B2(n7636), .C1(n7507), 
        .C2(n7635), .ZN(n7691) );
  NAND2_X1 U7874 ( .A1(n7693), .A2(n7694), .ZN(n7635) );
  NAND2_X1 U7875 ( .A1(n7698), .A2(n4804), .ZN(n7697) );
  MUX2_X1 U7876 ( .A(n4805), .B(n7674), .S(n7696), .Z(n7698) );
  XOR2_X1 U7877 ( .A(n7701), .B(n7702), .Z(n7636) );
  AOI222_X1 U7878 ( .A1(n7677), .A2(memAddr[13]), .B1(n4132), .B2(n4208), .C1(
        n4096), .C2(regWrData[13]), .ZN(n7690) );
  NAND2_X1 U7879 ( .A1(n7703), .A2(n7704), .ZN(n3966) );
  AOI222_X1 U7880 ( .A1(n7565), .A2(n7645), .B1(n7506), .B2(n7644), .C1(n7507), 
        .C2(n7647), .ZN(n7704) );
  NAND2_X1 U7881 ( .A1(n7708), .A2(n4804), .ZN(n7707) );
  MUX2_X1 U7882 ( .A(n7674), .B(n4805), .S(n7550), .Z(n7708) );
  XOR2_X1 U7883 ( .A(n7710), .B(n7711), .Z(n7644) );
  INV_X1 U7884 ( .A(n7712), .ZN(n7645) );
  AOI222_X1 U7885 ( .A1(n7677), .A2(memAddr[10]), .B1(n4132), .B2(n4209), .C1(
        n4096), .C2(regWrData[10]), .ZN(n7703) );
  NOR4_X1 U7886 ( .A1(n7716), .A2(n7717), .A3(n7718), .A4(n7719), .ZN(n7715)
         );
  NAND4_X1 U7887 ( .A1(n7547), .A2(n7528), .A3(n7504), .A4(n7503), .ZN(n7719)
         );
  OR4_X1 U7888 ( .A1(n7720), .A2(n7721), .A3(n7722), .A4(n7723), .ZN(n7718) );
  NAND4_X1 U7889 ( .A1(n7527), .A2(n7529), .A3(n7499), .A4(n7498), .ZN(n7717)
         );
  NAND4_X1 U7890 ( .A1(n7497), .A2(n7496), .A3(n7495), .A4(n7494), .ZN(n7716)
         );
  NOR4_X1 U7891 ( .A1(n7724), .A2(n7725), .A3(n7661), .A4(n7663), .ZN(n7714)
         );
  MUX2_X1 U7892 ( .A(n7727), .B(n4545), .S(n4813), .Z(n3898) );
  OAI21_X1 U7893 ( .B1(n7728), .B2(n4611), .A(n4809), .ZN(n3894) );
  INV_X1 U7894 ( .A(n7729), .ZN(n3893) );
  AOI22_X1 U7895 ( .A1(n4811), .A2(n4275), .B1(instruction[31]), .B2(n4806), 
        .ZN(n7729) );
  OAI22_X1 U7896 ( .A1(n7728), .A2(n8959), .B1(n7730), .B2(n4808), .ZN(n3892)
         );
  INV_X1 U7897 ( .A(instruction[30]), .ZN(n7730) );
  INV_X1 U7898 ( .A(n7731), .ZN(n3891) );
  AOI22_X1 U7899 ( .A1(n4811), .A2(n4119), .B1(instruction[29]), .B2(n4806), 
        .ZN(n7731) );
  OAI22_X1 U7900 ( .A1(n8845), .A2(n4824), .B1(n4119), .B2(n7733), .ZN(n3890)
         );
  INV_X1 U7901 ( .A(n7734), .ZN(n3889) );
  AOI22_X1 U7902 ( .A1(n4811), .A2(n4538), .B1(instruction[28]), .B2(n4806), 
        .ZN(n7734) );
  INV_X1 U7903 ( .A(n7735), .ZN(n3888) );
  AOI22_X1 U7904 ( .A1(n4811), .A2(n4120), .B1(instruction[27]), .B2(n4806), 
        .ZN(n7735) );
  MUX2_X1 U7905 ( .A(n7736), .B(n4629), .S(n4813), .Z(n3887) );
  NOR2_X1 U7906 ( .A1(n7737), .A2(n7738), .ZN(n7736) );
  MUX2_X1 U7907 ( .A(n7739), .B(n4630), .S(n4813), .Z(n3886) );
  NOR2_X1 U7908 ( .A1(n8959), .A2(n7740), .ZN(n7739) );
  INV_X1 U7909 ( .A(n7741), .ZN(n3885) );
  AOI22_X1 U7910 ( .A1(n4811), .A2(op0_1), .B1(instruction[26]), .B2(n4806), 
        .ZN(n7741) );
  OAI221_X1 U7911 ( .B1(n8954), .B2(n7733), .C1(n8842), .C2(n4824), .A(n7742), 
        .ZN(n3882) );
  OAI221_X1 U7912 ( .B1(n4323), .B2(n7733), .C1(n8841), .C2(n4824), .A(n7742), 
        .ZN(n3881) );
  NAND4_X1 U7913 ( .A1(n7743), .A2(n7744), .A3(n4538), .A4(n4119), .ZN(n7742)
         );
  INV_X1 U7914 ( .A(n7733), .ZN(n7743) );
  OAI22_X1 U7915 ( .A1(n8964), .A2(n4824), .B1(n7610), .B2(n7745), .ZN(n3880)
         );
  OAI22_X1 U7916 ( .A1(n8840), .A2(n4824), .B1(n7611), .B2(n7745), .ZN(n3879)
         );
  OAI22_X1 U7917 ( .A1(n8839), .A2(n4824), .B1(n7612), .B2(n7745), .ZN(n3878)
         );
  OAI21_X1 U7918 ( .B1(n8838), .B2(n4822), .A(n7746), .ZN(n3877) );
  INV_X1 U7919 ( .A(n7747), .ZN(n7746) );
  MUX2_X1 U7920 ( .A(n7748), .B(n4452), .S(n4813), .Z(n3876) );
  NAND3_X1 U7921 ( .A1(n7749), .A2(n7750), .A3(n7751), .ZN(n7748) );
  INV_X1 U7922 ( .A(n7752), .ZN(n3875) );
  AOI22_X1 U7923 ( .A1(n4811), .A2(rs1[4]), .B1(instruction[25]), .B2(n4806), 
        .ZN(n7752) );
  INV_X1 U7924 ( .A(n7753), .ZN(n3874) );
  AOI22_X1 U7925 ( .A1(n4811), .A2(rs1[3]), .B1(instruction[24]), .B2(n4806), 
        .ZN(n7753) );
  INV_X1 U7926 ( .A(n7754), .ZN(n3873) );
  AOI22_X1 U7927 ( .A1(n4811), .A2(rs1[2]), .B1(instruction[23]), .B2(n4806), 
        .ZN(n7754) );
  INV_X1 U7928 ( .A(n7755), .ZN(n3872) );
  AOI22_X1 U7929 ( .A1(n4811), .A2(rs1[1]), .B1(instruction[22]), .B2(n4806), 
        .ZN(n7755) );
  INV_X1 U7930 ( .A(n7756), .ZN(n3871) );
  AOI22_X1 U7931 ( .A1(n4811), .A2(rs1[0]), .B1(instruction[21]), .B2(n4806), 
        .ZN(n7756) );
  INV_X1 U7932 ( .A(n7757), .ZN(n3870) );
  AOI22_X1 U7933 ( .A1(n4811), .A2(n4332), .B1(instruction[20]), .B2(n4806), 
        .ZN(n7757) );
  INV_X1 U7934 ( .A(n7758), .ZN(n3869) );
  AOI22_X1 U7935 ( .A1(n4811), .A2(n4548), .B1(instruction[19]), .B2(n4806), 
        .ZN(n7758) );
  INV_X1 U7936 ( .A(n7759), .ZN(n3868) );
  AOI22_X1 U7937 ( .A1(n4811), .A2(n4547), .B1(instruction[18]), .B2(n4806), 
        .ZN(n7759) );
  INV_X1 U7938 ( .A(n7760), .ZN(n3867) );
  AOI22_X1 U7939 ( .A1(n4811), .A2(n4328), .B1(instruction[17]), .B2(n4806), 
        .ZN(n7760) );
  INV_X1 U7940 ( .A(n7761), .ZN(n3866) );
  AOI22_X1 U7941 ( .A1(n4811), .A2(n4329), .B1(instruction[16]), .B2(n4806), 
        .ZN(n7761) );
  INV_X1 U7942 ( .A(n7762), .ZN(n3865) );
  AOI22_X1 U7943 ( .A1(n4811), .A2(n4546), .B1(instruction[15]), .B2(n4806), 
        .ZN(n7762) );
  OAI22_X1 U7944 ( .A1(n8837), .A2(n4824), .B1(n8945), .B2(n7745), .ZN(n3864)
         );
  OAI221_X1 U7945 ( .B1(n8945), .B2(n7763), .C1(n8836), .C2(n4824), .A(n7764), 
        .ZN(n3863) );
  OAI211_X1 U7946 ( .C1(n7610), .C2(n7763), .A(n7765), .B(n7766), .ZN(n3862)
         );
  AOI22_X1 U7947 ( .A1(n7747), .A2(n4332), .B1(n4813), .B2(n4557), .ZN(n7766)
         );
  OAI211_X1 U7948 ( .C1(n7611), .C2(n7763), .A(n7765), .B(n7767), .ZN(n3861)
         );
  AOI22_X1 U7949 ( .A1(n7747), .A2(n4547), .B1(n4814), .B2(n4138), .ZN(n7767)
         );
  OAI211_X1 U7950 ( .C1(n7612), .C2(n7763), .A(n7765), .B(n7768), .ZN(n3860)
         );
  AOI22_X1 U7951 ( .A1(n7747), .A2(n4329), .B1(n4815), .B2(n4564), .ZN(n7768)
         );
  OAI22_X1 U7952 ( .A1(n7728), .A2(n8835), .B1(n7769), .B2(n4807), .ZN(n3859)
         );
  INV_X1 U7953 ( .A(instruction[14]), .ZN(n7769) );
  OAI221_X1 U7954 ( .B1(n8835), .B2(n7763), .C1(n8834), .C2(n4824), .A(n7764), 
        .ZN(n3858) );
  OAI22_X1 U7955 ( .A1(n8833), .A2(n4824), .B1(n8835), .B2(n7745), .ZN(n3857)
         );
  OAI22_X1 U7956 ( .A1(n7728), .A2(n8832), .B1(n7770), .B2(n4807), .ZN(n3856)
         );
  INV_X1 U7957 ( .A(instruction[13]), .ZN(n7770) );
  OAI221_X1 U7958 ( .B1(n8832), .B2(n7763), .C1(n8831), .C2(n4824), .A(n7764), 
        .ZN(n3855) );
  OAI22_X1 U7959 ( .A1(n8830), .A2(n4824), .B1(n8832), .B2(n7745), .ZN(n3854)
         );
  OAI22_X1 U7960 ( .A1(n7728), .A2(n8829), .B1(n7771), .B2(n4807), .ZN(n3853)
         );
  INV_X1 U7961 ( .A(instruction[12]), .ZN(n7771) );
  OAI221_X1 U7962 ( .B1(n8829), .B2(n7763), .C1(n8966), .C2(n4824), .A(n7764), 
        .ZN(n3852) );
  OAI22_X1 U7963 ( .A1(n8828), .A2(n4824), .B1(n8829), .B2(n7745), .ZN(n3851)
         );
  OAI22_X1 U7964 ( .A1(n7728), .A2(n8827), .B1(n7772), .B2(n4807), .ZN(n3850)
         );
  INV_X1 U7965 ( .A(instruction[11]), .ZN(n7772) );
  OAI221_X1 U7966 ( .B1(n8827), .B2(n7763), .C1(n8826), .C2(n4824), .A(n7764), 
        .ZN(n3849) );
  OAI22_X1 U7967 ( .A1(n8825), .A2(n4824), .B1(n8827), .B2(n7745), .ZN(n3848)
         );
  OAI22_X1 U7968 ( .A1(n7728), .A2(n8824), .B1(n7773), .B2(n4807), .ZN(n3847)
         );
  INV_X1 U7969 ( .A(instruction[10]), .ZN(n7773) );
  OAI221_X1 U7970 ( .B1(n8824), .B2(n7763), .C1(n8968), .C2(n4824), .A(n7764), 
        .ZN(n3846) );
  OAI22_X1 U7971 ( .A1(n8823), .A2(n4824), .B1(n8824), .B2(n7745), .ZN(n3845)
         );
  OAI22_X1 U7972 ( .A1(n7728), .A2(n8934), .B1(n7774), .B2(n4807), .ZN(n3844)
         );
  INV_X1 U7973 ( .A(instruction[9]), .ZN(n7774) );
  OAI22_X1 U7974 ( .A1(n8822), .A2(n4824), .B1(n8934), .B2(n7745), .ZN(n3843)
         );
  OAI211_X1 U7975 ( .C1(n8934), .C2(n7763), .A(n7765), .B(n7775), .ZN(n3842)
         );
  AOI22_X1 U7976 ( .A1(n7747), .A2(rs1[4]), .B1(n4816), .B2(n4565), .ZN(n7775)
         );
  OAI22_X1 U7977 ( .A1(n7728), .A2(n8936), .B1(n7776), .B2(n4807), .ZN(n3841)
         );
  INV_X1 U7978 ( .A(instruction[8]), .ZN(n7776) );
  OAI22_X1 U7979 ( .A1(n8960), .A2(n4822), .B1(n8936), .B2(n7745), .ZN(n3840)
         );
  OAI211_X1 U7980 ( .C1(n8936), .C2(n7763), .A(n7765), .B(n7777), .ZN(n3839)
         );
  AOI22_X1 U7981 ( .A1(n7747), .A2(rs1[3]), .B1(n4816), .B2(n4566), .ZN(n7777)
         );
  OAI22_X1 U7982 ( .A1(n4810), .A2(n8938), .B1(n7778), .B2(n4807), .ZN(n3838)
         );
  INV_X1 U7983 ( .A(instruction[7]), .ZN(n7778) );
  OAI22_X1 U7984 ( .A1(n8821), .A2(n4822), .B1(n8938), .B2(n7745), .ZN(n3837)
         );
  OAI211_X1 U7985 ( .C1(n8938), .C2(n7763), .A(n7765), .B(n7779), .ZN(n3836)
         );
  AOI22_X1 U7986 ( .A1(n7747), .A2(rs1[2]), .B1(n4817), .B2(n4467), .ZN(n7779)
         );
  OAI22_X1 U7987 ( .A1(n4810), .A2(n8940), .B1(n7780), .B2(n4807), .ZN(n3835)
         );
  INV_X1 U7988 ( .A(instruction[6]), .ZN(n7780) );
  OAI22_X1 U7989 ( .A1(n8962), .A2(n4822), .B1(n8940), .B2(n7745), .ZN(n3834)
         );
  OAI211_X1 U7990 ( .C1(n8940), .C2(n7763), .A(n7765), .B(n7781), .ZN(n3833)
         );
  AOI22_X1 U7991 ( .A1(n7747), .A2(rs1[1]), .B1(n4818), .B2(n4407), .ZN(n7781)
         );
  INV_X1 U7992 ( .A(n7782), .ZN(n3832) );
  AOI22_X1 U7993 ( .A1(n4811), .A2(n4525), .B1(instruction[5]), .B2(n4806), 
        .ZN(n7782) );
  OAI22_X1 U7994 ( .A1(n8820), .A2(n4822), .B1(n8956), .B2(n7745), .ZN(n3831)
         );
  OAI211_X1 U7995 ( .C1(n8956), .C2(n7763), .A(n7765), .B(n7783), .ZN(n3830)
         );
  AOI22_X1 U7996 ( .A1(n7747), .A2(rs1[0]), .B1(n4812), .B2(n4175), .ZN(n7783)
         );
  INV_X1 U7997 ( .A(n7784), .ZN(n3829) );
  MUX2_X1 U7998 ( .A(n7785), .B(n4091), .S(n4814), .Z(n7784) );
  INV_X1 U7999 ( .A(n7786), .ZN(n3828) );
  AOI22_X1 U8000 ( .A1(n4811), .A2(n4318), .B1(instruction[3]), .B2(n4806), 
        .ZN(n7786) );
  OAI22_X1 U8001 ( .A1(n8819), .A2(n4822), .B1(n8955), .B2(n7745), .ZN(n3827)
         );
  OAI211_X1 U8002 ( .C1(n8955), .C2(n7763), .A(n7765), .B(n7787), .ZN(n3826)
         );
  AOI22_X1 U8003 ( .A1(n7747), .A2(n4548), .B1(n4819), .B2(n4176), .ZN(n7787)
         );
  MUX2_X1 U8004 ( .A(n7788), .B(n4133), .S(n4814), .Z(n3825) );
  NAND3_X1 U8005 ( .A1(n7789), .A2(n7790), .A3(n7791), .ZN(n7788) );
  AOI21_X1 U8006 ( .B1(n7792), .B2(n7793), .A(n7794), .ZN(n7791) );
  INV_X1 U8007 ( .A(n7795), .ZN(n3824) );
  AOI22_X1 U8008 ( .A1(n4811), .A2(n4524), .B1(instruction[1]), .B2(n4806), 
        .ZN(n7795) );
  OAI22_X1 U8009 ( .A1(n8818), .A2(n4822), .B1(n8944), .B2(n7745), .ZN(n3823)
         );
  OAI211_X1 U8010 ( .C1(n8944), .C2(n7763), .A(n7765), .B(n7797), .ZN(n3822)
         );
  AOI22_X1 U8011 ( .A1(n7747), .A2(n4328), .B1(n4820), .B2(n4567), .ZN(n7797)
         );
  NAND4_X1 U8012 ( .A1(n7796), .A2(n7800), .A3(n7801), .A4(n4546), .ZN(n7764)
         );
  NAND3_X1 U8013 ( .A1(op0_1), .A2(n8957), .A3(n7802), .ZN(n7801) );
  OAI21_X1 U8014 ( .B1(n7803), .B2(n7804), .A(n4321), .ZN(n7800) );
  NOR2_X1 U8015 ( .A1(n7805), .A2(n4826), .ZN(n7796) );
  MUX2_X1 U8016 ( .A(n7806), .B(n4136), .S(n4815), .Z(n3821) );
  MUX2_X1 U8017 ( .A(n7807), .B(setInv_2), .S(n4815), .Z(n3820) );
  OAI211_X1 U8018 ( .C1(n7808), .C2(n7809), .A(n7810), .B(n7811), .ZN(n7807)
         );
  NOR2_X1 U8019 ( .A1(n7812), .A2(n7813), .ZN(n7811) );
  NOR3_X1 U8020 ( .A1(n7814), .A2(n7815), .A3(n4539), .ZN(n7813) );
  AOI21_X1 U8021 ( .B1(n7744), .B2(n4538), .A(n7816), .ZN(n7808) );
  OAI222_X1 U8022 ( .A1(n7817), .A2(n7818), .B1(n8945), .B2(n7819), .C1(n4533), 
        .C2(n4824), .ZN(n3819) );
  OAI222_X1 U8023 ( .A1(n7820), .A2(n7818), .B1(n8835), .B2(n7819), .C1(n4324), 
        .C2(n4824), .ZN(n3818) );
  OAI222_X1 U8024 ( .A1(n7821), .A2(n7818), .B1(n8832), .B2(n7819), .C1(n4095), 
        .C2(n4824), .ZN(n3817) );
  OAI222_X1 U8025 ( .A1(n7822), .A2(n7818), .B1(n8829), .B2(n7819), .C1(n4322), 
        .C2(n4824), .ZN(n3816) );
  OAI222_X1 U8026 ( .A1(n7823), .A2(n7818), .B1(n8827), .B2(n7819), .C1(n4094), 
        .C2(n4824), .ZN(n3815) );
  NAND2_X1 U8027 ( .A1(n4821), .A2(n7824), .ZN(n7819) );
  NAND3_X1 U8028 ( .A1(n7825), .A2(n4822), .A3(n7826), .ZN(n7818) );
  INV_X1 U8029 ( .A(n7824), .ZN(n7826) );
  OAI21_X1 U8030 ( .B1(n7610), .B2(n7827), .A(n7828), .ZN(n7824) );
  NAND3_X1 U8031 ( .A1(n4275), .A2(n4119), .A3(n8959), .ZN(n7825) );
  MUX2_X1 U8032 ( .A(n7829), .B(n4121), .S(n4815), .Z(n3814) );
  INV_X1 U8033 ( .A(n7830), .ZN(n3813) );
  MUX2_X1 U8034 ( .A(n7609), .B(n9055), .S(n4796), .Z(n7830) );
  INV_X1 U8035 ( .A(n7831), .ZN(n3812) );
  MUX2_X1 U8036 ( .A(n7608), .B(n8989), .S(n4797), .Z(n7831) );
  INV_X1 U8037 ( .A(n7832), .ZN(n3811) );
  MUX2_X1 U8038 ( .A(n7607), .B(n9000), .S(n4797), .Z(n7832) );
  MUX2_X1 U8039 ( .A(n4621), .B(memAddr[10]), .S(n4797), .Z(n3810) );
  MUX2_X1 U8040 ( .A(n4622), .B(memAddr[11]), .S(n4797), .Z(n3809) );
  INV_X1 U8041 ( .A(n7833), .ZN(n3808) );
  MUX2_X1 U8042 ( .A(n7606), .B(n9009), .S(n4797), .Z(n7833) );
  INV_X1 U8043 ( .A(n7834), .ZN(n3807) );
  MUX2_X1 U8044 ( .A(n7605), .B(n9013), .S(n4797), .Z(n7834) );
  INV_X1 U8045 ( .A(n7835), .ZN(n3806) );
  MUX2_X1 U8046 ( .A(n7604), .B(n9016), .S(n4797), .Z(n7835) );
  INV_X1 U8047 ( .A(n7836), .ZN(n3805) );
  MUX2_X1 U8048 ( .A(n7603), .B(n9024), .S(n4797), .Z(n7836) );
  INV_X1 U8049 ( .A(n7837), .ZN(n3804) );
  MUX2_X1 U8050 ( .A(n7602), .B(n9031), .S(n4797), .Z(n7837) );
  MUX2_X1 U8051 ( .A(n4613), .B(memAddr[24]), .S(n4797), .Z(n3803) );
  INV_X1 U8052 ( .A(n7838), .ZN(n3802) );
  MUX2_X1 U8053 ( .A(n7600), .B(n9039), .S(n4797), .Z(n7838) );
  INV_X1 U8054 ( .A(n7839), .ZN(n3801) );
  MUX2_X1 U8055 ( .A(n7599), .B(n9043), .S(n4798), .Z(n7839) );
  MUX2_X1 U8056 ( .A(n4623), .B(memAddr[30]), .S(n4798), .Z(n3800) );
  MUX2_X1 U8057 ( .A(n4614), .B(memAddr[31]), .S(n4798), .Z(n3799) );
  MUX2_X1 U8058 ( .A(dSize[0]), .B(n4633), .S(n7840), .Z(n3767) );
  MUX2_X1 U8059 ( .A(n4105), .B(dSize[0]), .S(n4798), .Z(n3766) );
  MUX2_X1 U8060 ( .A(dSize[1]), .B(n4634), .S(n7840), .Z(n3765) );
  NOR2_X1 U8061 ( .A1(n4892), .A2(n4789), .ZN(n7840) );
  MUX2_X1 U8062 ( .A(n4086), .B(dSize[1]), .S(n4798), .Z(n3764) );
  MUX2_X1 U8063 ( .A(rd[0]), .B(rd_3[0]), .S(n4798), .Z(n3760) );
  MUX2_X1 U8064 ( .A(rd[1]), .B(rd_3[1]), .S(n4798), .Z(n3758) );
  MUX2_X1 U8065 ( .A(rd[2]), .B(rd_3[2]), .S(n4798), .Z(n3756) );
  MUX2_X1 U8066 ( .A(rd[4]), .B(rd_3[4]), .S(n4798), .Z(n3749) );
  MUX2_X1 U8067 ( .A(rd[3]), .B(rd_3[3]), .S(n4798), .Z(n3747) );
  MUX2_X1 U8068 ( .A(n4104), .B(n4631), .S(n4798), .Z(n3744) );
  NOR2_X1 U8069 ( .A1(n8838), .A2(n4789), .ZN(n3741) );
  MUX2_X1 U8070 ( .A(n4670), .B(n4362), .S(n4799), .Z(n3739) );
  OAI221_X1 U8071 ( .B1(n7594), .B2(n4828), .C1(n7612), .C2(n4820), .A(n7841), 
        .ZN(n3695) );
  OAI22_X1 U8072 ( .A1(n8944), .A2(n4820), .B1(n8800), .B2(n4827), .ZN(n3693)
         );
  OAI221_X1 U8073 ( .B1(n7592), .B2(n4828), .C1(n7611), .C2(n4820), .A(n7841), 
        .ZN(n3691) );
  OAI22_X1 U8074 ( .A1(n8955), .A2(n4820), .B1(n8915), .B2(n4828), .ZN(n3689)
         );
  OAI221_X1 U8075 ( .B1(n7590), .B2(n4828), .C1(n7610), .C2(n4820), .A(n7841), 
        .ZN(n3687) );
  OAI22_X1 U8076 ( .A1(n8956), .A2(n4820), .B1(n8926), .B2(n4828), .ZN(n3685)
         );
  OAI22_X1 U8077 ( .A1(n4818), .A2(n4323), .B1(n8929), .B2(n4828), .ZN(n3683)
         );
  OAI22_X1 U8078 ( .A1(n8954), .A2(n4820), .B1(n8930), .B2(n4828), .ZN(n3681)
         );
  OAI22_X1 U8079 ( .A1(n8957), .A2(n4820), .B1(n8928), .B2(n4828), .ZN(n3679)
         );
  OAI22_X1 U8080 ( .A1(n8953), .A2(n4820), .B1(n8918), .B2(n4828), .ZN(n3677)
         );
  OAI22_X1 U8081 ( .A1(n8959), .A2(n4820), .B1(n8917), .B2(n4828), .ZN(n3675)
         );
  OAI22_X1 U8082 ( .A1(n8791), .A2(n4827), .B1(n8953), .B2(n7733), .ZN(n3673)
         );
  OAI221_X1 U8083 ( .B1(n4119), .B2(n7733), .C1(n4827), .C2(n4610), .A(n7842), 
        .ZN(n3671) );
  OAI21_X1 U8084 ( .B1(n7843), .B2(n7844), .A(n4822), .ZN(n7842) );
  OAI221_X1 U8085 ( .B1(n4321), .B2(n7785), .C1(n7827), .C2(n7845), .A(n7828), 
        .ZN(n7844) );
  AOI21_X1 U8086 ( .B1(n7793), .B2(n7846), .A(n7803), .ZN(n7828) );
  INV_X1 U8087 ( .A(n7789), .ZN(n7803) );
  AND2_X1 U8088 ( .A1(n7847), .A2(n7845), .ZN(n7846) );
  OAI21_X1 U8089 ( .B1(n7848), .B2(n4525), .A(n4129), .ZN(n7847) );
  NOR3_X1 U8090 ( .A1(n4318), .A2(n7611), .A3(n7814), .ZN(n7848) );
  INV_X1 U8091 ( .A(n7849), .ZN(n7814) );
  INV_X1 U8092 ( .A(n7850), .ZN(n7845) );
  NAND3_X1 U8093 ( .A1(n4129), .A2(n4525), .A3(n7793), .ZN(n7785) );
  NAND4_X1 U8094 ( .A1(n7751), .A2(n7750), .A3(n7851), .A4(n7852), .ZN(n7843)
         );
  NAND3_X1 U8095 ( .A1(n4823), .A2(n4275), .A3(n8959), .ZN(n7733) );
  OAI221_X1 U8096 ( .B1(n4820), .B2(n7854), .C1(n4827), .C2(n4650), .A(n7841), 
        .ZN(n3668) );
  NOR3_X1 U8097 ( .A1(n7804), .A2(n7855), .A3(n7856), .ZN(n7854) );
  NAND4_X1 U8098 ( .A1(n7857), .A2(n7751), .A3(n7827), .A4(n7740), .ZN(n7804)
         );
  NAND4_X1 U8099 ( .A1(n7858), .A2(n7749), .A3(n7827), .A4(n7740), .ZN(n7751)
         );
  NAND2_X1 U8100 ( .A1(n7816), .A2(n7859), .ZN(n7858) );
  NAND2_X1 U8101 ( .A1(n7860), .A2(n7861), .ZN(n7857) );
  XOR2_X1 U8102 ( .A(n4532), .B(n4137), .Z(n7862) );
  INV_X1 U8103 ( .A(n7863), .ZN(n3664) );
  MUX2_X1 U8104 ( .A(n8789), .B(n8788), .S(n4815), .Z(n7863) );
  MUX2_X1 U8105 ( .A(reg31Val_0[0]), .B(reg31Val_3[0]), .S(n4799), .Z(n3662)
         );
  OAI21_X1 U8106 ( .B1(n4829), .B2(n4087), .A(n7763), .ZN(n3661) );
  OAI22_X1 U8107 ( .A1(n4817), .A2(n4528), .B1(n8931), .B2(n4828), .ZN(n3660)
         );
  OAI22_X1 U8108 ( .A1(n4819), .A2(n4529), .B1(n8786), .B2(n4828), .ZN(n3658)
         );
  OAI22_X1 U8109 ( .A1(n4818), .A2(n4527), .B1(n8919), .B2(n4828), .ZN(n3656)
         );
  OAI22_X1 U8110 ( .A1(n4819), .A2(n4531), .B1(n8920), .B2(n4828), .ZN(n3654)
         );
  OAI22_X1 U8111 ( .A1(n4816), .A2(n4530), .B1(n8921), .B2(n4828), .ZN(n3652)
         );
  OAI22_X1 U8112 ( .A1(n8904), .A2(n4820), .B1(n8922), .B2(n4829), .ZN(n3650)
         );
  OAI22_X1 U8113 ( .A1(n8905), .A2(n4820), .B1(n8924), .B2(n4828), .ZN(n3648)
         );
  OAI22_X1 U8114 ( .A1(n8906), .A2(n4820), .B1(n8923), .B2(n4829), .ZN(n3646)
         );
  OAI22_X1 U8115 ( .A1(n8907), .A2(n4820), .B1(n8925), .B2(n4828), .ZN(n3644)
         );
  OAI22_X1 U8116 ( .A1(n8908), .A2(n4820), .B1(n8909), .B2(n4829), .ZN(n3642)
         );
  OAI22_X1 U8117 ( .A1(n8945), .A2(n4820), .B1(n8911), .B2(n4829), .ZN(n3640)
         );
  OAI22_X1 U8118 ( .A1(n8835), .A2(n4820), .B1(n8912), .B2(n4829), .ZN(n3638)
         );
  OAI22_X1 U8119 ( .A1(n8832), .A2(n4820), .B1(n8913), .B2(n4829), .ZN(n3636)
         );
  OAI22_X1 U8120 ( .A1(n8829), .A2(n4817), .B1(n8914), .B2(n4829), .ZN(n3634)
         );
  OAI22_X1 U8121 ( .A1(n8827), .A2(n4820), .B1(n8772), .B2(n4829), .ZN(n3632)
         );
  OAI22_X1 U8122 ( .A1(n8824), .A2(n4820), .B1(n8770), .B2(n4829), .ZN(n3630)
         );
  OAI22_X1 U8123 ( .A1(n8934), .A2(n4818), .B1(n8768), .B2(n4829), .ZN(n3628)
         );
  OAI22_X1 U8124 ( .A1(n8936), .A2(n4817), .B1(n8766), .B2(n4829), .ZN(n3626)
         );
  OAI22_X1 U8125 ( .A1(n8938), .A2(n4819), .B1(n8910), .B2(n4829), .ZN(n3624)
         );
  OAI22_X1 U8126 ( .A1(n8940), .A2(n4819), .B1(n8927), .B2(n4829), .ZN(n3622)
         );
  OAI22_X1 U8127 ( .A1(n4818), .A2(n4611), .B1(n4361), .B2(n4829), .ZN(n3620)
         );
  OAI22_X1 U8128 ( .A1(n9057), .A2(n4827), .B1(n7864), .B2(n7865), .ZN(n3618)
         );
  NAND4_X1 U8129 ( .A1(n7493), .A2(n7866), .A3(n7867), .A4(n7868), .ZN(n7865)
         );
  XNOR2_X1 U8130 ( .A(rd_3[0]), .B(rs2[0]), .ZN(n7868) );
  XNOR2_X1 U8131 ( .A(rd_3[4]), .B(rs2[4]), .ZN(n7867) );
  NAND4_X1 U8132 ( .A1(n7869), .A2(n7870), .A3(n7871), .A4(n7872), .ZN(n7864)
         );
  XNOR2_X1 U8133 ( .A(rd_3[3]), .B(rs2[3]), .ZN(n7871) );
  XNOR2_X1 U8134 ( .A(rd_3[2]), .B(rs2[2]), .ZN(n7870) );
  XNOR2_X1 U8135 ( .A(rd_3[1]), .B(rs2[1]), .ZN(n7869) );
  OAI22_X1 U8136 ( .A1(n9052), .A2(n4827), .B1(n7873), .B2(n7874), .ZN(n3617)
         );
  NAND4_X1 U8137 ( .A1(n7875), .A2(n7876), .A3(n7877), .A4(n7878), .ZN(n7874)
         );
  XNOR2_X1 U8138 ( .A(n4530), .B(n4319), .ZN(n7878) );
  XNOR2_X1 U8139 ( .A(n4531), .B(n4093), .ZN(n7877) );
  XNOR2_X1 U8140 ( .A(n4527), .B(n4081), .ZN(n7876) );
  XNOR2_X1 U8141 ( .A(n4528), .B(n4320), .ZN(n7875) );
  NAND4_X1 U8142 ( .A1(n7879), .A2(n7493), .A3(n7866), .A4(n7880), .ZN(n7873)
         );
  XNOR2_X1 U8143 ( .A(n4529), .B(n4092), .ZN(n7879) );
  OAI22_X1 U8144 ( .A1(n9058), .A2(n4827), .B1(n7881), .B2(n7872), .ZN(n3616)
         );
  OAI22_X1 U8145 ( .A1(n9053), .A2(n4827), .B1(n7881), .B2(n7880), .ZN(n3614)
         );
  XOR2_X1 U8146 ( .A(n7883), .B(n7884), .Z(n7882) );
  NOR2_X1 U8147 ( .A1(n8901), .A2(n4532), .ZN(n7883) );
  INV_X1 U8148 ( .A(n7885), .ZN(n3610) );
  MUX2_X1 U8149 ( .A(n8760), .B(n8759), .S(n4817), .Z(n7885) );
  MUX2_X1 U8150 ( .A(reg31Val_0[1]), .B(reg31Val_3[1]), .S(n4799), .Z(n3608)
         );
  INV_X1 U8151 ( .A(n7886), .ZN(n3605) );
  MUX2_X1 U8152 ( .A(n7588), .B(n9028), .S(n4799), .Z(n7886) );
  XOR2_X1 U8153 ( .A(n7889), .B(n7890), .Z(n7651) );
  MUX2_X1 U8154 ( .A(n4615), .B(memAddr[9]), .S(n4799), .Z(n3602) );
  AOI22_X1 U8155 ( .A1(n7897), .A2(n7895), .B1(n7492), .B2(n7898), .ZN(n7893)
         );
  NAND3_X1 U8156 ( .A1(n4091), .A2(n7896), .A3(n7899), .ZN(n7897) );
  MUX2_X1 U8157 ( .A(n7674), .B(n7894), .S(n7518), .Z(n7899) );
  AOI22_X1 U8158 ( .A1(n7491), .A2(n7699), .B1(n7490), .B2(n7700), .ZN(n7892)
         );
  AOI22_X1 U8159 ( .A1(n7489), .A2(n7900), .B1(n4729), .B2(n7901), .ZN(n7891)
         );
  MUX2_X1 U8160 ( .A(n4616), .B(memAddr[17]), .S(n4799), .Z(n3599) );
  NAND2_X1 U8161 ( .A1(n7902), .A2(n7903), .ZN(n3597) );
  AOI222_X1 U8162 ( .A1(n7565), .A2(n7626), .B1(n7506), .B2(n7625), .C1(n7507), 
        .C2(n7629), .ZN(n7903) );
  NAND2_X1 U8163 ( .A1(n7904), .A2(n7905), .ZN(n7629) );
  NAND2_X1 U8164 ( .A1(n7908), .A2(n4804), .ZN(n7907) );
  MUX2_X1 U8165 ( .A(n7674), .B(n4805), .S(n7537), .Z(n7908) );
  XNOR2_X1 U8166 ( .A(n7909), .B(n7910), .ZN(n7625) );
  INV_X1 U8167 ( .A(n7911), .ZN(n7626) );
  AOI222_X1 U8168 ( .A1(n7677), .A2(memAddr[12]), .B1(n4132), .B2(n4334), .C1(
        n4096), .C2(regWrData[12]), .ZN(n7902) );
  MUX2_X1 U8169 ( .A(n4624), .B(memAddr[12]), .S(n4799), .Z(n3596) );
  MUX2_X1 U8170 ( .A(n4625), .B(memAddr[29]), .S(n4799), .Z(n3593) );
  MUX2_X1 U8171 ( .A(n4617), .B(memAddr[8]), .S(n4799), .Z(n3590) );
  MUX2_X1 U8172 ( .A(n4618), .B(memAddr[25]), .S(n4799), .Z(n3587) );
  MUX2_X1 U8173 ( .A(n4619), .B(memAddr[18]), .S(n4799), .Z(n3584) );
  MUX2_X1 U8174 ( .A(n4626), .B(memAddr[27]), .S(n4800), .Z(n3581) );
  NAND2_X1 U8175 ( .A1(n7915), .A2(n7916), .ZN(n3579) );
  NAND2_X1 U8176 ( .A1(n7920), .A2(n4804), .ZN(n7919) );
  MUX2_X1 U8177 ( .A(n4805), .B(n7674), .S(n7918), .Z(n7920) );
  AOI222_X1 U8178 ( .A1(n7677), .A2(memAddr[4]), .B1(n4132), .B2(n4335), .C1(
        n4096), .C2(regWrData[4]), .ZN(n7915) );
  MUX2_X1 U8179 ( .A(n4620), .B(memAddr[4]), .S(n4800), .Z(n3578) );
  INV_X1 U8180 ( .A(n7922), .ZN(n3575) );
  MUX2_X1 U8181 ( .A(n7581), .B(n9022), .S(n4800), .Z(n7922) );
  INV_X1 U8182 ( .A(n7923), .ZN(n3573) );
  MUX2_X1 U8183 ( .A(n7924), .B(n8756), .S(n7666), .Z(n7923) );
  OAI22_X1 U8184 ( .A1(n8755), .A2(n4810), .B1(n4807), .B2(n7924), .ZN(n3572)
         );
  INV_X1 U8185 ( .A(n7926), .ZN(n3571) );
  MUX2_X1 U8186 ( .A(n8755), .B(n8754), .S(n4817), .Z(n7926) );
  INV_X1 U8187 ( .A(n7927), .ZN(n3569) );
  MUX2_X1 U8188 ( .A(n7928), .B(n8753), .S(n7666), .Z(n7927) );
  OAI22_X1 U8189 ( .A1(n8752), .A2(n4810), .B1(n4809), .B2(n7928), .ZN(n3568)
         );
  INV_X1 U8190 ( .A(n7929), .ZN(n3567) );
  MUX2_X1 U8191 ( .A(n8752), .B(n8751), .S(n4817), .Z(n7929) );
  INV_X1 U8192 ( .A(n7930), .ZN(n3565) );
  MUX2_X1 U8193 ( .A(n7931), .B(n8750), .S(n7666), .Z(n7930) );
  OAI22_X1 U8194 ( .A1(n8749), .A2(n4810), .B1(n4808), .B2(n7931), .ZN(n3564)
         );
  INV_X1 U8195 ( .A(n7932), .ZN(n3563) );
  MUX2_X1 U8196 ( .A(n8749), .B(n8748), .S(n4818), .Z(n7932) );
  INV_X1 U8197 ( .A(n7933), .ZN(n3561) );
  MUX2_X1 U8198 ( .A(n7934), .B(n8747), .S(n7666), .Z(n7933) );
  OAI22_X1 U8199 ( .A1(n8746), .A2(n4810), .B1(n4809), .B2(n7934), .ZN(n3560)
         );
  INV_X1 U8200 ( .A(n7935), .ZN(n3559) );
  MUX2_X1 U8201 ( .A(n8746), .B(n8745), .S(n4818), .Z(n7935) );
  INV_X1 U8202 ( .A(n7936), .ZN(n3557) );
  MUX2_X1 U8203 ( .A(n7937), .B(n8744), .S(n7666), .Z(n7936) );
  OAI22_X1 U8204 ( .A1(n8743), .A2(n4810), .B1(n4808), .B2(n7937), .ZN(n3556)
         );
  INV_X1 U8205 ( .A(n7938), .ZN(n3555) );
  MUX2_X1 U8206 ( .A(n8743), .B(n8742), .S(n4818), .Z(n7938) );
  INV_X1 U8207 ( .A(n7939), .ZN(n3553) );
  MUX2_X1 U8208 ( .A(n7940), .B(n8741), .S(n7666), .Z(n7939) );
  OAI22_X1 U8209 ( .A1(n8740), .A2(n4810), .B1(n4809), .B2(n7940), .ZN(n3552)
         );
  INV_X1 U8210 ( .A(n7941), .ZN(n3551) );
  MUX2_X1 U8211 ( .A(n8740), .B(n8739), .S(n4818), .Z(n7941) );
  INV_X1 U8212 ( .A(n7942), .ZN(n3549) );
  MUX2_X1 U8213 ( .A(n7943), .B(n8738), .S(n7666), .Z(n7942) );
  OAI22_X1 U8214 ( .A1(n8737), .A2(n4810), .B1(n4808), .B2(n7943), .ZN(n3548)
         );
  INV_X1 U8215 ( .A(n7944), .ZN(n3547) );
  MUX2_X1 U8216 ( .A(n8737), .B(n8736), .S(n4818), .Z(n7944) );
  INV_X1 U8217 ( .A(n7945), .ZN(n3545) );
  MUX2_X1 U8218 ( .A(n8735), .B(n7946), .S(n7487), .Z(n7945) );
  OAI22_X1 U8219 ( .A1(n8734), .A2(n4810), .B1(n4809), .B2(n7946), .ZN(n3544)
         );
  INV_X1 U8220 ( .A(n7947), .ZN(n3543) );
  MUX2_X1 U8221 ( .A(n8734), .B(n8733), .S(n4818), .Z(n7947) );
  INV_X1 U8222 ( .A(n7948), .ZN(n3541) );
  MUX2_X1 U8223 ( .A(n8732), .B(n7949), .S(n4793), .Z(n7948) );
  OAI22_X1 U8224 ( .A1(n8731), .A2(n4810), .B1(n4809), .B2(n7949), .ZN(n3540)
         );
  INV_X1 U8225 ( .A(n7950), .ZN(n3539) );
  MUX2_X1 U8226 ( .A(n8731), .B(n8730), .S(n4818), .Z(n7950) );
  INV_X1 U8227 ( .A(n7951), .ZN(n3537) );
  MUX2_X1 U8228 ( .A(n8729), .B(n7952), .S(n4793), .Z(n7951) );
  OAI22_X1 U8229 ( .A1(n8728), .A2(n4810), .B1(n4809), .B2(n7952), .ZN(n3536)
         );
  INV_X1 U8230 ( .A(n7953), .ZN(n3535) );
  MUX2_X1 U8231 ( .A(n8728), .B(n8727), .S(n4818), .Z(n7953) );
  INV_X1 U8232 ( .A(n7954), .ZN(n3533) );
  MUX2_X1 U8233 ( .A(n8726), .B(n4271), .S(n4793), .Z(n7954) );
  OAI22_X1 U8234 ( .A1(n8725), .A2(n4810), .B1(n4809), .B2(n4271), .ZN(n3532)
         );
  INV_X1 U8235 ( .A(n7955), .ZN(n3531) );
  MUX2_X1 U8236 ( .A(n8725), .B(n8724), .S(n4818), .Z(n7955) );
  MUX2_X1 U8237 ( .A(reg31Val_0[30]), .B(n7956), .S(n4800), .Z(n3529) );
  XOR2_X1 U8238 ( .A(n4526), .B(n7957), .Z(n7956) );
  NAND2_X1 U8239 ( .A1(n7958), .A2(n7959), .ZN(n3527) );
  NAND2_X1 U8240 ( .A1(n7961), .A2(n4804), .ZN(n7960) );
  MUX2_X1 U8241 ( .A(n7674), .B(n4805), .S(n7548), .Z(n7961) );
  AOI222_X1 U8242 ( .A1(n7677), .A2(memAddr[2]), .B1(n4132), .B2(n4336), .C1(
        n4096), .C2(regWrData[2]), .ZN(n7958) );
  INV_X1 U8243 ( .A(n7963), .ZN(n3526) );
  MUX2_X1 U8244 ( .A(n7580), .B(n8991), .S(n4800), .Z(n7963) );
  INV_X1 U8245 ( .A(n7964), .ZN(n3522) );
  MUX2_X1 U8246 ( .A(n8723), .B(n8722), .S(n4818), .Z(n7964) );
  MUX2_X1 U8247 ( .A(reg31Val_0[2]), .B(n8900), .S(n4800), .Z(n3520) );
  NAND2_X1 U8248 ( .A1(n7965), .A2(n7966), .ZN(n3518) );
  NAND2_X1 U8249 ( .A1(n7970), .A2(n4804), .ZN(n7969) );
  MUX2_X1 U8250 ( .A(n7674), .B(n4805), .S(n7539), .Z(n7970) );
  AOI222_X1 U8251 ( .A1(n7677), .A2(memAddr[5]), .B1(n4132), .B2(n4337), .C1(
        n4096), .C2(regWrData[5]), .ZN(n7965) );
  INV_X1 U8252 ( .A(n7973), .ZN(n3517) );
  MUX2_X1 U8253 ( .A(n7579), .B(n8996), .S(n4800), .Z(n7973) );
  NAND2_X1 U8254 ( .A1(n7974), .A2(n7975), .ZN(n3515) );
  NAND2_X1 U8255 ( .A1(n7979), .A2(n4804), .ZN(n7978) );
  MUX2_X1 U8256 ( .A(n7674), .B(n4805), .S(n7540), .Z(n7979) );
  AOI222_X1 U8257 ( .A1(n7677), .A2(memAddr[6]), .B1(n4132), .B2(n4338), .C1(
        n4096), .C2(regWrData[6]), .ZN(n7974) );
  INV_X1 U8258 ( .A(n7981), .ZN(n3514) );
  MUX2_X1 U8259 ( .A(n7578), .B(n8998), .S(n4800), .Z(n7981) );
  OAI211_X1 U8260 ( .C1(n7638), .C2(n7982), .A(n7983), .B(n7984), .ZN(n3512)
         );
  AOI222_X1 U8261 ( .A1(n7677), .A2(memAddr[14]), .B1(n4132), .B2(n4339), .C1(
        n4096), .C2(regWrData[14]), .ZN(n7984) );
  AOI22_X1 U8262 ( .A1(n7506), .A2(n7985), .B1(n7507), .B2(n7642), .ZN(n7983)
         );
  NAND2_X1 U8263 ( .A1(n7986), .A2(n7987), .ZN(n7642) );
  NAND2_X1 U8264 ( .A1(n7990), .A2(n4804), .ZN(n7989) );
  MUX2_X1 U8265 ( .A(n7674), .B(n4805), .S(n7541), .Z(n7990) );
  INV_X1 U8266 ( .A(n7637), .ZN(n7985) );
  XNOR2_X1 U8267 ( .A(n7486), .B(n7991), .ZN(n7637) );
  INV_X1 U8268 ( .A(n7992), .ZN(n3511) );
  MUX2_X1 U8269 ( .A(n7577), .B(n9011), .S(n4800), .Z(n7992) );
  INV_X1 U8270 ( .A(n7993), .ZN(n3509) );
  MUX2_X1 U8271 ( .A(n8719), .B(n7994), .S(n4793), .Z(n7993) );
  OAI22_X1 U8272 ( .A1(n8718), .A2(n4810), .B1(n4808), .B2(n7994), .ZN(n3508)
         );
  INV_X1 U8273 ( .A(n7995), .ZN(n3507) );
  MUX2_X1 U8274 ( .A(n8718), .B(n8717), .S(n4818), .Z(n7995) );
  INV_X1 U8275 ( .A(n7996), .ZN(n3505) );
  MUX2_X1 U8276 ( .A(n8716), .B(n7997), .S(n4793), .Z(n7996) );
  OAI22_X1 U8277 ( .A1(n8715), .A2(n4810), .B1(n4808), .B2(n7997), .ZN(n3504)
         );
  NAND2_X1 U8278 ( .A1(n7998), .A2(n7999), .ZN(n7997) );
  INV_X1 U8279 ( .A(n8001), .ZN(n3503) );
  MUX2_X1 U8280 ( .A(n8715), .B(n8714), .S(n4819), .Z(n8001) );
  INV_X1 U8281 ( .A(n8002), .ZN(n3501) );
  MUX2_X1 U8282 ( .A(n8713), .B(n8003), .S(n4793), .Z(n8002) );
  OAI22_X1 U8283 ( .A1(n8712), .A2(n4810), .B1(n4808), .B2(n8003), .ZN(n3500)
         );
  INV_X1 U8284 ( .A(n8004), .ZN(n3499) );
  MUX2_X1 U8285 ( .A(n8712), .B(n8711), .S(n4819), .Z(n8004) );
  INV_X1 U8286 ( .A(n8005), .ZN(n3497) );
  MUX2_X1 U8287 ( .A(n8710), .B(n8006), .S(n4793), .Z(n8005) );
  OAI22_X1 U8288 ( .A1(n8709), .A2(n7728), .B1(n4808), .B2(n8006), .ZN(n3496)
         );
  NAND2_X1 U8289 ( .A1(n7925), .A2(n8007), .ZN(n8006) );
  INV_X1 U8290 ( .A(n8008), .ZN(n3495) );
  MUX2_X1 U8291 ( .A(n8709), .B(n8708), .S(n4819), .Z(n8008) );
  INV_X1 U8292 ( .A(n8009), .ZN(n3493) );
  MUX2_X1 U8293 ( .A(n8707), .B(n8010), .S(n4793), .Z(n8009) );
  OAI22_X1 U8294 ( .A1(n8706), .A2(n7728), .B1(n4808), .B2(n8010), .ZN(n3492)
         );
  INV_X1 U8295 ( .A(n8011), .ZN(n3491) );
  MUX2_X1 U8296 ( .A(n8706), .B(n8705), .S(n4819), .Z(n8011) );
  MUX2_X1 U8297 ( .A(reg31Val_0[29]), .B(n8012), .S(n4800), .Z(n3489) );
  XNOR2_X1 U8298 ( .A(n8013), .B(n4534), .ZN(n8012) );
  MUX2_X1 U8299 ( .A(reg31Val_0[28]), .B(n8014), .S(n4800), .Z(n3488) );
  XNOR2_X1 U8300 ( .A(n8856), .B(n8015), .ZN(n8014) );
  NAND2_X1 U8301 ( .A1(n8016), .A2(n8017), .ZN(n3486) );
  NAND2_X1 U8302 ( .A1(n8021), .A2(n4804), .ZN(n8020) );
  MUX2_X1 U8303 ( .A(n4805), .B(n7674), .S(n8019), .Z(n8021) );
  NAND2_X1 U8304 ( .A1(n7507), .A2(n7562), .ZN(n7982) );
  AOI222_X1 U8305 ( .A1(n7677), .A2(memAddr[3]), .B1(n4132), .B2(n4340), .C1(
        n4096), .C2(regWrData[3]), .ZN(n8016) );
  INV_X1 U8306 ( .A(n8023), .ZN(n3485) );
  MUX2_X1 U8307 ( .A(n7576), .B(n8993), .S(n4801), .Z(n8023) );
  INV_X1 U8308 ( .A(n8024), .ZN(n3483) );
  MUX2_X1 U8309 ( .A(n8704), .B(n8025), .S(n4793), .Z(n8024) );
  OAI22_X1 U8310 ( .A1(n8703), .A2(n7728), .B1(n4808), .B2(n8025), .ZN(n3482)
         );
  INV_X1 U8311 ( .A(n8026), .ZN(n3481) );
  MUX2_X1 U8312 ( .A(n8703), .B(n8702), .S(n4819), .Z(n8026) );
  MUX2_X1 U8313 ( .A(reg31Val_0[3]), .B(n8027), .S(n4801), .Z(n3479) );
  XOR2_X1 U8314 ( .A(n4174), .B(n4109), .Z(n8027) );
  INV_X1 U8315 ( .A(n8028), .ZN(n3478) );
  MUX2_X1 U8316 ( .A(n8701), .B(n8029), .S(n4793), .Z(n8028) );
  OAI22_X1 U8317 ( .A1(n8700), .A2(n7728), .B1(n4808), .B2(n8029), .ZN(n3477)
         );
  INV_X1 U8318 ( .A(n8030), .ZN(n3476) );
  MUX2_X1 U8319 ( .A(n8700), .B(n8699), .S(n4819), .Z(n8030) );
  MUX2_X1 U8320 ( .A(reg31Val_0[4]), .B(n8031), .S(n4801), .Z(n3474) );
  XOR2_X1 U8321 ( .A(n4401), .B(n8032), .Z(n8031) );
  INV_X1 U8322 ( .A(n8033), .ZN(n3472) );
  MUX2_X1 U8323 ( .A(n8698), .B(n8034), .S(n4793), .Z(n8033) );
  OAI22_X1 U8324 ( .A1(n8697), .A2(n7728), .B1(n4808), .B2(n8034), .ZN(n3471)
         );
  INV_X1 U8325 ( .A(n8035), .ZN(n3470) );
  MUX2_X1 U8326 ( .A(n8697), .B(n8696), .S(n4819), .Z(n8035) );
  MUX2_X1 U8327 ( .A(reg31Val_0[5]), .B(n8036), .S(n4801), .Z(n3468) );
  XNOR2_X1 U8328 ( .A(n8037), .B(n4173), .ZN(n8036) );
  INV_X1 U8329 ( .A(n8038), .ZN(n3466) );
  MUX2_X1 U8330 ( .A(n8695), .B(n8039), .S(n7487), .Z(n8038) );
  OAI22_X1 U8331 ( .A1(n8694), .A2(n7728), .B1(n4808), .B2(n8039), .ZN(n3465)
         );
  NAND2_X1 U8332 ( .A1(n8040), .A2(n8041), .ZN(n8039) );
  INV_X1 U8333 ( .A(n8042), .ZN(n3464) );
  MUX2_X1 U8334 ( .A(n8694), .B(n8693), .S(n4819), .Z(n8042) );
  MUX2_X1 U8335 ( .A(reg31Val_0[6]), .B(n8043), .S(n4801), .Z(n3462) );
  XOR2_X1 U8336 ( .A(n4400), .B(n8044), .Z(n8043) );
  INV_X1 U8337 ( .A(n8045), .ZN(n3461) );
  MUX2_X1 U8338 ( .A(n8692), .B(n8046), .S(n7487), .Z(n8045) );
  OAI22_X1 U8339 ( .A1(n8691), .A2(n7728), .B1(n4808), .B2(n8046), .ZN(n3460)
         );
  INV_X1 U8340 ( .A(n8047), .ZN(n3459) );
  MUX2_X1 U8341 ( .A(n8691), .B(n8690), .S(n4819), .Z(n8047) );
  MUX2_X1 U8342 ( .A(reg31Val_0[7]), .B(n8048), .S(n4801), .Z(n3457) );
  XNOR2_X1 U8343 ( .A(n8049), .B(n4172), .ZN(n8048) );
  INV_X1 U8344 ( .A(n8050), .ZN(n3455) );
  MUX2_X1 U8345 ( .A(n8689), .B(n8051), .S(n7487), .Z(n8050) );
  OAI22_X1 U8346 ( .A1(n8688), .A2(n7728), .B1(n4808), .B2(n8051), .ZN(n3454)
         );
  NAND2_X1 U8347 ( .A1(n8052), .A2(n8053), .ZN(n8051) );
  INV_X1 U8348 ( .A(n8054), .ZN(n3453) );
  MUX2_X1 U8349 ( .A(n8688), .B(n8687), .S(n4819), .Z(n8054) );
  MUX2_X1 U8350 ( .A(reg31Val_0[8]), .B(n8055), .S(n4801), .Z(n3451) );
  XOR2_X1 U8351 ( .A(n4399), .B(n8056), .Z(n8055) );
  INV_X1 U8352 ( .A(n8057), .ZN(n3450) );
  MUX2_X1 U8353 ( .A(n8686), .B(n8058), .S(n7487), .Z(n8057) );
  OAI22_X1 U8354 ( .A1(n8685), .A2(n4810), .B1(n4809), .B2(n8058), .ZN(n3449)
         );
  INV_X1 U8355 ( .A(n8059), .ZN(n3448) );
  MUX2_X1 U8356 ( .A(n8685), .B(n8684), .S(n4819), .Z(n8059) );
  MUX2_X1 U8357 ( .A(reg31Val_0[9]), .B(n8060), .S(n4801), .Z(n3446) );
  XNOR2_X1 U8358 ( .A(n8061), .B(n4171), .ZN(n8060) );
  INV_X1 U8359 ( .A(n8062), .ZN(n3444) );
  MUX2_X1 U8360 ( .A(n8683), .B(n8063), .S(n7487), .Z(n8062) );
  OAI22_X1 U8361 ( .A1(n8682), .A2(n7728), .B1(n4809), .B2(n8063), .ZN(n3443)
         );
  NAND2_X1 U8362 ( .A1(n8064), .A2(n8065), .ZN(n8063) );
  INV_X1 U8363 ( .A(n8066), .ZN(n3442) );
  MUX2_X1 U8364 ( .A(n8682), .B(n8681), .S(n4820), .Z(n8066) );
  MUX2_X1 U8365 ( .A(reg31Val_0[10]), .B(n8067), .S(n4801), .Z(n3440) );
  XOR2_X1 U8366 ( .A(n4398), .B(n8068), .Z(n8067) );
  INV_X1 U8367 ( .A(n8069), .ZN(n3439) );
  MUX2_X1 U8368 ( .A(n8680), .B(n8070), .S(n4793), .Z(n8069) );
  OAI22_X1 U8369 ( .A1(n8679), .A2(n7728), .B1(n4809), .B2(n8070), .ZN(n3438)
         );
  INV_X1 U8370 ( .A(n8071), .ZN(n3437) );
  MUX2_X1 U8371 ( .A(n8679), .B(n8678), .S(n4820), .Z(n8071) );
  MUX2_X1 U8372 ( .A(reg31Val_0[11]), .B(n8072), .S(n4801), .Z(n3435) );
  XNOR2_X1 U8373 ( .A(n8073), .B(n4170), .ZN(n8072) );
  INV_X1 U8374 ( .A(n8074), .ZN(n3433) );
  MUX2_X1 U8375 ( .A(n8677), .B(n8075), .S(n7487), .Z(n8074) );
  OAI22_X1 U8376 ( .A1(n8676), .A2(n7728), .B1(n4809), .B2(n8075), .ZN(n3432)
         );
  NAND2_X1 U8377 ( .A1(n8076), .A2(n8077), .ZN(n8075) );
  INV_X1 U8378 ( .A(n8078), .ZN(n3431) );
  MUX2_X1 U8379 ( .A(n8676), .B(n8675), .S(n4820), .Z(n8078) );
  MUX2_X1 U8380 ( .A(reg31Val_0[12]), .B(n8079), .S(n4801), .Z(n3429) );
  XOR2_X1 U8381 ( .A(n4397), .B(n8080), .Z(n8079) );
  INV_X1 U8382 ( .A(n8081), .ZN(n3428) );
  MUX2_X1 U8383 ( .A(n8674), .B(n8082), .S(n7487), .Z(n8081) );
  OAI22_X1 U8384 ( .A1(n8673), .A2(n7728), .B1(n4809), .B2(n8082), .ZN(n3427)
         );
  INV_X1 U8385 ( .A(n8083), .ZN(n3426) );
  MUX2_X1 U8386 ( .A(n8673), .B(n8672), .S(n4820), .Z(n8083) );
  MUX2_X1 U8387 ( .A(reg31Val_0[13]), .B(n8084), .S(n4802), .Z(n3424) );
  XNOR2_X1 U8388 ( .A(n8085), .B(n4277), .ZN(n8084) );
  INV_X1 U8389 ( .A(n8086), .ZN(n3422) );
  MUX2_X1 U8390 ( .A(n8671), .B(n8087), .S(n7487), .Z(n8086) );
  OAI22_X1 U8391 ( .A1(n8670), .A2(n4810), .B1(n4809), .B2(n8087), .ZN(n3421)
         );
  NAND2_X1 U8392 ( .A1(n8000), .A2(n8088), .ZN(n8087) );
  INV_X1 U8393 ( .A(n8089), .ZN(n3420) );
  MUX2_X1 U8394 ( .A(n8670), .B(n8669), .S(n4820), .Z(n8089) );
  MUX2_X1 U8395 ( .A(reg31Val_0[21]), .B(n8090), .S(n4802), .Z(n3418) );
  XNOR2_X1 U8396 ( .A(n8091), .B(n4457), .ZN(n8090) );
  MUX2_X1 U8397 ( .A(reg31Val_0[20]), .B(n8092), .S(n4802), .Z(n3417) );
  XNOR2_X1 U8398 ( .A(n8870), .B(n8093), .ZN(n8092) );
  MUX2_X1 U8399 ( .A(reg31Val_0[19]), .B(n8094), .S(n4802), .Z(n3416) );
  XNOR2_X1 U8400 ( .A(n8095), .B(n4458), .ZN(n8094) );
  MUX2_X1 U8401 ( .A(reg31Val_0[18]), .B(n8096), .S(n4802), .Z(n3415) );
  XNOR2_X1 U8402 ( .A(n8874), .B(n8097), .ZN(n8096) );
  MUX2_X1 U8403 ( .A(reg31Val_0[17]), .B(n8098), .S(n4802), .Z(n3414) );
  XNOR2_X1 U8404 ( .A(n8099), .B(n4459), .ZN(n8098) );
  MUX2_X1 U8405 ( .A(reg31Val_0[16]), .B(n8100), .S(n4802), .Z(n3413) );
  XOR2_X1 U8406 ( .A(n4453), .B(n8101), .Z(n8100) );
  MUX2_X1 U8407 ( .A(reg31Val_0[15]), .B(n8102), .S(n4802), .Z(n3411) );
  XNOR2_X1 U8408 ( .A(n8103), .B(n4276), .ZN(n8102) );
  MUX2_X1 U8409 ( .A(reg31Val_0[14]), .B(n8104), .S(n4802), .Z(n3410) );
  XOR2_X1 U8410 ( .A(n4454), .B(n8105), .Z(n8104) );
  MUX2_X1 U8411 ( .A(reg31Val_0[27]), .B(n8106), .S(n4802), .Z(n3408) );
  XNOR2_X1 U8412 ( .A(n8107), .B(n4535), .ZN(n8106) );
  MUX2_X1 U8413 ( .A(reg31Val_0[26]), .B(n8108), .S(n4802), .Z(n3407) );
  XNOR2_X1 U8414 ( .A(n8859), .B(n8109), .ZN(n8108) );
  MUX2_X1 U8415 ( .A(reg31Val_0[25]), .B(n8110), .S(n4797), .Z(n3405) );
  XNOR2_X1 U8416 ( .A(n8111), .B(n4536), .ZN(n8110) );
  MUX2_X1 U8417 ( .A(reg31Val_0[24]), .B(n8112), .S(n4801), .Z(n3404) );
  XNOR2_X1 U8418 ( .A(n8863), .B(n8113), .ZN(n8112) );
  MUX2_X1 U8419 ( .A(reg31Val_0[23]), .B(n8114), .S(n4801), .Z(n3402) );
  XNOR2_X1 U8420 ( .A(n8115), .B(n4456), .ZN(n8114) );
  MUX2_X1 U8421 ( .A(reg31Val_0[22]), .B(n8117), .S(n4801), .Z(n3400) );
  XNOR2_X1 U8422 ( .A(n8867), .B(n8118), .ZN(n8117) );
  INV_X1 U8423 ( .A(n8119), .ZN(n3397) );
  MUX2_X1 U8424 ( .A(n8665), .B(n8120), .S(n7487), .Z(n8119) );
  OAI22_X1 U8425 ( .A1(n8664), .A2(n4810), .B1(n4809), .B2(n8120), .ZN(n3396)
         );
  INV_X1 U8426 ( .A(n8121), .ZN(n3395) );
  MUX2_X1 U8427 ( .A(n8664), .B(n8663), .S(n4820), .Z(n8121) );
  MUX2_X1 U8428 ( .A(reg31Val_0[31]), .B(n8122), .S(n4801), .Z(n3393) );
  XOR2_X1 U8429 ( .A(n8123), .B(n8851), .Z(n8122) );
  NAND2_X1 U8430 ( .A1(n7957), .A2(n4526), .ZN(n8123) );
  NOR2_X1 U8431 ( .A1(n8013), .A2(n8854), .ZN(n7957) );
  NAND2_X1 U8432 ( .A1(n8015), .A2(n4326), .ZN(n8013) );
  NOR2_X1 U8433 ( .A1(n8107), .A2(n8857), .ZN(n8015) );
  NAND2_X1 U8434 ( .A1(n8109), .A2(n4327), .ZN(n8107) );
  NOR2_X1 U8435 ( .A1(n8111), .A2(n8860), .ZN(n8109) );
  NAND2_X1 U8436 ( .A1(n8113), .A2(n4325), .ZN(n8111) );
  NOR2_X1 U8437 ( .A1(n8115), .A2(n8864), .ZN(n8113) );
  NAND2_X1 U8438 ( .A1(n8118), .A2(n4278), .ZN(n8115) );
  NOR2_X1 U8439 ( .A1(n8091), .A2(n8868), .ZN(n8118) );
  NAND2_X1 U8440 ( .A1(n8093), .A2(n4279), .ZN(n8091) );
  NOR2_X1 U8441 ( .A1(n8095), .A2(n8872), .ZN(n8093) );
  NAND2_X1 U8442 ( .A1(n8097), .A2(n4280), .ZN(n8095) );
  NOR2_X1 U8443 ( .A1(n8099), .A2(n8875), .ZN(n8097) );
  NAND2_X1 U8444 ( .A1(n8101), .A2(n4453), .ZN(n8099) );
  NOR2_X1 U8445 ( .A1(n8103), .A2(n8878), .ZN(n8101) );
  NAND2_X1 U8446 ( .A1(n8105), .A2(n4454), .ZN(n8103) );
  NOR2_X1 U8447 ( .A1(n8085), .A2(n8882), .ZN(n8105) );
  NAND2_X1 U8448 ( .A1(n8080), .A2(n4397), .ZN(n8085) );
  NOR2_X1 U8449 ( .A1(n8073), .A2(n8886), .ZN(n8080) );
  NAND2_X1 U8450 ( .A1(n8068), .A2(n4398), .ZN(n8073) );
  NOR2_X1 U8451 ( .A1(n8061), .A2(n8890), .ZN(n8068) );
  NAND2_X1 U8452 ( .A1(n8056), .A2(n4399), .ZN(n8061) );
  NOR2_X1 U8453 ( .A1(n8049), .A2(n8893), .ZN(n8056) );
  NAND2_X1 U8454 ( .A1(n8044), .A2(n4400), .ZN(n8049) );
  NOR2_X1 U8455 ( .A1(n8037), .A2(n8896), .ZN(n8044) );
  NAND2_X1 U8456 ( .A1(n8032), .A2(n4401), .ZN(n8037) );
  NOR2_X1 U8457 ( .A1(n8847), .A2(n8900), .ZN(n8032) );
  INV_X1 U8458 ( .A(n8124), .ZN(n3382) );
  MUX2_X1 U8459 ( .A(n7575), .B(n9026), .S(n4801), .Z(n8124) );
  OAI22_X1 U8460 ( .A1(n8958), .A2(n4817), .B1(n8916), .B2(n4829), .ZN(n3380)
         );
  OAI22_X1 U8461 ( .A1(n4591), .A2(n4818), .B1(n8652), .B2(n4829), .ZN(n3379)
         );
  NAND4_X1 U8462 ( .A1(n8927), .A2(n8928), .A3(n8929), .A4(n8930), .ZN(n8127)
         );
  NAND4_X1 U8463 ( .A1(n8921), .A2(n8922), .A3(n8920), .A4(n8130), .ZN(n8126)
         );
  AND4_X1 U8464 ( .A1(n8926), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(n8130)
         );
  NAND4_X1 U8465 ( .A1(n8131), .A2(n8132), .A3(n8133), .A4(n8134), .ZN(n8125)
         );
  AND4_X1 U8466 ( .A1(n8919), .A2(n8916), .A3(n8915), .A4(n8914), .ZN(n8134)
         );
  AND3_X1 U8467 ( .A1(n8911), .A2(n8913), .A3(n8912), .ZN(n8133) );
  AND4_X1 U8468 ( .A1(n8910), .A2(n8909), .A3(n8814), .A4(n8800), .ZN(n8132)
         );
  NOR3_X1 U8469 ( .A1(n4131), .A2(n4330), .A3(n4544), .ZN(n8131) );
  OAI21_X1 U8470 ( .B1(n8651), .B2(n4829), .A(n8135), .ZN(n3377) );
  NAND4_X1 U8471 ( .A1(n8136), .A2(n8137), .A3(n8138), .A4(n8139), .ZN(n8135)
         );
  AND4_X1 U8472 ( .A1(n4592), .A2(n8928), .A3(n8930), .A4(n8929), .ZN(n8139)
         );
  AND4_X1 U8473 ( .A1(n8140), .A2(n8770), .A3(n8141), .A4(n8142), .ZN(n8129)
         );
  NOR4_X1 U8474 ( .A1(n8143), .A2(n8144), .A3(n8145), .A4(n8146), .ZN(n8142)
         );
  XNOR2_X1 U8475 ( .A(n4320), .B(rd_2[4]), .ZN(n8146) );
  XNOR2_X1 U8476 ( .A(n4092), .B(rd_2[3]), .ZN(n8145) );
  XOR2_X1 U8477 ( .A(n4081), .B(n4095), .Z(n8144) );
  XNOR2_X1 U8478 ( .A(n4093), .B(rd_2[1]), .ZN(n8143) );
  AND2_X1 U8479 ( .A1(n7866), .A2(n8772), .ZN(n8141) );
  INV_X1 U8480 ( .A(n8147), .ZN(n7866) );
  OAI21_X1 U8481 ( .B1(n8148), .B2(n8149), .A(valid_3), .ZN(n8147) );
  NAND2_X1 U8482 ( .A1(n4319), .A2(n4093), .ZN(n8149) );
  NAND3_X1 U8483 ( .A1(n4092), .A2(n4320), .A3(n4081), .ZN(n8148) );
  XOR2_X1 U8484 ( .A(rd_2[0]), .B(n4319), .Z(n8140) );
  AND4_X1 U8485 ( .A1(n8918), .A2(n4726), .A3(n8917), .A4(n8150), .ZN(n8128)
         );
  NOR3_X1 U8486 ( .A1(n7592), .A2(n8791), .A3(n7594), .ZN(n8150) );
  AND4_X1 U8487 ( .A1(n8151), .A2(n8921), .A3(n8923), .A4(n8922), .ZN(n8138)
         );
  AND4_X1 U8488 ( .A1(n8924), .A2(n8925), .A3(n8926), .A4(n8927), .ZN(n8151)
         );
  AND4_X1 U8489 ( .A1(n8152), .A2(n8912), .A3(n8914), .A4(n8913), .ZN(n8137)
         );
  AND4_X1 U8490 ( .A1(n8915), .A2(n8916), .A3(n8919), .A4(n8920), .ZN(n8152)
         );
  NOR4_X1 U8491 ( .A1(n8153), .A2(n4131), .A3(n4330), .A4(n4544), .ZN(n8136)
         );
  NAND4_X1 U8492 ( .A1(n8800), .A2(n8909), .A3(n8910), .A4(n8911), .ZN(n8153)
         );
  NAND2_X1 U8493 ( .A1(n8917), .A2(n8918), .ZN(n8155) );
  INV_X1 U8494 ( .A(n8156), .ZN(n8154) );
  AOI21_X1 U8495 ( .B1(n7880), .B2(n7872), .A(n8916), .ZN(n8156) );
  NAND4_X1 U8496 ( .A1(n8157), .A2(n8158), .A3(n8159), .A4(n8160), .ZN(n7872)
         );
  NOR3_X1 U8497 ( .A1(n8161), .A2(n8162), .A3(n8163), .ZN(n8160) );
  XNOR2_X1 U8498 ( .A(rd_2[4]), .B(n7817), .ZN(n8163) );
  INV_X1 U8499 ( .A(rs2[4]), .ZN(n7817) );
  XNOR2_X1 U8500 ( .A(rd_2[3]), .B(n7820), .ZN(n8162) );
  INV_X1 U8501 ( .A(rs2[3]), .ZN(n7820) );
  XOR2_X1 U8502 ( .A(rd_2[0]), .B(rs2[0]), .Z(n8161) );
  XOR2_X1 U8503 ( .A(rd_2[2]), .B(n7821), .Z(n8158) );
  INV_X1 U8504 ( .A(rs2[2]), .ZN(n7821) );
  XNOR2_X1 U8505 ( .A(rd_2[1]), .B(rs2[1]), .ZN(n8157) );
  NAND4_X1 U8506 ( .A1(n8164), .A2(n8159), .A3(n8165), .A4(n8166), .ZN(n7880)
         );
  NOR3_X1 U8507 ( .A1(n8167), .A2(n8168), .A3(n8169), .ZN(n8166) );
  XNOR2_X1 U8508 ( .A(n4527), .B(rd_2[2]), .ZN(n8169) );
  XNOR2_X1 U8509 ( .A(n4528), .B(rd_2[4]), .ZN(n8168) );
  XNOR2_X1 U8510 ( .A(n4529), .B(rd_2[3]), .ZN(n8167) );
  XNOR2_X1 U8511 ( .A(n4530), .B(n4094), .ZN(n8165) );
  INV_X1 U8512 ( .A(n8170), .ZN(n8159) );
  OAI21_X1 U8513 ( .B1(n8171), .B2(n8172), .A(valid_2), .ZN(n8170) );
  NAND2_X1 U8514 ( .A1(n4094), .A2(n4322), .ZN(n8172) );
  NAND3_X1 U8515 ( .A1(n4324), .A2(n4533), .A3(n4095), .ZN(n8171) );
  XNOR2_X1 U8516 ( .A(n4531), .B(n4322), .ZN(n8164) );
  OR2_X1 U8517 ( .A1(n4876), .A2(initPC[0]), .ZN(n3371) );
  NAND2_X1 U8518 ( .A1(initPC[0]), .A2(n4890), .ZN(n3370) );
  OR2_X1 U8519 ( .A1(n4867), .A2(initPC[1]), .ZN(n3369) );
  NAND2_X1 U8520 ( .A1(initPC[1]), .A2(n4889), .ZN(n3368) );
  OR2_X1 U8521 ( .A1(n4866), .A2(initPC[19]), .ZN(n3367) );
  NAND2_X1 U8522 ( .A1(initPC[19]), .A2(n4888), .ZN(n3366) );
  OR2_X1 U8523 ( .A1(n4865), .A2(initPC[20]), .ZN(n3365) );
  NAND2_X1 U8524 ( .A1(initPC[20]), .A2(n4887), .ZN(n3364) );
  OR2_X1 U8525 ( .A1(n4870), .A2(initPC[21]), .ZN(n3363) );
  NAND2_X1 U8526 ( .A1(initPC[21]), .A2(n4886), .ZN(n3362) );
  OR2_X1 U8527 ( .A1(n4869), .A2(initPC[23]), .ZN(n3361) );
  NAND2_X1 U8528 ( .A1(initPC[23]), .A2(n4885), .ZN(n3360) );
  OR2_X1 U8529 ( .A1(n4868), .A2(initPC[24]), .ZN(n3359) );
  NAND2_X1 U8530 ( .A1(initPC[24]), .A2(n4885), .ZN(n3358) );
  OR2_X1 U8531 ( .A1(n4873), .A2(initPC[25]), .ZN(n3357) );
  NAND2_X1 U8532 ( .A1(initPC[25]), .A2(n4884), .ZN(n3356) );
  OR2_X1 U8533 ( .A1(n4872), .A2(initPC[26]), .ZN(n3355) );
  NAND2_X1 U8534 ( .A1(initPC[26]), .A2(n4883), .ZN(n3354) );
  OR2_X1 U8535 ( .A1(n4871), .A2(initPC[27]), .ZN(n3353) );
  NAND2_X1 U8536 ( .A1(initPC[27]), .A2(n4882), .ZN(n3352) );
  OR2_X1 U8537 ( .A1(n4875), .A2(initPC[28]), .ZN(n3351) );
  NAND2_X1 U8538 ( .A1(initPC[28]), .A2(n4881), .ZN(n3350) );
  OR2_X1 U8539 ( .A1(n4874), .A2(initPC[29]), .ZN(n3349) );
  NAND2_X1 U8540 ( .A1(initPC[29]), .A2(n4880), .ZN(n3348) );
  OR2_X1 U8541 ( .A1(n4864), .A2(initPC[30]), .ZN(n3347) );
  NAND2_X1 U8542 ( .A1(initPC[30]), .A2(n4879), .ZN(n3346) );
  OR2_X1 U8543 ( .A1(n4863), .A2(initPC[2]), .ZN(n3345) );
  NAND2_X1 U8544 ( .A1(initPC[2]), .A2(n4891), .ZN(n3344) );
  OR2_X1 U8545 ( .A1(n4862), .A2(initPC[15]), .ZN(n3343) );
  NAND2_X1 U8546 ( .A1(initPC[15]), .A2(n4890), .ZN(n3342) );
  OR2_X1 U8547 ( .A1(n4861), .A2(initPC[16]), .ZN(n3341) );
  NAND2_X1 U8548 ( .A1(initPC[16]), .A2(n4889), .ZN(n3340) );
  OR2_X1 U8549 ( .A1(n4861), .A2(initPC[17]), .ZN(n3339) );
  NAND2_X1 U8550 ( .A1(initPC[17]), .A2(n4888), .ZN(n3338) );
  OR2_X1 U8551 ( .A1(n4860), .A2(initPC[18]), .ZN(n3337) );
  NAND2_X1 U8552 ( .A1(initPC[18]), .A2(n4887), .ZN(n3336) );
  OR2_X1 U8553 ( .A1(n4857), .A2(initPC[22]), .ZN(n3335) );
  NAND2_X1 U8554 ( .A1(initPC[22]), .A2(n4886), .ZN(n3334) );
  OR2_X1 U8555 ( .A1(n4856), .A2(initPC[3]), .ZN(n3333) );
  NAND2_X1 U8556 ( .A1(initPC[3]), .A2(n4885), .ZN(n3332) );
  OR2_X1 U8557 ( .A1(n4878), .A2(initPC[4]), .ZN(n3331) );
  NAND2_X1 U8558 ( .A1(initPC[4]), .A2(n4888), .ZN(n3330) );
  OR2_X1 U8559 ( .A1(n4878), .A2(initPC[5]), .ZN(n3329) );
  NAND2_X1 U8560 ( .A1(initPC[5]), .A2(n4892), .ZN(n3328) );
  OR2_X1 U8561 ( .A1(n4878), .A2(initPC[6]), .ZN(n3327) );
  NAND2_X1 U8562 ( .A1(initPC[6]), .A2(n4892), .ZN(n3326) );
  OR2_X1 U8563 ( .A1(n4878), .A2(initPC[7]), .ZN(n3325) );
  NAND2_X1 U8564 ( .A1(initPC[7]), .A2(n4891), .ZN(n3324) );
  OR2_X1 U8565 ( .A1(n4878), .A2(initPC[8]), .ZN(n3323) );
  NAND2_X1 U8566 ( .A1(initPC[8]), .A2(n4892), .ZN(n3322) );
  OR2_X1 U8567 ( .A1(n4878), .A2(initPC[9]), .ZN(n3321) );
  NAND2_X1 U8568 ( .A1(initPC[9]), .A2(n4892), .ZN(n3320) );
  OR2_X1 U8569 ( .A1(n4878), .A2(initPC[10]), .ZN(n3319) );
  NAND2_X1 U8570 ( .A1(initPC[10]), .A2(n4892), .ZN(n3318) );
  OR2_X1 U8571 ( .A1(n4878), .A2(initPC[11]), .ZN(n3317) );
  NAND2_X1 U8572 ( .A1(initPC[11]), .A2(n4892), .ZN(n3316) );
  OR2_X1 U8573 ( .A1(n4878), .A2(initPC[12]), .ZN(n3315) );
  NAND2_X1 U8574 ( .A1(initPC[12]), .A2(n4892), .ZN(n3314) );
  OR2_X1 U8575 ( .A1(n4878), .A2(initPC[13]), .ZN(n3313) );
  NAND2_X1 U8576 ( .A1(initPC[13]), .A2(n4892), .ZN(n3312) );
  OR2_X1 U8577 ( .A1(n4878), .A2(initPC[14]), .ZN(n3311) );
  NAND2_X1 U8578 ( .A1(initPC[14]), .A2(n4892), .ZN(n3310) );
  OR2_X1 U8579 ( .A1(n4878), .A2(initPC[31]), .ZN(n3309) );
  NAND2_X1 U8580 ( .A1(initPC[31]), .A2(n4892), .ZN(n3308) );
  OAI222_X1 U8581 ( .A1(n8758), .A2(n4831), .B1(n9004), .B2(n4833), .C1(n4635), 
        .C2(n4834), .ZN(memWrData[9]) );
  OAI222_X1 U8582 ( .A1(n8658), .A2(n4831), .B1(n9002), .B2(n4833), .C1(n4636), 
        .C2(n4835), .ZN(memWrData[8]) );
  OAI222_X1 U8583 ( .A1(n8802), .A2(n4831), .B1(n9000), .B2(n4833), .C1(n4638), 
        .C2(n4834), .ZN(memWrData[7]) );
  OAI222_X1 U8584 ( .A1(n8666), .A2(n4831), .B1(n8998), .B2(n4833), .C1(n4639), 
        .C2(n4835), .ZN(memWrData[6]) );
  OAI222_X1 U8585 ( .A1(n8720), .A2(n4831), .B1(n8996), .B2(n4833), .C1(n4640), 
        .C2(n4834), .ZN(memWrData[5]) );
  OAI222_X1 U8586 ( .A1(n8757), .A2(n4831), .B1(n8995), .B2(n4833), .C1(n4641), 
        .C2(n4835), .ZN(memWrData[4]) );
  OAI222_X1 U8587 ( .A1(n8668), .A2(n4831), .B1(n8993), .B2(n4833), .C1(n4642), 
        .C2(n4834), .ZN(memWrData[3]) );
  OAI222_X1 U8588 ( .A1(n8811), .A2(n4831), .B1(n8988), .B2(n4833), .C1(n4702), 
        .C2(n4835), .ZN(memWrData[31]) );
  OAI222_X1 U8589 ( .A1(n8810), .A2(n4831), .B1(n9049), .B2(n4833), .C1(n4363), 
        .C2(n4834), .ZN(memWrData[30]) );
  OAI222_X1 U8590 ( .A1(n8721), .A2(n4831), .B1(n8991), .B2(n4833), .C1(n4643), 
        .C2(n4835), .ZN(memWrData[2]) );
  OAI222_X1 U8591 ( .A1(n8657), .A2(n4830), .B1(n9045), .B2(n4832), .C1(n4364), 
        .C2(n4835), .ZN(memWrData[29]) );
  OAI222_X1 U8592 ( .A1(n8809), .A2(n4830), .B1(n9043), .B2(n4832), .C1(n4365), 
        .C2(n4835), .ZN(memWrData[28]) );
  OAI222_X1 U8593 ( .A1(n8661), .A2(n4830), .B1(n9041), .B2(n4832), .C1(n4366), 
        .C2(n4835), .ZN(memWrData[27]) );
  OAI222_X1 U8594 ( .A1(n8808), .A2(n4830), .B1(n9039), .B2(n4832), .C1(n4367), 
        .C2(n4835), .ZN(memWrData[26]) );
  OAI222_X1 U8595 ( .A1(n8659), .A2(n4830), .B1(n9037), .B2(n4832), .C1(n4703), 
        .C2(n4835), .ZN(memWrData[25]) );
  OAI222_X1 U8596 ( .A1(n8807), .A2(n4830), .B1(n9034), .B2(n4832), .C1(n4674), 
        .C2(n4835), .ZN(memWrData[24]) );
  OAI222_X1 U8597 ( .A1(n8806), .A2(n4830), .B1(n9031), .B2(n4832), .C1(n4717), 
        .C2(n4835), .ZN(memWrData[23]) );
  OAI222_X1 U8598 ( .A1(n8654), .A2(n4830), .B1(n9028), .B2(n4832), .C1(n4718), 
        .C2(n4835), .ZN(memWrData[22]) );
  OAI222_X1 U8599 ( .A1(n8653), .A2(n4830), .B1(n9026), .B2(n4832), .C1(n4719), 
        .C2(n4835), .ZN(memWrData[21]) );
  OAI222_X1 U8600 ( .A1(n8649), .A2(n4830), .B1(n9024), .B2(n4832), .C1(n4720), 
        .C2(n4835), .ZN(memWrData[20]) );
  OAI222_X1 U8601 ( .A1(n8801), .A2(n4830), .B1(n8989), .B2(n4832), .C1(n4644), 
        .C2(n4835), .ZN(memWrData[1]) );
  OAI222_X1 U8602 ( .A1(n8662), .A2(n4831), .B1(n9022), .B2(n4833), .C1(n4721), 
        .C2(n4834), .ZN(memWrData[19]) );
  OAI222_X1 U8603 ( .A1(n8660), .A2(n4830), .B1(n9020), .B2(n4832), .C1(n4722), 
        .C2(n4834), .ZN(memWrData[18]) );
  OAI222_X1 U8604 ( .A1(n8655), .A2(n4831), .B1(n9018), .B2(n4833), .C1(n4723), 
        .C2(n4834), .ZN(memWrData[17]) );
  OAI222_X1 U8605 ( .A1(n8805), .A2(n4830), .B1(n9016), .B2(n4832), .C1(n4724), 
        .C2(n4834), .ZN(memWrData[16]) );
  OAI222_X1 U8606 ( .A1(n8647), .A2(n4831), .B1(n9013), .B2(n4833), .C1(n4637), 
        .C2(n4834), .ZN(memWrData[15]) );
  OAI222_X1 U8607 ( .A1(n8667), .A2(n4830), .B1(n9011), .B2(n4832), .C1(n4645), 
        .C2(n4834), .ZN(memWrData[14]) );
  OAI222_X1 U8608 ( .A1(n8804), .A2(n4831), .B1(n9009), .B2(n4833), .C1(n4646), 
        .C2(n4834), .ZN(memWrData[13]) );
  OAI222_X1 U8609 ( .A1(n8656), .A2(n4830), .B1(n9008), .B2(n4832), .C1(n4647), 
        .C2(n4834), .ZN(memWrData[12]) );
  OAI222_X1 U8610 ( .A1(n8803), .A2(n4831), .B1(n9007), .B2(n4833), .C1(n4648), 
        .C2(n4834), .ZN(memWrData[11]) );
  OAI222_X1 U8611 ( .A1(n8648), .A2(n4830), .B1(n9006), .B2(n4832), .C1(n4649), 
        .C2(n4834), .ZN(memWrData[10]) );
  OAI222_X1 U8612 ( .A1(n8762), .A2(n4831), .B1(n9055), .B2(n4833), .C1(n4632), 
        .C2(n4834), .ZN(memWrData[0]) );
  XNOR2_X1 U8613 ( .A(n8175), .B(n8176), .ZN(n8174) );
  XNOR2_X1 U8614 ( .A(n8178), .B(n8179), .ZN(n8177) );
  XNOR2_X1 U8615 ( .A(n8181), .B(n8182), .ZN(n8180) );
  XNOR2_X1 U8616 ( .A(n8184), .B(n8185), .ZN(n8183) );
  XNOR2_X1 U8617 ( .A(n8187), .B(n8188), .ZN(n8186) );
  XNOR2_X1 U8618 ( .A(n8190), .B(n8191), .ZN(n8189) );
  XNOR2_X1 U8619 ( .A(n8193), .B(n8194), .ZN(n8192) );
  XOR2_X1 U8620 ( .A(n8196), .B(n8197), .Z(n8195) );
  XNOR2_X1 U8621 ( .A(n8851), .B(n8850), .ZN(n8197) );
  OAI22_X1 U8622 ( .A1(n8852), .A2(n8853), .B1(n8198), .B2(n8199), .ZN(n8196)
         );
  INV_X1 U8623 ( .A(n8200), .ZN(n8198) );
  XOR2_X1 U8624 ( .A(n8200), .B(n8199), .Z(n8201) );
  XOR2_X1 U8625 ( .A(n8853), .B(n4526), .Z(n8199) );
  OAI22_X1 U8626 ( .A1(n8854), .A2(n8855), .B1(n8202), .B2(n8203), .ZN(n8200)
         );
  XNOR2_X1 U8627 ( .A(n8205), .B(n8206), .ZN(n8204) );
  XNOR2_X1 U8628 ( .A(n4408), .B(n4109), .ZN(n8206) );
  XNOR2_X1 U8629 ( .A(n8202), .B(n8203), .ZN(n8207) );
  XOR2_X1 U8630 ( .A(n8855), .B(n4534), .Z(n8203) );
  AOI22_X1 U8631 ( .A1(n4540), .A2(n4326), .B1(n8208), .B2(n8209), .ZN(n8202)
         );
  XNOR2_X1 U8632 ( .A(n8208), .B(n8209), .ZN(n8210) );
  XOR2_X1 U8633 ( .A(n4540), .B(n4326), .Z(n8209) );
  OAI22_X1 U8634 ( .A1(n8857), .A2(n8858), .B1(n8211), .B2(n8212), .ZN(n8208)
         );
  XNOR2_X1 U8635 ( .A(n8211), .B(n8212), .ZN(n8213) );
  XOR2_X1 U8636 ( .A(n8858), .B(n4535), .Z(n8212) );
  AOI22_X1 U8637 ( .A1(n4541), .A2(n4327), .B1(n8214), .B2(n8215), .ZN(n8211)
         );
  XNOR2_X1 U8638 ( .A(n8214), .B(n8215), .ZN(n8216) );
  XOR2_X1 U8639 ( .A(n4541), .B(n4327), .Z(n8215) );
  OAI22_X1 U8640 ( .A1(n8860), .A2(n8861), .B1(n8217), .B2(n8218), .ZN(n8214)
         );
  XNOR2_X1 U8641 ( .A(n8217), .B(n8218), .ZN(n8219) );
  XOR2_X1 U8642 ( .A(n8861), .B(n4536), .Z(n8218) );
  AOI22_X1 U8643 ( .A1(n4325), .A2(n4542), .B1(n8220), .B2(n8221), .ZN(n8217)
         );
  XNOR2_X1 U8644 ( .A(n8220), .B(n8221), .ZN(n8222) );
  XOR2_X1 U8645 ( .A(n4542), .B(n4325), .Z(n8221) );
  OAI22_X1 U8646 ( .A1(n8864), .A2(n8865), .B1(n8223), .B2(n8224), .ZN(n8220)
         );
  XNOR2_X1 U8647 ( .A(n8223), .B(n8224), .ZN(n8225) );
  XOR2_X1 U8648 ( .A(n8865), .B(n4456), .Z(n8224) );
  AOI22_X1 U8649 ( .A1(n4278), .A2(n4464), .B1(n8226), .B2(n8227), .ZN(n8223)
         );
  XNOR2_X1 U8650 ( .A(n8226), .B(n8227), .ZN(n8228) );
  XOR2_X1 U8651 ( .A(n4464), .B(n4278), .Z(n8227) );
  OAI22_X1 U8652 ( .A1(n8868), .A2(n8869), .B1(n8229), .B2(n8230), .ZN(n8226)
         );
  XNOR2_X1 U8653 ( .A(n8229), .B(n8230), .ZN(n8231) );
  XOR2_X1 U8654 ( .A(n8869), .B(n4457), .Z(n8230) );
  AOI22_X1 U8655 ( .A1(n4462), .A2(n4279), .B1(n8232), .B2(n8233), .ZN(n8229)
         );
  XNOR2_X1 U8656 ( .A(n8232), .B(n8233), .ZN(n8234) );
  XOR2_X1 U8657 ( .A(n4462), .B(n4279), .Z(n8233) );
  OAI22_X1 U8658 ( .A1(n8872), .A2(n8873), .B1(n8235), .B2(n8236), .ZN(n8232)
         );
  XNOR2_X1 U8659 ( .A(n8235), .B(n8236), .ZN(n8237) );
  XOR2_X1 U8660 ( .A(n8873), .B(n4458), .Z(n8236) );
  AOI22_X1 U8661 ( .A1(n4463), .A2(n4280), .B1(n8238), .B2(n8239), .ZN(n8235)
         );
  XNOR2_X1 U8662 ( .A(n8238), .B(n8239), .ZN(n8240) );
  XOR2_X1 U8663 ( .A(n4463), .B(n4280), .Z(n8239) );
  OAI22_X1 U8664 ( .A1(n8875), .A2(n8876), .B1(n8241), .B2(n8242), .ZN(n8238)
         );
  INV_X1 U8665 ( .A(n8243), .ZN(n8241) );
  XOR2_X1 U8666 ( .A(n8243), .B(n8242), .Z(n8244) );
  XOR2_X1 U8667 ( .A(n8876), .B(n4459), .Z(n8242) );
  OAI22_X1 U8668 ( .A1(n8975), .A2(n8877), .B1(n8245), .B2(n8246), .ZN(n8243)
         );
  XNOR2_X1 U8669 ( .A(n8245), .B(n8246), .ZN(n8247) );
  XOR2_X1 U8670 ( .A(n8975), .B(n4453), .Z(n8246) );
  AOI22_X1 U8671 ( .A1(n4276), .A2(n4465), .B1(n8248), .B2(n8249), .ZN(n8245)
         );
  XNOR2_X1 U8672 ( .A(n8248), .B(n8249), .ZN(n8250) );
  XOR2_X1 U8673 ( .A(n4465), .B(n4276), .Z(n8249) );
  OAI22_X1 U8674 ( .A1(n8881), .A2(n8880), .B1(n8251), .B2(n8252), .ZN(n8248)
         );
  XNOR2_X1 U8675 ( .A(n8251), .B(n8252), .ZN(n8253) );
  XOR2_X1 U8676 ( .A(n8880), .B(n4454), .Z(n8252) );
  AOI22_X1 U8677 ( .A1(n4277), .A2(n4466), .B1(n8254), .B2(n8255), .ZN(n8251)
         );
  XNOR2_X1 U8678 ( .A(n8254), .B(n8255), .ZN(n8256) );
  XOR2_X1 U8679 ( .A(n4466), .B(n4277), .Z(n8255) );
  OAI22_X1 U8680 ( .A1(n8885), .A2(n8884), .B1(n8257), .B2(n8258), .ZN(n8254)
         );
  XNOR2_X1 U8681 ( .A(n8257), .B(n8258), .ZN(n8259) );
  XOR2_X1 U8682 ( .A(n8884), .B(n4397), .Z(n8258) );
  AOI22_X1 U8683 ( .A1(n4170), .A2(n4403), .B1(n8260), .B2(n8261), .ZN(n8257)
         );
  XNOR2_X1 U8684 ( .A(n8260), .B(n8261), .ZN(n8262) );
  XOR2_X1 U8685 ( .A(n4403), .B(n4170), .Z(n8261) );
  OAI22_X1 U8686 ( .A1(n8889), .A2(n8888), .B1(n8263), .B2(n8264), .ZN(n8260)
         );
  XNOR2_X1 U8687 ( .A(n8263), .B(n8264), .ZN(n8265) );
  XOR2_X1 U8688 ( .A(n8888), .B(n4398), .Z(n8264) );
  AOI22_X1 U8689 ( .A1(n4171), .A2(n4404), .B1(n8175), .B2(n8176), .ZN(n8263)
         );
  XOR2_X1 U8690 ( .A(n4404), .B(n4171), .Z(n8176) );
  OAI22_X1 U8691 ( .A1(n8961), .A2(n8892), .B1(n8178), .B2(n8179), .ZN(n8175)
         );
  XOR2_X1 U8692 ( .A(n8961), .B(n4399), .Z(n8179) );
  AOI22_X1 U8693 ( .A1(n4172), .A2(n4405), .B1(n8181), .B2(n8182), .ZN(n8178)
         );
  XOR2_X1 U8694 ( .A(n4405), .B(n4172), .Z(n8182) );
  OAI22_X1 U8695 ( .A1(n8963), .A2(n8895), .B1(n8184), .B2(n8185), .ZN(n8181)
         );
  XOR2_X1 U8696 ( .A(n8963), .B(n4400), .Z(n8185) );
  AOI22_X1 U8697 ( .A1(n4173), .A2(n4406), .B1(n8187), .B2(n8188), .ZN(n8184)
         );
  XOR2_X1 U8698 ( .A(n4406), .B(n4173), .Z(n8188) );
  OAI22_X1 U8699 ( .A1(n8965), .A2(n8898), .B1(n8190), .B2(n8191), .ZN(n8187)
         );
  XOR2_X1 U8700 ( .A(n8965), .B(n4401), .Z(n8191) );
  AOI22_X1 U8701 ( .A1(n4402), .A2(n4174), .B1(n8194), .B2(n8193), .ZN(n8190)
         );
  AOI21_X1 U8702 ( .B1(n8205), .B2(n8900), .A(n8266), .ZN(n8193) );
  AOI21_X1 U8703 ( .B1(n8267), .B2(n4109), .A(n4408), .ZN(n8266) );
  INV_X1 U8704 ( .A(n8267), .ZN(n8205) );
  OAI22_X1 U8705 ( .A1(n8812), .A2(n4368), .B1(n7884), .B2(n8268), .ZN(n8267)
         );
  NAND2_X1 U8706 ( .A1(reg31Val_3[0]), .A2(n4137), .ZN(n8268) );
  XNOR2_X1 U8707 ( .A(n8812), .B(n4368), .ZN(n7884) );
  XOR2_X1 U8708 ( .A(n4402), .B(n4174), .Z(n8194) );
  AOI21_X1 U8709 ( .B1(n8269), .B2(n7573), .A(n4135), .ZN(
        hazard_detect_multiplier_fsm_N19) );
  INV_X1 U8710 ( .A(n7649), .ZN(n8269) );
  MUX2_X1 U8711 ( .A(n8270), .B(n4135), .S(n4537), .Z(
        hazard_detect_multiplier_fsm_N18) );
  NOR2_X1 U8712 ( .A1(n4135), .A2(n7649), .ZN(n8270) );
  NAND3_X1 U8713 ( .A1(n7727), .A2(n7806), .A3(n7829), .ZN(n7649) );
  NAND4_X1 U8714 ( .A1(n8271), .A2(n7789), .A3(n8272), .A4(n8273), .ZN(n7829)
         );
  AOI221_X1 U8715 ( .B1(n8274), .B2(op0_1), .C1(n8275), .C2(n7793), .A(n8276), 
        .ZN(n8273) );
  AOI211_X1 U8716 ( .C1(n7851), .C2(n8277), .A(n4538), .B(n8954), .ZN(n8276)
         );
  NAND2_X1 U8717 ( .A1(n8278), .A2(op0_1), .ZN(n8277) );
  INV_X1 U8718 ( .A(n8279), .ZN(n8275) );
  OAI21_X1 U8719 ( .B1(n7792), .B2(n7850), .A(n4321), .ZN(n8279) );
  INV_X1 U8720 ( .A(n7790), .ZN(n8274) );
  NAND3_X1 U8721 ( .A1(n7611), .A2(n8280), .A3(n8281), .ZN(n8272) );
  AOI21_X1 U8722 ( .B1(n7612), .B2(n4318), .A(n8944), .ZN(n8281) );
  INV_X1 U8723 ( .A(n7812), .ZN(n8271) );
  NOR4_X1 U8724 ( .A1(n4524), .A2(n4321), .A3(n7815), .A4(n7611), .ZN(n7812)
         );
  NAND4_X1 U8725 ( .A1(n8282), .A2(n7810), .A3(n8283), .A4(n7789), .ZN(n7806)
         );
  NAND2_X1 U8726 ( .A1(n7855), .A2(n7859), .ZN(n7789) );
  OAI21_X1 U8727 ( .B1(n8284), .B2(n8285), .A(n7793), .ZN(n8283) );
  INV_X1 U8728 ( .A(n7827), .ZN(n7793) );
  MUX2_X1 U8729 ( .A(n7850), .B(n7792), .S(n4524), .Z(n8285) );
  NOR4_X1 U8730 ( .A1(n4318), .A2(n4129), .A3(n7611), .A4(n8956), .ZN(n7792)
         );
  NOR3_X1 U8731 ( .A1(n4318), .A2(n4129), .A3(n4525), .ZN(n7850) );
  NOR4_X1 U8732 ( .A1(n8286), .A2(n7611), .A3(n8955), .A4(n8956), .ZN(n8284)
         );
  NAND2_X1 U8733 ( .A1(n7849), .A2(n7610), .ZN(n8286) );
  NOR2_X1 U8734 ( .A1(n4524), .A2(n7612), .ZN(n7849) );
  INV_X1 U8735 ( .A(n8287), .ZN(n7810) );
  OAI33_X1 U8736 ( .A1(n8288), .A2(n4538), .A3(n7809), .B1(n8289), .B2(n8944), 
        .B3(n7815), .ZN(n8287) );
  NAND2_X1 U8737 ( .A1(n7612), .A2(n7611), .ZN(n8289) );
  NAND2_X1 U8738 ( .A1(n4120), .A2(n4323), .ZN(n8288) );
  MUX2_X1 U8739 ( .A(n7790), .B(n8290), .S(n8954), .Z(n8282) );
  NAND3_X1 U8740 ( .A1(op0_1), .A2(n4538), .A3(n8278), .ZN(n8290) );
  NAND3_X1 U8741 ( .A1(n8291), .A2(n4538), .A3(n7802), .ZN(n7790) );
  INV_X1 U8742 ( .A(n7851), .ZN(n7802) );
  NAND2_X1 U8743 ( .A1(n8292), .A2(n8293), .ZN(n7727) );
  NOR4_X1 U8744 ( .A1(n7799), .A2(n7798), .A3(n7855), .A4(n8294), .ZN(n8293)
         );
  INV_X1 U8745 ( .A(n7749), .ZN(n8294) );
  OAI21_X1 U8746 ( .B1(n7860), .B2(n7856), .A(n8959), .ZN(n7749) );
  OAI21_X1 U8747 ( .B1(n8953), .B2(n4538), .A(n8958), .ZN(n7856) );
  INV_X1 U8748 ( .A(n7738), .ZN(n7860) );
  NAND3_X1 U8749 ( .A1(n8953), .A2(n4538), .A3(n8954), .ZN(n7738) );
  AND2_X1 U8750 ( .A1(n8959), .A2(n7816), .ZN(n7855) );
  INV_X1 U8751 ( .A(n7750), .ZN(n7799) );
  NAND3_X1 U8752 ( .A1(n7859), .A2(n4554), .A3(n7816), .ZN(n7750) );
  NOR3_X1 U8753 ( .A1(n4323), .A2(n4538), .A3(n4120), .ZN(n7816) );
  AOI211_X1 U8754 ( .C1(n7611), .C2(n8280), .A(n7794), .B(n7805), .ZN(n8292)
         );
  NOR3_X1 U8755 ( .A1(n7851), .A2(n8957), .A3(n8291), .ZN(n7805) );
  NAND2_X1 U8756 ( .A1(op0_1), .A2(n4120), .ZN(n8291) );
  NAND2_X1 U8757 ( .A1(n7861), .A2(n4119), .ZN(n7851) );
  INV_X1 U8758 ( .A(n7737), .ZN(n7861) );
  NAND2_X1 U8759 ( .A1(n8959), .A2(n8958), .ZN(n7737) );
  NAND2_X1 U8760 ( .A1(n7815), .A2(n8295), .ZN(n7794) );
  INV_X1 U8761 ( .A(n8296), .ZN(n8295) );
  AOI21_X1 U8762 ( .B1(n4538), .B2(n7744), .A(n7809), .ZN(n8296) );
  INV_X1 U8763 ( .A(n8278), .ZN(n7809) );
  NOR3_X1 U8764 ( .A1(n8959), .A2(n8953), .A3(n4275), .ZN(n8278) );
  NAND2_X1 U8765 ( .A1(n8280), .A2(n4318), .ZN(n7815) );
  NOR3_X1 U8766 ( .A1(n7827), .A2(n8956), .A3(n4129), .ZN(n8280) );
  NAND3_X1 U8767 ( .A1(n8959), .A2(n8297), .A3(n7744), .ZN(n7827) );
  NOR2_X1 U8768 ( .A1(n4120), .A2(op0_1), .ZN(n7744) );
  NAND2_X1 U8769 ( .A1(n8904), .A2(n7852), .ZN(rs2[4]) );
  NAND2_X1 U8770 ( .A1(n8905), .A2(n7852), .ZN(rs2[3]) );
  NAND2_X1 U8771 ( .A1(n8906), .A2(n7852), .ZN(rs2[2]) );
  INV_X1 U8772 ( .A(n7822), .ZN(rs2[1]) );
  NOR2_X1 U8773 ( .A1(n4328), .A2(n7614), .ZN(n7822) );
  INV_X1 U8774 ( .A(n7823), .ZN(rs2[0]) );
  NOR2_X1 U8775 ( .A1(n4329), .A2(n7614), .ZN(n7823) );
  INV_X1 U8776 ( .A(n7852), .ZN(n7614) );
  NAND2_X1 U8777 ( .A1(op0_1), .A2(n7798), .ZN(n7852) );
  INV_X1 U8778 ( .A(n7740), .ZN(n7798) );
  NAND2_X1 U8779 ( .A1(n8297), .A2(n4120), .ZN(n7740) );
  AND2_X1 U8780 ( .A1(n8957), .A2(n7859), .ZN(n8297) );
  NOR2_X1 U8781 ( .A1(n4119), .A2(n4275), .ZN(n7859) );
  XOR2_X1 U8782 ( .A(n8300), .B(n8301), .Z(n8299) );
  XOR2_X1 U8783 ( .A(n8302), .B(n8303), .Z(n8301) );
  NAND2_X1 U8784 ( .A1(n4442), .A2(n8305), .ZN(n8302) );
  XOR2_X1 U8785 ( .A(n8307), .B(n8308), .Z(n8298) );
  XOR2_X1 U8786 ( .A(n8309), .B(n8310), .Z(n8308) );
  OAI21_X1 U8787 ( .B1(n8311), .B2(n8312), .A(n8313), .ZN(n8310) );
  XOR2_X1 U8788 ( .A(n8314), .B(n8315), .Z(n8307) );
  AOI221_X1 U8789 ( .B1(n7489), .B2(n7713), .C1(n7554), .C2(n8321), .A(n8322), 
        .ZN(n8320) );
  XNOR2_X1 U8790 ( .A(n8305), .B(n4442), .ZN(n8311) );
  OAI21_X1 U8791 ( .B1(n8327), .B2(n8328), .A(n8306), .ZN(n8319) );
  MUX2_X1 U8792 ( .A(n4077), .B(n4731), .S(n8325), .Z(n8328) );
  AOI221_X1 U8793 ( .B1(n7489), .B2(n7962), .C1(n8331), .C2(n4729), .A(n8332), 
        .ZN(n8330) );
  INV_X1 U8794 ( .A(n8334), .ZN(n8331) );
  OAI21_X1 U8795 ( .B1(n8327), .B2(n8337), .A(n8304), .ZN(n8329) );
  MUX2_X1 U8796 ( .A(n4077), .B(n4731), .S(n8335), .Z(n8337) );
  OR2_X1 U8797 ( .A1(n4728), .A2(n8342), .ZN(n8339) );
  OAI21_X1 U8798 ( .B1(n8327), .B2(n8343), .A(n8316), .ZN(n8338) );
  MUX2_X1 U8799 ( .A(n4731), .B(n4077), .S(n7544), .Z(n8343) );
  AOI221_X1 U8800 ( .B1(n7492), .B2(n7971), .C1(n7491), .C2(n7921), .A(n8347), 
        .ZN(n8346) );
  OAI22_X1 U8801 ( .A1(n7488), .A2(n8340), .B1(n8022), .B2(n8323), .ZN(n8347)
         );
  NAND2_X1 U8802 ( .A1(n4729), .A2(n8350), .ZN(n8345) );
  OAI21_X1 U8803 ( .B1(n8327), .B2(n8351), .A(n7720), .ZN(n8344) );
  MUX2_X1 U8804 ( .A(n4731), .B(n4077), .S(n7535), .Z(n8351) );
  AOI221_X1 U8805 ( .B1(n7489), .B2(n7972), .C1(n7554), .C2(n8354), .A(n8355), 
        .ZN(n8353) );
  OAI22_X1 U8806 ( .A1(n7488), .A2(n8323), .B1(n7917), .B2(n8324), .ZN(n8355)
         );
  OAI21_X1 U8807 ( .B1(n8327), .B2(n8356), .A(n7721), .ZN(n8352) );
  MUX2_X1 U8808 ( .A(n4731), .B(n4077), .S(n7543), .Z(n8356) );
  AOI221_X1 U8809 ( .B1(n7489), .B2(n7670), .C1(n8359), .C2(n4729), .A(n8360), 
        .ZN(n8358) );
  OAI22_X1 U8810 ( .A1(n8361), .A2(n8323), .B1(n7967), .B2(n8324), .ZN(n8360)
         );
  INV_X1 U8811 ( .A(n8363), .ZN(n8359) );
  OAI21_X1 U8812 ( .B1(n8327), .B2(n8365), .A(n7722), .ZN(n8357) );
  MUX2_X1 U8813 ( .A(n4731), .B(n4077), .S(n7517), .Z(n8365) );
  AOI221_X1 U8814 ( .B1(n7489), .B2(n7676), .C1(n7554), .C2(n8368), .A(n8369), 
        .ZN(n8367) );
  OAI22_X1 U8815 ( .A1(n8370), .A2(n8323), .B1(n7976), .B2(n8324), .ZN(n8369)
         );
  OAI21_X1 U8816 ( .B1(n8327), .B2(n8372), .A(n7723), .ZN(n8366) );
  MUX2_X1 U8817 ( .A(n4731), .B(n4077), .S(n7522), .Z(n8372) );
  AOI221_X1 U8818 ( .B1(n7489), .B2(n7888), .C1(n8375), .C2(n7554), .A(n8376), 
        .ZN(n8374) );
  OAI22_X1 U8819 ( .A1(n8377), .A2(n8323), .B1(n7669), .B2(n8324), .ZN(n8376)
         );
  INV_X1 U8820 ( .A(n8383), .ZN(n8375) );
  OAI21_X1 U8821 ( .B1(n8327), .B2(n8384), .A(n8326), .ZN(n8373) );
  MUX2_X1 U8822 ( .A(n4731), .B(n4077), .S(n7510), .Z(n8384) );
  AOI221_X1 U8823 ( .B1(n7489), .B2(n7706), .C1(n8387), .C2(n7554), .A(n8388), 
        .ZN(n8386) );
  OAI22_X1 U8824 ( .A1(n7912), .A2(n8323), .B1(n8389), .B2(n8324), .ZN(n8388)
         );
  OAI21_X1 U8825 ( .B1(n8380), .B2(n8394), .A(n8382), .ZN(n8341) );
  INV_X1 U8826 ( .A(n8395), .ZN(n8387) );
  OAI21_X1 U8827 ( .B1(n8327), .B2(n8396), .A(n8364), .ZN(n8385) );
  MUX2_X1 U8828 ( .A(n4731), .B(n4077), .S(n7511), .Z(n8396) );
  AOI221_X1 U8829 ( .B1(n7492), .B2(n7686), .C1(n7491), .C2(n7709), .A(n8400), 
        .ZN(n8399) );
  OAI22_X1 U8830 ( .A1(n7526), .A2(n8340), .B1(n8401), .B2(n8323), .ZN(n8400)
         );
  OAI21_X1 U8831 ( .B1(n8380), .B2(n8403), .A(n8382), .ZN(n8402) );
  OAI22_X1 U8832 ( .A1(n7563), .A2(n8406), .B1(n8407), .B2(n8408), .ZN(n8405)
         );
  NAND2_X1 U8833 ( .A1(n4729), .A2(n8410), .ZN(n8398) );
  OAI21_X1 U8834 ( .B1(n8327), .B2(n8411), .A(n8336), .ZN(n8397) );
  MUX2_X1 U8835 ( .A(n4731), .B(n4077), .S(n7534), .Z(n8411) );
  AOI221_X1 U8836 ( .B1(n7489), .B2(n7685), .C1(n8414), .C2(n7554), .A(n8415), 
        .ZN(n8413) );
  OAI22_X1 U8837 ( .A1(n7526), .A2(n8323), .B1(n7705), .B2(n8324), .ZN(n8415)
         );
  OAI21_X1 U8838 ( .B1(n8380), .B2(n8419), .A(n8382), .ZN(n8393) );
  INV_X1 U8839 ( .A(n8421), .ZN(n8414) );
  OAI21_X1 U8840 ( .B1(n8327), .B2(n8422), .A(n8348), .ZN(n8412) );
  MUX2_X1 U8841 ( .A(n4731), .B(n4077), .S(n7542), .Z(n8422) );
  AOI221_X1 U8842 ( .B1(n7492), .B2(n7695), .C1(n7491), .C2(n7687), .A(n8426), 
        .ZN(n8425) );
  OAI22_X1 U8843 ( .A1(n7505), .A2(n8340), .B1(n8427), .B2(n8323), .ZN(n8426)
         );
  OAI21_X1 U8844 ( .B1(n8380), .B2(n8429), .A(n8382), .ZN(n8362) );
  NAND2_X1 U8845 ( .A1(n4729), .A2(n8434), .ZN(n8424) );
  OAI21_X1 U8846 ( .B1(n8327), .B2(n8435), .A(n8349), .ZN(n8423) );
  MUX2_X1 U8847 ( .A(n4731), .B(n4077), .S(n7533), .Z(n8435) );
  AOI221_X1 U8848 ( .B1(n7489), .B2(n7700), .C1(n8438), .C2(n4729), .A(n8439), 
        .ZN(n8437) );
  OAI22_X1 U8849 ( .A1(n7505), .A2(n8323), .B1(n8433), .B2(n8324), .ZN(n8439)
         );
  AOI22_X1 U8850 ( .A1(n8391), .A2(n8442), .B1(n7560), .B2(n8394), .ZN(n8441)
         );
  OAI21_X1 U8851 ( .B1(n8380), .B2(n8445), .A(n8382), .ZN(n8371) );
  INV_X1 U8852 ( .A(n8446), .ZN(n8438) );
  OAI21_X1 U8853 ( .B1(n8380), .B2(n7561), .A(n8382), .ZN(n8379) );
  OAI21_X1 U8854 ( .B1(n8327), .B2(n8449), .A(n8448), .ZN(n8436) );
  MUX2_X1 U8855 ( .A(n4731), .B(n4077), .S(n7519), .Z(n8449) );
  AOI222_X1 U8856 ( .A1(n7554), .A2(n8456), .B1(n7491), .B2(n7898), .C1(n7490), 
        .C2(n7900), .ZN(n8455) );
  AOI22_X1 U8857 ( .A1(n8457), .A2(n8458), .B1(n8459), .B2(n8460), .ZN(n8454)
         );
  NAND2_X1 U8858 ( .A1(n8461), .A2(n8450), .ZN(n8459) );
  MUX2_X1 U8859 ( .A(n4805), .B(n7674), .S(n8458), .Z(n8461) );
  OAI21_X1 U8860 ( .B1(n7894), .B2(n8460), .A(n7896), .ZN(n8457) );
  OAI21_X1 U8861 ( .B1(n7492), .B2(n7489), .A(n8462), .ZN(n8453) );
  NAND4_X1 U8862 ( .A1(n8465), .A2(n8466), .A3(n8467), .A4(n8468), .ZN(
        aluRes_2[15]) );
  AOI222_X1 U8863 ( .A1(n4729), .A2(n8469), .B1(n7492), .B2(n7900), .C1(n7489), 
        .C2(n7898), .ZN(n8468) );
  AOI22_X1 U8864 ( .A1(n8391), .A2(n8472), .B1(n7560), .B2(n8473), .ZN(n8471)
         );
  NOR2_X1 U8865 ( .A1(n8474), .A2(n7525), .ZN(n8392) );
  AOI221_X1 U8866 ( .B1(n8445), .B2(n8391), .C1(n8390), .C2(n7558), .A(n7564), 
        .ZN(n8416) );
  OAI221_X1 U8867 ( .B1(n8418), .B2(n8476), .C1(n8420), .C2(n7563), .A(n8474), 
        .ZN(n8443) );
  AOI221_X1 U8868 ( .B1(n8394), .B2(n8391), .C1(n8442), .C2(n7558), .A(n7564), 
        .ZN(n8444) );
  AOI22_X1 U8869 ( .A1(n8478), .A2(n8479), .B1(n8480), .B2(n7726), .ZN(n8467)
         );
  NAND2_X1 U8870 ( .A1(n8481), .A2(n8450), .ZN(n8480) );
  NOR2_X1 U8871 ( .A1(n4130), .A2(n4082), .ZN(n8450) );
  MUX2_X1 U8872 ( .A(n4805), .B(n7674), .S(n8479), .Z(n8481) );
  OAI21_X1 U8873 ( .B1(n7726), .B2(n7894), .A(n7896), .ZN(n8478) );
  OAI21_X1 U8874 ( .B1(n7491), .B2(n7490), .A(n8462), .ZN(n8466) );
  OAI221_X1 U8875 ( .B1(n8378), .B2(n8476), .C1(n8447), .C2(n7563), .A(n8474), 
        .ZN(n8404) );
  OAI221_X1 U8876 ( .B1(n8408), .B2(n7563), .C1(n8406), .C2(n8476), .A(n8474), 
        .ZN(n8430) );
  AOI221_X1 U8877 ( .B1(n8432), .B2(n7558), .C1(n8403), .C2(n8391), .A(n7564), 
        .ZN(n8428) );
  NAND2_X1 U8878 ( .A1(n7546), .A2(n7918), .ZN(n8474) );
  NAND2_X1 U8879 ( .A1(n8483), .A2(n4794), .ZN(n8465) );
  XOR2_X1 U8880 ( .A(n8463), .B(n8464), .Z(n8483) );
  NAND2_X1 U8881 ( .A1(n9047), .A2(n4545), .ZN(n8477) );
  OR2_X1 U8882 ( .A1(n7558), .A2(n8380), .ZN(n8382) );
  NOR3_X1 U8883 ( .A1(n4545), .A2(n4136), .A3(n4133), .ZN(n8475) );
  AOI221_X1 U8884 ( .B1(n7560), .B2(n8432), .C1(n8431), .C2(n8019), .A(n8488), 
        .ZN(n8487) );
  OAI221_X1 U8885 ( .B1(n7553), .B2(n8489), .C1(n7497), .C2(n8490), .A(n8491), 
        .ZN(n8431) );
  AOI21_X1 U8886 ( .B1(n7918), .B2(n8403), .A(n7532), .ZN(n8491) );
  OAI221_X1 U8887 ( .B1(n7504), .B2(n8492), .C1(n7516), .C2(n8493), .A(n8494), 
        .ZN(n8403) );
  OAI221_X1 U8888 ( .B1(n7498), .B2(n8492), .C1(n5700), .C2(n8493), .A(n8494), 
        .ZN(n8432) );
  AOI211_X1 U8889 ( .C1(n7559), .C2(n8304), .A(n8496), .B(n8497), .ZN(n8495)
         );
  OAI22_X1 U8890 ( .A1(n7520), .A2(n8485), .B1(n8406), .B2(n8407), .ZN(n8497)
         );
  AOI221_X1 U8891 ( .B1(n8448), .B2(n7530), .C1(n7634), .C2(n7531), .A(n7532), 
        .ZN(n8406) );
  OAI221_X1 U8892 ( .B1(n8408), .B2(n8498), .C1(n7525), .C2(n8409), .A(n8499), 
        .ZN(n8496) );
  AOI221_X1 U8893 ( .B1(n7648), .B2(n7523), .C1(n8336), .C2(n4468), .A(n7532), 
        .ZN(n8409) );
  AOI221_X1 U8894 ( .B1(n7721), .B2(n7530), .C1(n7659), .C2(n7531), .A(n7532), 
        .ZN(n8408) );
  AOI221_X1 U8895 ( .B1(n7560), .B2(n8452), .C1(n8451), .C2(n8019), .A(n8488), 
        .ZN(n8500) );
  OAI221_X1 U8896 ( .B1(n7551), .B2(n8489), .C1(n7496), .C2(n8490), .A(n8501), 
        .ZN(n8451) );
  AOI21_X1 U8897 ( .B1(n7918), .B2(n8381), .A(n7532), .ZN(n8501) );
  INV_X1 U8898 ( .A(n4468), .ZN(n8490) );
  AOI221_X1 U8899 ( .B1(n8460), .B2(n7530), .C1(n7726), .C2(n7531), .A(n7532), 
        .ZN(n8378) );
  AOI221_X1 U8900 ( .B1(n7723), .B2(n7530), .C1(n7617), .C2(n7531), .A(n7532), 
        .ZN(n8447) );
  OAI221_X1 U8901 ( .B1(n8418), .B2(n8407), .C1(n8417), .C2(n7525), .A(n8504), 
        .ZN(n8503) );
  AOI221_X1 U8902 ( .B1(n7559), .B2(n8316), .C1(n8502), .C2(n7663), .A(n8488), 
        .ZN(n8504) );
  AOI221_X1 U8903 ( .B1(n7623), .B2(n7523), .C1(n8348), .C2(n4468), .A(n8505), 
        .ZN(n8417) );
  OAI21_X1 U8904 ( .B1(n7524), .B2(n8420), .A(n8494), .ZN(n8505) );
  AOI221_X1 U8905 ( .B1(n7720), .B2(n7530), .C1(n7661), .C2(n7531), .A(n7532), 
        .ZN(n8420) );
  AOI221_X1 U8906 ( .B1(n8349), .B2(n7530), .C1(n7628), .C2(n7531), .A(n7532), 
        .ZN(n8418) );
  AOI222_X1 U8907 ( .A1(n7559), .A2(n7723), .B1(n7560), .B2(n8472), .C1(n8502), 
        .C2(n7617), .ZN(n8507) );
  AOI21_X1 U8908 ( .B1(n8508), .B2(n8473), .A(n8488), .ZN(n8506) );
  AOI221_X1 U8909 ( .B1(n7726), .B2(n7523), .C1(n8460), .C2(n4468), .A(n7532), 
        .ZN(n8470) );
  OAI221_X1 U8910 ( .B1(n7501), .B2(n8492), .C1(n7513), .C2(n8493), .A(n8494), 
        .ZN(n8445) );
  OAI221_X1 U8911 ( .B1(n7496), .B2(n8492), .C1(n7551), .C2(n8493), .A(n8494), 
        .ZN(n8390) );
  AOI222_X1 U8912 ( .A1(n7559), .A2(n7721), .B1(n7560), .B2(n8442), .C1(n8502), 
        .C2(n7659), .ZN(n8510) );
  NOR2_X1 U8913 ( .A1(n8476), .A2(n8492), .ZN(n8502) );
  OAI221_X1 U8914 ( .B1(n7499), .B2(n8492), .C1(n7549), .C2(n8493), .A(n8494), 
        .ZN(n8442) );
  NAND2_X1 U8915 ( .A1(n7525), .A2(n7918), .ZN(n8407) );
  NAND2_X1 U8916 ( .A1(n7558), .A2(n7531), .ZN(n8486) );
  AOI21_X1 U8917 ( .B1(n8508), .B2(n8394), .A(n8488), .ZN(n8509) );
  INV_X1 U8918 ( .A(n8499), .ZN(n8488) );
  NAND2_X1 U8919 ( .A1(n7532), .A2(n7558), .ZN(n8499) );
  NAND2_X1 U8920 ( .A1(n7525), .A2(n7524), .ZN(n8476) );
  OAI221_X1 U8921 ( .B1(n7503), .B2(n8492), .C1(n7520), .C2(n8493), .A(n8494), 
        .ZN(n8394) );
  INV_X1 U8922 ( .A(n8498), .ZN(n8508) );
  NAND2_X1 U8923 ( .A1(n7918), .A2(n8019), .ZN(n8498) );
  AOI221_X1 U8924 ( .B1(n7634), .B2(n7523), .C1(n8448), .C2(n4468), .A(n7532), 
        .ZN(n8440) );
  NAND4_X1 U8925 ( .A1(n7519), .A2(n7518), .A3(n7521), .A4(n7509), .ZN(n8511)
         );
  NAND4_X1 U8926 ( .A1(n7517), .A2(n7522), .A3(n7510), .A4(n7511), .ZN(n8512)
         );
  NOR3_X1 U8927 ( .A1(n9051), .A2(n9047), .A3(n4121), .ZN(n8482) );
  XOR2_X1 U8928 ( .A(n8514), .B(setInv_2), .Z(n8513) );
  OR2_X1 U8929 ( .A1(n8515), .A2(n8516), .ZN(n8514) );
  NAND4_X1 U8930 ( .A1(n8517), .A2(n9051), .A3(n4545), .A4(n4133), .ZN(n8484)
         );
  MUX2_X1 U8931 ( .A(n8518), .B(n8519), .S(setInv_2), .Z(n8517) );
  OAI21_X1 U8932 ( .B1(n8515), .B2(n4121), .A(n8520), .ZN(n8519) );
  INV_X1 U8933 ( .A(n8521), .ZN(n8518) );
  AOI22_X1 U8934 ( .A1(n8515), .A2(n8522), .B1(n4121), .B2(n8520), .ZN(n8521)
         );
  NOR2_X1 U8935 ( .A1(n8524), .A2(n7509), .ZN(n8516) );
  INV_X1 U8936 ( .A(n8523), .ZN(n8522) );
  NAND4_X1 U8937 ( .A1(n8525), .A2(n8526), .A3(n8527), .A4(n8528), .ZN(n8523)
         );
  NOR4_X1 U8938 ( .A1(n8529), .A2(n8530), .A3(n8531), .A4(n8532), .ZN(n8528)
         );
  NAND4_X1 U8939 ( .A1(n8342), .A2(n7662), .A3(n4469), .A4(n7664), .ZN(n8532)
         );
  XOR2_X1 U8940 ( .A(n8537), .B(n8538), .Z(n8018) );
  XNOR2_X1 U8941 ( .A(n8539), .B(n8540), .ZN(n8342) );
  NAND4_X1 U8942 ( .A1(n7660), .A2(n7656), .A3(n7914), .A4(n7712), .ZN(n8531)
         );
  OAI21_X1 U8943 ( .B1(n8541), .B2(n8542), .A(n8543), .ZN(n7712) );
  OAI21_X1 U8944 ( .B1(n7484), .B2(n8544), .A(n8545), .ZN(n7914) );
  OAI21_X1 U8945 ( .B1(n8546), .B2(n8547), .A(n8548), .ZN(n7656) );
  OAI21_X1 U8946 ( .B1(n8549), .B2(n7555), .A(n8550), .ZN(n7660) );
  NAND4_X1 U8947 ( .A1(n7638), .A2(n7911), .A3(n8334), .A4(n8363), .ZN(n8530)
         );
  OAI21_X1 U8948 ( .B1(n8551), .B2(n8552), .A(n8553), .ZN(n8363) );
  OAI21_X1 U8949 ( .B1(n8554), .B2(n8555), .A(n8556), .ZN(n8334) );
  OAI21_X1 U8950 ( .B1(n8557), .B2(n8558), .A(n8559), .ZN(n7911) );
  OAI21_X1 U8951 ( .B1(n8560), .B2(n8561), .A(n8562), .ZN(n7638) );
  NAND4_X1 U8952 ( .A1(n8383), .A2(n8395), .A3(n8421), .A4(n8446), .ZN(n8529)
         );
  OAI21_X1 U8953 ( .B1(n8563), .B2(n8564), .A(n8565), .ZN(n8446) );
  OAI21_X1 U8954 ( .B1(n8566), .B2(n8567), .A(n8568), .ZN(n8421) );
  OAI21_X1 U8955 ( .B1(n8569), .B2(n8570), .A(n8571), .ZN(n8395) );
  OAI21_X1 U8956 ( .B1(n8572), .B2(n8573), .A(n8574), .ZN(n8383) );
  NOR4_X1 U8957 ( .A1(n8575), .A2(n8469), .A3(n8456), .A4(n8434), .ZN(n8527)
         );
  XOR2_X1 U8958 ( .A(n8576), .B(n8577), .Z(n8434) );
  XOR2_X1 U8959 ( .A(n8578), .B(n8579), .Z(n8456) );
  XOR2_X1 U8960 ( .A(n8580), .B(n8581), .Z(n8469) );
  OR4_X1 U8961 ( .A1(n8368), .A2(n8410), .A3(n8350), .A4(n8354), .ZN(n8575) );
  XNOR2_X1 U8962 ( .A(n8582), .B(n8583), .ZN(n8354) );
  XOR2_X1 U8963 ( .A(n8584), .B(n8585), .Z(n8350) );
  XNOR2_X1 U8964 ( .A(n8586), .B(n8587), .ZN(n8410) );
  XNOR2_X1 U8965 ( .A(n8588), .B(n8589), .ZN(n8368) );
  NOR4_X1 U8966 ( .A1(n7652), .A2(n7557), .A3(n7901), .A4(n4498), .ZN(n8526)
         );
  XOR2_X1 U8967 ( .A(n8590), .B(n8591), .Z(n7901) );
  XOR2_X1 U8968 ( .A(n8592), .B(n8593), .Z(n7658) );
  XOR2_X1 U8969 ( .A(n8594), .B(n8595), .Z(n7652) );
  NOR4_X1 U8970 ( .A1(n7620), .A2(n7692), .A3(n8321), .A4(n7556), .ZN(n8525)
         );
  XOR2_X1 U8971 ( .A(n8596), .B(n8597), .Z(n7616) );
  XOR2_X1 U8972 ( .A(n8598), .B(n8599), .Z(n8321) );
  INV_X1 U8973 ( .A(n7631), .ZN(n7692) );
  XOR2_X1 U8974 ( .A(n8600), .B(n8601), .Z(n7631) );
  XOR2_X1 U8975 ( .A(n8602), .B(n8603), .Z(n7620) );
  XOR2_X1 U8976 ( .A(n8605), .B(n8606), .Z(n8604) );
  AOI22_X1 U8977 ( .A1(n8599), .A2(n8598), .B1(n8607), .B2(n8306), .ZN(n8606)
         );
  OAI21_X1 U8978 ( .B1(n7503), .B2(n8608), .A(n8556), .ZN(n8598) );
  NAND2_X1 U8979 ( .A1(n8554), .A2(n8555), .ZN(n8556) );
  XOR2_X1 U8980 ( .A(n8609), .B(n8316), .Z(n8540) );
  XOR2_X1 U8981 ( .A(n8610), .B(n7720), .Z(n8585) );
  XOR2_X1 U8982 ( .A(n8611), .B(n7721), .Z(n8583) );
  OAI21_X1 U8983 ( .B1(n7501), .B2(n8613), .A(n8553), .ZN(n8582) );
  NAND2_X1 U8984 ( .A1(n8551), .A2(n8552), .ZN(n8553) );
  XNOR2_X1 U8985 ( .A(n8614), .B(n7500), .ZN(n8589) );
  OAI21_X1 U8986 ( .B1(n7527), .B2(n8616), .A(n8574), .ZN(n8588) );
  NAND2_X1 U8987 ( .A1(n8572), .A2(n8573), .ZN(n8574) );
  OAI21_X1 U8988 ( .B1(n7529), .B2(n8617), .A(n8571), .ZN(n8573) );
  NAND2_X1 U8989 ( .A1(n8569), .A2(n8570), .ZN(n8571) );
  XOR2_X1 U8990 ( .A(n8618), .B(n8336), .Z(n8587) );
  OAI21_X1 U8991 ( .B1(n7498), .B2(n8620), .A(n8568), .ZN(n8586) );
  NAND2_X1 U8992 ( .A1(n8566), .A2(n8567), .ZN(n8568) );
  XOR2_X1 U8993 ( .A(n8621), .B(n8349), .Z(n8577) );
  OAI21_X1 U8994 ( .B1(n7495), .B2(n8623), .A(n8565), .ZN(n8622) );
  NAND2_X1 U8995 ( .A1(n8563), .A2(n8564), .ZN(n8565) );
  XOR2_X1 U8996 ( .A(n8624), .B(n7895), .Z(n8591) );
  OAI22_X1 U8997 ( .A1(n7494), .A2(n8626), .B1(n8578), .B2(n8579), .ZN(n8625)
         );
  XOR2_X1 U8998 ( .A(n8626), .B(n8460), .Z(n8579) );
  INV_X1 U8999 ( .A(n8627), .ZN(n8578) );
  OAI22_X1 U9000 ( .A1(n7485), .A2(n8628), .B1(n8580), .B2(n8581), .ZN(n8627)
         );
  XOR2_X1 U9001 ( .A(n7726), .B(n8628), .Z(n8581) );
  NAND2_X1 U9002 ( .A1(n8560), .A2(n8561), .ZN(n8562) );
  XOR2_X1 U9003 ( .A(n7634), .B(n8631), .Z(n8601) );
  OAI21_X1 U9004 ( .B1(n7553), .B2(n8633), .A(n8559), .ZN(n8600) );
  NAND2_X1 U9005 ( .A1(n8557), .A2(n8558), .ZN(n8559) );
  INV_X1 U9006 ( .A(n8634), .ZN(n8558) );
  AOI22_X1 U9007 ( .A1(n7623), .A2(n8635), .B1(n8602), .B2(n8603), .ZN(n8634)
         );
  XOR2_X1 U9008 ( .A(n7623), .B(n8635), .Z(n8603) );
  XOR2_X1 U9009 ( .A(n8637), .B(n7617), .Z(n8597) );
  OAI21_X1 U9010 ( .B1(n7513), .B2(n8639), .A(n8548), .ZN(n8596) );
  NAND2_X1 U9011 ( .A1(n8546), .A2(n8547), .ZN(n8548) );
  XNOR2_X1 U9012 ( .A(n8640), .B(n7514), .ZN(n8593) );
  OAI21_X1 U9013 ( .B1(n7515), .B2(n8642), .A(n8550), .ZN(n8592) );
  NAND2_X1 U9014 ( .A1(n8549), .A2(n7555), .ZN(n8550) );
  XOR2_X1 U9015 ( .A(n7663), .B(n8644), .Z(n8538) );
  NAND2_X1 U9016 ( .A1(n8533), .A2(n8534), .ZN(n8535) );
  XNOR2_X1 U9017 ( .A(n8645), .B(n7665), .ZN(n8533) );
  XOR2_X1 U9018 ( .A(n8536), .B(n7548), .Z(n8645) );
  XNOR2_X1 U9019 ( .A(n8536), .B(n7525), .ZN(n8644) );
  XNOR2_X1 U9020 ( .A(n7661), .B(n8642), .ZN(n8549) );
  XNOR2_X1 U9021 ( .A(n8605), .B(n7524), .ZN(n8642) );
  XOR2_X1 U9022 ( .A(n8605), .B(n7968), .Z(n8640) );
  XNOR2_X1 U9023 ( .A(n8639), .B(n7657), .ZN(n8546) );
  XOR2_X1 U9024 ( .A(n8605), .B(n7977), .Z(n8639) );
  XNOR2_X1 U9025 ( .A(n8536), .B(n7671), .ZN(n8637) );
  XNOR2_X1 U9026 ( .A(n7648), .B(n8636), .ZN(n8541) );
  XNOR2_X1 U9027 ( .A(n7550), .B(n8605), .ZN(n8636) );
  XOR2_X1 U9028 ( .A(n7682), .B(n8536), .Z(n8635) );
  XNOR2_X1 U9029 ( .A(n7628), .B(n8633), .ZN(n8557) );
  XOR2_X1 U9030 ( .A(n7906), .B(n8605), .Z(n8633) );
  XOR2_X1 U9031 ( .A(n7696), .B(n8605), .Z(n8631) );
  XOR2_X1 U9032 ( .A(n7641), .B(n8629), .Z(n8560) );
  XOR2_X1 U9033 ( .A(n7988), .B(n8536), .Z(n8629) );
  OAI22_X1 U9034 ( .A1(n4837), .A2(n9012), .B1(n4838), .B2(n8833), .ZN(n8646)
         );
  XOR2_X1 U9035 ( .A(n8479), .B(n8605), .Z(n8628) );
  XOR2_X1 U9036 ( .A(n8536), .B(n7521), .Z(n8626) );
  XOR2_X1 U9037 ( .A(n8536), .B(n7518), .Z(n8624) );
  XNOR2_X1 U9038 ( .A(n8623), .B(n8448), .ZN(n8563) );
  XOR2_X1 U9039 ( .A(n8536), .B(n7519), .Z(n8623) );
  XOR2_X1 U9040 ( .A(n8536), .B(n7533), .Z(n8621) );
  XNOR2_X1 U9041 ( .A(n8620), .B(n8348), .ZN(n8566) );
  XOR2_X1 U9042 ( .A(n8536), .B(n7542), .Z(n8620) );
  XOR2_X1 U9043 ( .A(n8536), .B(n7534), .Z(n8618) );
  XNOR2_X1 U9044 ( .A(n8617), .B(n8364), .ZN(n8569) );
  XOR2_X1 U9045 ( .A(n8536), .B(n7511), .Z(n8617) );
  XNOR2_X1 U9046 ( .A(n8616), .B(n8326), .ZN(n8572) );
  XNOR2_X1 U9047 ( .A(n8605), .B(n7510), .ZN(n8616) );
  XNOR2_X1 U9048 ( .A(n8605), .B(n7522), .ZN(n8614) );
  XNOR2_X1 U9049 ( .A(n8613), .B(n7722), .ZN(n8551) );
  XNOR2_X1 U9050 ( .A(n8605), .B(n7517), .ZN(n8613) );
  XNOR2_X1 U9051 ( .A(n8605), .B(n7543), .ZN(n8611) );
  XNOR2_X1 U9052 ( .A(n8536), .B(n7535), .ZN(n8610) );
  XNOR2_X1 U9053 ( .A(n8605), .B(n7544), .ZN(n8609) );
  XOR2_X1 U9054 ( .A(n7503), .B(n8608), .Z(n8554) );
  XNOR2_X1 U9055 ( .A(n8605), .B(n7545), .ZN(n8608) );
  XOR2_X1 U9056 ( .A(n8306), .B(n8607), .Z(n8599) );
  XNOR2_X1 U9057 ( .A(n8605), .B(n8325), .ZN(n8607) );
  AND2_X1 U9058 ( .A1(n9057), .A2(n9058), .ZN(n8173) );
  NOR2_X1 U9059 ( .A1(n4156), .A2(n4373), .ZN(n8116) );
  DFFS_X1 hazard_detect_multiplier_fsm_if_id_mult_ctrl_reg_1_ ( .D(
        hazard_detect_multiplier_fsm_N19), .CK(clk), .SN(n4877), .Q(n4593) );
  DFFS_X1 hazard_detect_multiplier_fsm_id_ex_mult_ctrl_reg_1_ ( .D(
        hazard_detect_multiplier_fsm_N19), .CK(clk), .SN(n4877), .QN(n4898) );
  DFFS_X1 hazard_detect_multiplier_fsm_ex_mem_mult_ctrl_reg_1_ ( .D(
        hazard_detect_multiplier_fsm_N19), .CK(clk), .SN(n4877), .Q(n4569) );
endmodule

