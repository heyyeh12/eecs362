
module pipeline ( clk, rst, initPC, instruction, iAddr, memAddr, memRdData, 
        memWrData, dSize, memWr, busA, busB, busFP, rs1, rs2, rd, regWrData, 
        regWr, fp );
  input [31:0] initPC;
  input [31:0] instruction;
  output [31:0] iAddr;
  output [31:0] memAddr;
  input [31:0] memRdData;
  output [31:0] memWrData;
  output [1:0] dSize;
  input [31:0] busA;
  input [31:0] busB;
  input [31:0] busFP;
  output [4:0] rs1;
  output [4:0] rs2;
  output [4:0] rd;
  output [31:0] regWrData;
  input clk, rst;
  output memWr, regWr, fp;
  wire   n7908, op0_1, valid_2, valid_3, setInv_2, op0_2, zeroExt_2, link_3,
         fp_3, \id_ex/N45 , \id_ex/N42 , \id_ex/N41 , \id_ex/N40 , \id_ex/N38 ,
         \id_ex/N37 , \id_ex/N33 , \id_ex/N31 , \id_ex/N4 , \ex_mem/N247 ,
         \ex_mem/N246 , \ex_mem/N245 , \ex_mem/N244 , \ex_mem/N243 ,
         \ex_mem/N242 , \ex_mem/N241 , \ex_mem/N240 , \ex_mem/N239 ,
         \ex_mem/N237 , \ex_mem/N236 , \ex_mem/N235 , \ex_mem/N234 ,
         \ex_mem/N233 , \ex_mem/N232 , \ex_mem/N231 , \ex_mem/N230 ,
         \ex_mem/N229 , \ex_mem/N227 , \ex_mem/N226 , \ex_mem/N225 ,
         \ex_mem/N224 , \ex_mem/N223 , \ex_mem/N222 , \ex_mem/N221 ,
         \ex_mem/N220 , \ex_mem/N219 , \ex_mem/N218 , \ex_mem/N217 ,
         \ex_mem/N216 , \ex_mem/N215 , \ex_mem/N214 , \ex_mem/N213 ,
         \ex_mem/N212 , \ex_mem/N211 , \ex_mem/N210 , \ex_mem/N209 ,
         \ex_mem/N208 , \ex_mem/N207 , \ex_mem/N206 , \ex_mem/N205 ,
         \ex_mem/N204 , \ex_mem/N203 , \ex_mem/N202 , \ex_mem/N200 ,
         \ex_mem/N199 , \ex_mem/N198 , \ex_mem/N197 , \ex_mem/N196 ,
         \ex_mem/N162 , \ex_mem/N161 , \ex_mem/N160 , \ex_mem/N159 ,
         \ex_mem/N158 , \ex_mem/N157 , \ex_mem/N156 , \ex_mem/N155 ,
         \ex_mem/N154 , \ex_mem/N153 , \ex_mem/N152 , \ex_mem/N151 ,
         \ex_mem/N150 , \ex_mem/N149 , \ex_mem/N148 , \ex_mem/N147 ,
         \ex_mem/N146 , \ex_mem/N145 , \ex_mem/N144 , \ex_mem/N143 ,
         \ex_mem/N142 , \ex_mem/N141 , \ex_mem/N140 , \ex_mem/N139 ,
         \ex_mem/N138 , \ex_mem/N137 , \ex_mem/N136 , \ex_mem/N135 ,
         \ex_mem/N134 , \ex_mem/N133 , \ex_mem/N132 , \ex_mem/N131 ,
         \ex_mem/N130 , \ex_mem/N129 , \ex_mem/N128 , \ex_mem/N127 ,
         \ex_mem/N126 , \ex_mem/N125 , \ex_mem/N124 , \ex_mem/N123 ,
         \ex_mem/N122 , \ex_mem/N121 , \ex_mem/N120 , \ex_mem/N119 ,
         \ex_mem/N118 , \ex_mem/N117 , \ex_mem/N116 , \ex_mem/N115 ,
         \ex_mem/N114 , \ex_mem/N113 , \ex_mem/N112 , \ex_mem/N111 ,
         \ex_mem/N110 , \ex_mem/N109 , \ex_mem/N108 , \ex_mem/N107 ,
         \ex_mem/N106 , \ex_mem/N105 , \ex_mem/N104 , \ex_mem/N103 ,
         \ex_mem/N102 , \ex_mem/N101 , \ex_mem/N100 , \ex_mem/N99 ,
         \ex_mem/N66 , \ex_mem/N65 , \ex_mem/N64 , \ex_mem/N63 , \ex_mem/N62 ,
         \ex_mem/N61 , \ex_mem/N60 , \ex_mem/N59 , \ex_mem/N58 , \ex_mem/N57 ,
         \ex_mem/N56 , \ex_mem/N55 , \ex_mem/N54 , \ex_mem/N53 , \ex_mem/N52 ,
         \ex_mem/N51 , \ex_mem/N50 , \ex_mem/N49 , \ex_mem/N48 , \ex_mem/N47 ,
         \ex_mem/N46 , \ex_mem/N45 , \ex_mem/N44 , \ex_mem/N43 , \ex_mem/N42 ,
         \ex_mem/N41 , \ex_mem/N40 , \ex_mem/N39 , \ex_mem/N38 , \ex_mem/N37 ,
         \ex_mem/N36 , \ex_mem/N35 , \mem_wb/N41 , \mem_wb/N36 ,
         \mem/addImm/mux_map1/M3/z2[31] , n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1950, n1952,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1986, n1990,
         n1992, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2083, n2084, n2086, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2116,
         n2118, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2133, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2220, n2222, n2223, n2224, n2225, n2227, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n8108, n7907, n7906, n2528, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2544, n2545, n2546,
         n2547, n2548, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, net33021, \hazard_detect/eq_83/A[0] ,
         \hazard_detect/eq_83/A[1] , \hazard_detect/eq_83/A[2] ,
         \hazard_detect/eq_83/A[3] , \hazard_detect/eq_83/A[4] , net33193,
         net33197, net33204, net33205, net33207, net33219, net33230, net33276,
         net33280, net36084, net35542, net35483, net35052, net35047, net35037,
         net35036, net34763, net34726, net34717, net34613, net133771,
         net220285, net220292, net220293, net220294, net220295, net220297,
         net220305, net220307, net220310, net220312, net220313, net220315,
         net220319, net220320, net220354, net220403, net220405, net220409,
         net220517, net220535, net220536, net220537, net220539, net220540,
         net220601, net220632, net220637, net220638, net220640, net220644,
         net220646, net220651, net220656, net220663, net220714, net220720,
         net220728, net220729, net220746, net220753, net220757, net220766,
         net220767, net220769, net220775, net220778, net220780, net220838,
         net220849, net220851, net220865, net220874, net220875, net220876,
         net220882, net220885, net220888, net220889, net220890, net220894,
         net220895, net220921, net221152, net221153, net221157, net221163,
         net221165, net221340, net221411, net221416, net221424, net221426,
         net221431, net221442, net221477, net221479, net221481, net221487,
         net221489, net221490, net221491, net221492, net221494, net221531,
         net221648, net221652, net221754, net221757, net221758, net221759,
         net221761, net221762, net221763, net221765, net221766, net221791,
         net221792, net221793, net221798, net221800, net221802, net221806,
         net221807, net221812, net221813, net221818, net221819, net221820,
         net221856, net221858, net221862, net221864, net221874, net221878,
         net221881, net221888, net221905, net221922, net221924, net221929,
         net222151, net222155, net222370, net222371, net222515, net222672,
         net222745, net222840, net223209, net223242, net223245, net223262,
         net223300, net223329, net223337, net223338, net223345, net223346,
         net223348, net223437, net223657, net223721, net223781, net224727,
         net224725, net224723, net224721, net224719, net224717, net224713,
         net224711, net224703, net224699, net224693, net224691, net224685,
         net224683, net224681, net224679, net224675, net224673, net224671,
         net224669, net224663, net224661, net224659, net224657, net224655,
         net224653, net224645, net224643, net224641, net224639, net224637,
         net224635, net224633, net224631, net224629, net224627, net224625,
         net224623, net224621, net224619, net224617, net224615, net224613,
         net224611, net224753, net224751, net224749, net224747, net224745,
         net224743, net224741, net224737, net224735, net224733, net224731,
         net224759, net224755, net224767, net224765, net224777, net224773,
         net224789, net224787, net224785, net224783, net224781, net224835,
         net224833, net224843, net224855, net224853, net224851, net224849,
         net224869, net224865, net224861, net224859, net224871, net224919,
         net224915, net224913, net224909, net224903, net224901, net224899,
         net224897, net224895, net224893, net224891, net224929, net224925,
         net224957, net224955, net224953, net224947, net224943, net224939,
         net224937, net224933, net224967, net224965, net224999, net224997,
         net224995, net224993, net224991, net225003, net225001, net225013,
         net225011, net225017, net225015, net225029, net225051, net225049,
         net225047, net225045, net225053, net225084, net225083, net225082,
         net225091, net225096, net225102, net225101, net225216, net225214,
         net225226, net225230, net225238, net225237, net225243, net225251,
         net225378, net225434, net225520, net225580, net225588, net225587,
         net225601, net225605, net225622, net227791, net227817, net227828,
         net227884, net227945, net227982, net228018, net228029, net228058,
         net228074, net228087, net228081, net228080, net228094, net228093,
         net228150, net228149, net228148, net228159, net228233, net228276,
         net228280, net228287, net228326, net228323, net228341, net228345,
         net228359, net228407, net228479, net228541, net228552, net228597,
         net228610, net228697, net228700, net228710, net228707, net228720,
         net228735, net228809, net228816, net228858, net228869, net228909,
         net228915, net228921, net228936, net228942, net228941, net228949,
         net228982, net228981, net229005, net229037, net229061, net229071,
         net229173, net229239, net229271, net229270, net229307, net229330,
         net229367, net229370, net229393, net229454, net229482, net229481,
         net229522, net229575, net229579, net229596, net229606, net229624,
         net229628, net229646, net229656, net229691, net229719, net229782,
         net229784, net229952, net229958, net229988, net230040, net230088,
         net230097, net230103, net230130, net230145, net230144, net230143,
         net230142, net230157, net230181, net230191, net230199, net230226,
         net230225, net230231, net230245, net230488, net230493, net230611,
         net230622, net230683, net230730, net230733, net230741, net230760,
         net228768, net221817, net221488, net223341, net223340, net225242,
         net223342, net222771, net221875, net229291, net225600, net221892,
         net221890, net221889, net220619, net228677, net220314, net225229,
         net222698, net229486, net224873, net222156, net221473, net220524,
         net228495, net221805, net221799, net221770, net221432, net220322,
         net220318, net220316, net220299, net227823, net225581, net225055,
         net223347, net223339, net222353, net222161, net222158, net220323,
         net228940, net228715, net228056, net220747, net228615, net225095,
         net223343, net229737, net229736, net228708, net221876, net221863,
         net221769, net221425, net220301, net220300, net220298, net220296,
         net220289, net220288, net220287, net220286, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2664, n2665, n2666, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3144, n3146, n3147, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3252, n3253,
         n3254, n3255, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3610, n3611, n3612, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3784, n3785, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3884, n3885, n3887, n3888, n3891, n3892, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5314, n5315, n5316,
         n5317, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n8109, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7857, n7859, n7861, n7862, n7863, n7866, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107;
  wire   [27:0] instr_2;
  wire   [4:0] rd_2;
  wire   [4:0] rd_3;
  wire   [1:0] reg31Val_3;
  wire   [31:0] reg31Val_0;
  wire   [31:0] \wb/dsize_reg/z2 ;
  assign \mem_wb/N41  = rst;
  assign rs2[0] = \hazard_detect/eq_83/A[0] ;
  assign rs2[1] = \hazard_detect/eq_83/A[1] ;
  assign rs2[2] = \hazard_detect/eq_83/A[2] ;
  assign rs2[3] = \hazard_detect/eq_83/A[3] ;
  assign rs2[4] = \hazard_detect/eq_83/A[4] ;
  assign regWr = net230040;
  assign iAddr[27] = n3790;

  DFFR_X1 \ex_mem/aluRes_q_reg[0]  ( .D(net133771), .CK(clk), .RN(net224623), 
        .Q(memAddr[0]), .QN(n7542) );
  DFFR_X1 \ex_mem/aluRes_q_reg[16]  ( .D(\ex_mem/N212 ), .CK(clk), .RN(
        net224623), .Q(memAddr[16]), .QN(n7541) );
  DFFR_X1 \ex_mem/aluRes_q_reg[21]  ( .D(\ex_mem/N217 ), .CK(clk), .RN(
        net224623), .Q(memAddr[21]), .QN(n7540) );
  DFFR_X1 \ex_mem/aluRes_q_reg[22]  ( .D(\ex_mem/N218 ), .CK(clk), .RN(
        net224623), .Q(memAddr[22]), .QN(n7539) );
  DFFR_X1 \ex_mem/aluRes_q_reg[23]  ( .D(\ex_mem/N219 ), .CK(clk), .RN(
        net224623), .Q(memAddr[23]), .QN(n7538) );
  DFFR_X1 \ex_mem/aluRes_q_reg[24]  ( .D(\ex_mem/N220 ), .CK(clk), .RN(
        net224623), .Q(memAddr[24]), .QN(n7537) );
  DFFR_X1 \ex_mem/aluRes_q_reg[25]  ( .D(\ex_mem/N221 ), .CK(clk), .RN(
        net224623), .Q(memAddr[25]), .QN(n7536) );
  DFFR_X1 \ex_mem/aluRes_q_reg[31]  ( .D(\ex_mem/N227 ), .CK(clk), .RN(
        net224623), .Q(memAddr[31]), .QN(n7535) );
  DFFR_X1 \ex_mem/aluRes_q_reg[4]  ( .D(\ex_mem/N199 ), .CK(clk), .RN(
        net224621), .Q(memAddr[4]), .QN(n7534) );
  DFFR_X1 \ex_mem/aluRes_q_reg[9]  ( .D(\ex_mem/N205 ), .CK(clk), .RN(
        net224621), .Q(memAddr[9]), .QN(n7533) );
  DFFR_X1 \ex_mem/aluRes_q_reg[2]  ( .D(\ex_mem/N197 ), .CK(clk), .RN(
        net224621), .Q(memAddr[2]), .QN(n7532) );
  DFFR_X1 \ex_mem/aluRes_q_reg[1]  ( .D(\ex_mem/N196 ), .CK(clk), .RN(
        net224621), .Q(memAddr[1]), .QN(n7531) );
  DFFR_X1 \ex_mem/aluRes_q_reg[6]  ( .D(\ex_mem/N202 ), .CK(clk), .RN(
        net224621), .Q(memAddr[6]), .QN(n7529) );
  DFFR_X1 \ex_mem/aluRes_q_reg[11]  ( .D(\ex_mem/N207 ), .CK(clk), .RN(
        net224621), .Q(memAddr[11]), .QN(n7528) );
  DFFR_X1 \ex_mem/aluRes_q_reg[7]  ( .D(\ex_mem/N203 ), .CK(clk), .RN(
        net224621), .Q(memAddr[7]), .QN(n7527) );
  DFFR_X1 \ex_mem/aluRes_q_reg[29]  ( .D(\ex_mem/N225 ), .CK(clk), .RN(
        net224621), .Q(memAddr[29]), .QN(n7526) );
  DFFR_X1 \ex_mem/aluRes_q_reg[8]  ( .D(\ex_mem/N204 ), .CK(clk), .RN(
        net224621), .Q(memAddr[8]), .QN(n7525) );
  DFFR_X1 \ex_mem/aluRes_q_reg[12]  ( .D(\ex_mem/N208 ), .CK(clk), .RN(
        net224621), .Q(memAddr[12]), .QN(n7524) );
  DFFR_X1 \ex_mem/aluRes_q_reg[13]  ( .D(\ex_mem/N209 ), .CK(clk), .RN(
        net224621), .Q(memAddr[13]), .QN(n7523) );
  DFFR_X1 \ex_mem/aluRes_q_reg[10]  ( .D(\ex_mem/N206 ), .CK(clk), .RN(
        net224619), .Q(memAddr[10]), .QN(n7522) );
  DFFR_X1 \ex_mem/aluRes_q_reg[30]  ( .D(\ex_mem/N226 ), .CK(clk), .RN(
        net224617), .Q(memAddr[30]), .QN(n7500) );
  DFFR_X1 \ex_mem/fp_q_reg  ( .D(n7358), .CK(clk), .RN(net224615), .Q(fp_3) );
  DFFR_X1 \ex_mem/rd_q_reg[1]  ( .D(\ex_mem/N244 ), .CK(clk), .RN(net224615), 
        .Q(rd_3[1]) );
  DFFR_X1 \id_ex/instr_q_reg[5]  ( .D(n7378), .CK(clk), .RN(net224615), .Q(
        instr_2[5]) );
  DFFR_X1 \id_ex/instr_q_reg[3]  ( .D(n7362), .CK(clk), .RN(net224615), .QN(
        n7498) );
  DFFR_X1 \id_ex/instr_q_reg[27]  ( .D(\id_ex/N31 ), .CK(clk), .RN(net224613), 
        .Q(instr_2[27]) );
  DFFR_X1 \id_ex/instr_q_reg[26]  ( .D(n7359), .CK(clk), .RN(net224613), .Q(
        instr_2[26]) );
  DFFR_X1 \id_ex/instr_q_reg[23]  ( .D(n7371), .CK(clk), .RN(net224613), .QN(
        n7489) );
  DFFR_X1 \id_ex/instr_q_reg[22]  ( .D(n7370), .CK(clk), .RN(net224613), .QN(
        n7488) );
  DFFR_X1 \id_ex/instr_q_reg[21]  ( .D(n7369), .CK(clk), .RN(net224613), .QN(
        n7487) );
  DFFR_X1 \id_ex/instr_q_reg[20]  ( .D(n3074), .CK(clk), .RN(net224613), .QN(
        n7486) );
  DFFR_X1 \id_ex/instr_q_reg[19]  ( .D(n3073), .CK(clk), .RN(net224613), .Q(
        instr_2[19]) );
  DFFR_X1 \id_ex/instr_q_reg[18]  ( .D(n3072), .CK(clk), .RN(net224613), .Q(
        instr_2[18]) );
  DFFR_X1 \id_ex/instr_q_reg[17]  ( .D(n3071), .CK(clk), .RN(net224611), .Q(
        instr_2[17]) );
  DFFR_X1 \id_ex/instr_q_reg[16]  ( .D(n2835), .CK(clk), .RN(net224611), .QN(
        n3085) );
  DFFR_X1 \id_ex/instr_q_reg[14]  ( .D(n7375), .CK(clk), .RN(net224611), .QN(
        n7484) );
  DFFR_X1 \id_ex/instr_q_reg[13]  ( .D(n7374), .CK(clk), .RN(net224611), .QN(
        n7483) );
  DFFR_X1 \id_ex/instr_q_reg[12]  ( .D(n7373), .CK(clk), .RN(net224611), .QN(
        n7482) );
  DFFR_X1 \id_ex/instr_q_reg[11]  ( .D(n7368), .CK(clk), .RN(net224611), .QN(
        n7481) );
  DFFR_X1 \id_ex/instr_q_reg[9]  ( .D(n7366), .CK(clk), .RN(net224611), .Q(
        instr_2[9]) );
  DFFR_X1 \id_ex/instr_q_reg[8]  ( .D(n7365), .CK(clk), .RN(net224611), .Q(
        instr_2[8]) );
  DFFR_X1 \id_ex/instr_q_reg[7]  ( .D(n7364), .CK(clk), .RN(net224611), .Q(
        instr_2[7]) );
  DFFR_X1 \id_ex/instr_q_reg[6]  ( .D(n7363), .CK(clk), .RN(net224611), .Q(
        instr_2[6]) );
  DFFR_X1 \id_ex/instr_q_reg[31]  ( .D(n2795), .CK(clk), .RN(net224617), .Q(
        n2922) );
  DFFR_X1 \id_ex/regWr_q_reg  ( .D(\id_ex/N37 ), .CK(clk), .RN(net224633), 
        .QN(n7479) );
  DFFR_X1 \ex_mem/rd_q_reg[4]  ( .D(\ex_mem/N247 ), .CK(clk), .RN(net224655), 
        .Q(rd_3[4]) );
  DFFR_X1 \ex_mem/valid_q_reg  ( .D(\ex_mem/N241 ), .CK(clk), .RN(net224657), 
        .Q(valid_3) );
  DFFR_X1 \ex_mem/link_q_reg  ( .D(\ex_mem/N236 ), .CK(clk), .RN(net224643), 
        .Q(link_3) );
  DFFR_X1 \ex_mem/regWr_q_reg  ( .D(\ex_mem/N231 ), .CK(clk), .RN(net224661), 
        .Q(\mem_wb/N36 ) );
  DFFR_X1 \ex_mem/memWr_q_reg  ( .D(\ex_mem/N230 ), .CK(clk), .RN(net224663), 
        .Q(memWr) );
  DFFR_X1 \id_ex/memWrData_sel_q_reg[1]  ( .D(n7875), .CK(clk), .RN(net224633), 
        .QN(n7470) );
  DFFR_X1 \ex_mem/busA_q_reg[30]  ( .D(n2544), .CK(clk), .RN(net224633), .Q(
        n3111) );
  DFFR_X1 \ex_mem/busA_q_reg[29]  ( .D(n2533), .CK(clk), .RN(net224629), .Q(
        n3112) );
  DFFR_X1 \ex_mem/busA_q_reg[13]  ( .D(n2531), .CK(clk), .RN(net224653), .Q(
        n3103) );
  DFFR_X1 \ex_mem/busA_q_reg[12]  ( .D(n2553), .CK(clk), .RN(net224635), .Q(
        n3104) );
  DFFR_X1 \ex_mem/busA_q_reg[11]  ( .D(n2554), .CK(clk), .RN(net224659), .Q(
        n3115) );
  DFFR_X1 \ex_mem/busA_q_reg[9]  ( .D(n2539), .CK(clk), .RN(net224627), .Q(
        n3102) );
  DFFR_X1 \ex_mem/busA_q_reg[8]  ( .D(n2546), .CK(clk), .RN(net224625), .Q(
        n3100) );
  DFFR_X1 \ex_mem/busA_q_reg[6]  ( .D(n2542), .CK(clk), .RN(net224657), .Q(
        n3101) );
  DFFR_X1 \ex_mem/imm32_q_reg[31]  ( .D(\ex_mem/N162 ), .CK(clk), .RN(
        net224673), .Q(\mem/addImm/mux_map1/M3/z2[31] ) );
  DFFR_X1 \ex_mem/busA_q_reg[2]  ( .D(n2534), .CK(clk), .RN(net224639), .Q(
        n2991) );
  DFFR_X1 \ex_mem/busA_q_reg[3]  ( .D(n2558), .CK(clk), .RN(net224639), .Q(
        n2990) );
  DFFR_X1 \ex_mem/aluRes_q_reg[28]  ( .D(\ex_mem/N224 ), .CK(clk), .RN(
        net224639), .Q(memAddr[28]), .QN(n7424) );
  DFFR_X1 \ex_mem/busA_q_reg[27]  ( .D(n2556), .CK(clk), .RN(net224637), .Q(
        n3113) );
  DFFR_X1 \ex_mem/aluRes_q_reg[26]  ( .D(\ex_mem/N222 ), .CK(clk), .RN(
        net224637), .Q(memAddr[26]), .QN(n7421) );
  DFFR_X1 \ex_mem/busA_q_reg[26]  ( .D(n2535), .CK(clk), .RN(net224637), .Q(
        n3107) );
  DFFR_X1 \ex_mem/aluRes_q_reg[5]  ( .D(\ex_mem/N200 ), .CK(clk), .RN(
        net224637), .Q(memAddr[5]), .QN(n7420) );
  DFFR_X1 \ex_mem/busA_q_reg[5]  ( .D(n2536), .CK(clk), .RN(net224637), .Q(
        n3099) );
  DFFR_X1 \ex_mem/busA_q_reg[25]  ( .D(n2541), .CK(clk), .RN(net224637), .Q(
        n3108) );
  DFFR_X1 \ex_mem/busA_q_reg[24]  ( .D(n2550), .CK(clk), .RN(net224637), .Q(
        n3110) );
  DFFR_X1 \ex_mem/busA_q_reg[23]  ( .D(n2545), .CK(clk), .RN(net224637), .Q(
        n3109) );
  DFFR_X1 \ex_mem/busA_q_reg[22]  ( .D(n2540), .CK(clk), .RN(net224637), .Q(
        n3114) );
  DFFR_X1 \ex_mem/busA_q_reg[16]  ( .D(n2548), .CK(clk), .RN(net224635), .Q(
        n3098) );
  DFFR_X1 \ex_mem/aluRes_q_reg[14]  ( .D(\ex_mem/N210 ), .CK(clk), .RN(
        net224635), .Q(memAddr[14]), .QN(n7417) );
  DFFR_X1 \ex_mem/aluRes_q_reg[20]  ( .D(\ex_mem/N216 ), .CK(clk), .RN(
        net224635), .Q(memAddr[20]), .QN(n7415) );
  DFFR_X1 \ex_mem/busA_q_reg[20]  ( .D(n2555), .CK(clk), .RN(net224635), .Q(
        n2993) );
  DFFR_X1 \ex_mem/aluRes_q_reg[15]  ( .D(\ex_mem/N211 ), .CK(clk), .RN(
        net224635), .Q(memAddr[15]), .QN(n7414) );
  DFFR_X1 \ex_mem/aluRes_q_reg[18]  ( .D(\ex_mem/N214 ), .CK(clk), .RN(
        net224635), .Q(memAddr[18]), .QN(n7412) );
  DFFR_X1 \ex_mem/busA_q_reg[18]  ( .D(n2532), .CK(clk), .RN(net224635), .Q(
        n3116) );
  DFFR_X1 \ex_mem/aluRes_q_reg[17]  ( .D(\ex_mem/N213 ), .CK(clk), .RN(
        net224635), .Q(memAddr[17]), .QN(n7411) );
  DFFR_X1 \ex_mem/busA_q_reg[17]  ( .D(n2537), .CK(clk), .RN(net224635), .Q(
        n3105) );
  DFFR_X1 \ex_mem/busA_q_reg[19]  ( .D(n2552), .CK(clk), .RN(net224633), .Q(
        n3106) );
  DFFR_X1 \if_id/incPC_q_reg[10]  ( .D(n2214), .CK(clk), .RN(net224629), .Q(
        n3031) );
  DFFR_X1 \if_id/incPC_q_reg[11]  ( .D(n2212), .CK(clk), .RN(net224655), .Q(
        n2833) );
  DFFR_X1 \if_id/incPC_q_reg[13]  ( .D(n2210), .CK(clk), .RN(net224655), .Q(
        n3030) );
  DFFR_X1 \if_id/incPC_q_reg[14]  ( .D(n2208), .CK(clk), .RN(net224629), .Q(
        n3029) );
  DFFR_X1 \if_id/incPC_q_reg[15]  ( .D(n2206), .CK(clk), .RN(net224655), .Q(
        n2832) );
  DFFR_X1 \if_id/incPC_q_reg[16]  ( .D(n2204), .CK(clk), .RN(net224629), .Q(
        n3028) );
  DFFR_X1 \if_id/incPC_q_reg[17]  ( .D(n2202), .CK(clk), .RN(net224653), .Q(
        n2831) );
  DFFR_X1 \if_id/incPC_q_reg[18]  ( .D(n2200), .CK(clk), .RN(net224627), .Q(
        n2830) );
  DFFR_X1 \if_id/incPC_q_reg[19]  ( .D(n2198), .CK(clk), .RN(net224653), .Q(
        n3027) );
  DFFR_X1 \if_id/incPC_q_reg[20]  ( .D(n2196), .CK(clk), .RN(net224653), .Q(
        n3026) );
  DFFR_X1 \if_id/incPC_q_reg[21]  ( .D(n2194), .CK(clk), .RN(net224627), .Q(
        n3025) );
  DFFR_X1 \if_id/incPC_q_reg[22]  ( .D(n2192), .CK(clk), .RN(net224653), .Q(
        n3024) );
  DFFR_X1 \if_id/incPC_q_reg[23]  ( .D(n2190), .CK(clk), .RN(net224627), .Q(
        n2829) );
  DFFR_X1 \if_id/incPC_q_reg[24]  ( .D(n2188), .CK(clk), .RN(net224653), .Q(
        n3023) );
  DFFR_X1 \if_id/incPC_q_reg[25]  ( .D(n2186), .CK(clk), .RN(net224627), .Q(
        n3022) );
  DFFR_X1 \if_id/incPC_q_reg[26]  ( .D(n2184), .CK(clk), .RN(net224653), .Q(
        n3021) );
  DFFR_X1 \if_id/incPC_q_reg[27]  ( .D(n2182), .CK(clk), .RN(net224627), .Q(
        n3020) );
  DFFR_X1 \if_id/incPC_q_reg[28]  ( .D(n2180), .CK(clk), .RN(net224653), .Q(
        n3019) );
  DFFR_X1 \if_id/incPC_q_reg[29]  ( .D(n2178), .CK(clk), .RN(net224627), .Q(
        n3018) );
  DFFR_X1 \if_id/incPC_q_reg[30]  ( .D(n2176), .CK(clk), .RN(net224627), .Q(
        n2987) );
  DFFR_X1 \if_id/instr_q_reg[24]  ( .D(n2163), .CK(clk), .RN(net224627), .Q(
        rs1[3]) );
  DFFR_X1 \if_id/instr_q_reg[15]  ( .D(n2154), .CK(clk), .RN(net224661), .Q(
        n2939) );
  DFFR_X1 \if_id/instr_q_reg[14]  ( .D(n2153), .CK(clk), .RN(net224625), .Q(
        n2955) );
  DFFR_X1 \if_id/instr_q_reg[13]  ( .D(n2152), .CK(clk), .RN(net224645), .Q(
        n2956) );
  DFFR_X1 \if_id/instr_q_reg[12]  ( .D(n2151), .CK(clk), .RN(net224625), .Q(
        n2957) );
  DFFR_X1 \if_id/instr_q_reg[11]  ( .D(n2150), .CK(clk), .RN(net224657), .Q(
        n2958) );
  DFFR_X1 \if_id/instr_q_reg[10]  ( .D(n2149), .CK(clk), .RN(net224625), .Q(
        n2938) );
  DFFR_X1 \if_id/instr_q_reg[9]  ( .D(n2148), .CK(clk), .RN(net224623), .Q(
        n2936) );
  DFFR_X1 \if_id/instr_q_reg[8]  ( .D(n2147), .CK(clk), .RN(net224619), .Q(
        n2935) );
  DFFR_X1 \if_id/instr_q_reg[7]  ( .D(n2146), .CK(clk), .RN(net224623), .Q(
        n2934) );
  DFFR_X1 \if_id/instr_q_reg[6]  ( .D(n2145), .CK(clk), .RN(net224629), .Q(
        n2933) );
  DFFR_X1 \id_ex/rd_q_reg[0]  ( .D(n2138), .CK(clk), .RN(net224655), .Q(
        rd_2[0]), .QN(n2853) );
  DFFR_X1 \id_ex/setInv_q_reg  ( .D(n2135), .CK(clk), .RN(net224629), .Q(
        setInv_2), .QN(n2848) );
  DFFR_X1 \id_ex/memRd_q_reg  ( .D(n7882), .CK(clk), .RN(net224655), .QN(n7717) );
  DFFR_X1 \id_ex/branch_q_reg  ( .D(n2133), .CK(clk), .RN(net224623), .QN(
        n7644) );
  DFFR_X1 \id_ex/jr_q_reg  ( .D(n7881), .CK(clk), .RN(net224659), .QN(n7716)
         );
  DFFR_X1 \id_ex/op0_q_reg  ( .D(n2127), .CK(clk), .RN(net224619), .Q(op0_2), 
        .QN(n2945) );
  DFFR_X1 \id_ex/dSize_q_reg[0]  ( .D(n2126), .CK(clk), .RN(net224661), .Q(
        n2825) );
  DFFR_X1 \id_ex/dSize_q_reg[1]  ( .D(n2123), .CK(clk), .RN(net224671), .Q(
        n2824) );
  DFFR_X1 \id_ex/imm32_q_reg[0]  ( .D(n2120), .CK(clk), .RN(net224671), .Q(
        n2896), .QN(n7733) );
  DFFR_X1 \id_ex/imm32_q_reg[1]  ( .D(n7885), .CK(clk), .RN(net224659), .QN(
        n7749) );
  DFFR_X1 \id_ex/imm32_q_reg[2]  ( .D(n2118), .CK(clk), .RN(net224669), .QN(
        n7720) );
  DFFR_X1 \id_ex/imm32_q_reg[3]  ( .D(n7887), .CK(clk), .RN(net224659), .Q(
        n2918), .QN(n7748) );
  DFFR_X1 \id_ex/imm32_q_reg[4]  ( .D(n2116), .CK(clk), .RN(net224669), .QN(
        n7721) );
  DFFR_X1 \id_ex/imm32_q_reg[6]  ( .D(n7876), .CK(clk), .RN(net224669), .QN(
        n7746) );
  DFFR_X1 \id_ex/imm32_q_reg[7]  ( .D(n7877), .CK(clk), .RN(net224659), .QN(
        n7745) );
  DFFR_X1 \id_ex/imm32_q_reg[9]  ( .D(n7879), .CK(clk), .RN(net224659), .QN(
        n7743) );
  DFFR_X1 \id_ex/imm32_q_reg[11]  ( .D(n2109), .CK(clk), .RN(net224671), .QN(
        n7724) );
  DFFR_X1 \id_ex/imm32_q_reg[12]  ( .D(n2108), .CK(clk), .RN(net224661), .QN(
        n7725) );
  DFFR_X1 \id_ex/imm32_q_reg[13]  ( .D(n2107), .CK(clk), .RN(net224671), .Q(
        n2897), .QN(n7722) );
  DFFR_X1 \id_ex/imm32_q_reg[14]  ( .D(n2106), .CK(clk), .RN(net224661), .QN(
        n7726) );
  DFFR_X1 \id_ex/imm32_q_reg[15]  ( .D(n2105), .CK(clk), .RN(net224669), .Q(
        n2859), .QN(n7727) );
  DFFR_X1 \id_ex/imm32_q_reg[16]  ( .D(n2104), .CK(clk), .RN(net224661), .Q(
        n2932), .QN(n7742) );
  DFFR_X1 \id_ex/imm32_q_reg[17]  ( .D(n2103), .CK(clk), .RN(net224669), .Q(
        n2917), .QN(n7741) );
  DFFR_X1 \id_ex/imm32_q_reg[18]  ( .D(n2102), .CK(clk), .RN(net224661), .Q(
        n2931), .QN(n7740) );
  DFFR_X1 \id_ex/imm32_q_reg[19]  ( .D(n2101), .CK(clk), .RN(net224669), .Q(
        n2900), .QN(net33197) );
  DFFR_X1 \id_ex/imm32_q_reg[20]  ( .D(n2100), .CK(clk), .RN(net224669), .Q(
        n2901), .QN(n7739) );
  DFFR_X1 \id_ex/imm32_q_reg[21]  ( .D(n2099), .CK(clk), .RN(net224659), .Q(
        n2906), .QN(n7738) );
  DFFR_X1 \id_ex/imm32_q_reg[22]  ( .D(n2098), .CK(clk), .RN(net224669), .Q(
        n2764), .QN(n7737) );
  DFFR_X1 \id_ex/imm32_q_reg[23]  ( .D(n2097), .CK(clk), .RN(net224659), .Q(
        n2763), .QN(n7736) );
  DFFR_X1 \id_ex/imm32_q_reg[24]  ( .D(n2096), .CK(clk), .RN(net224669), .Q(
        n2773), .QN(n7735) );
  DFFR_X1 \id_ex/imm32_q_reg[25]  ( .D(n2095), .CK(clk), .RN(net224659), .Q(
        n2930), .QN(n7734) );
  DFFR_X1 \id_ex/imm32_q_reg[26]  ( .D(n2094), .CK(clk), .RN(net224669), .Q(
        n2915), .QN(n7729) );
  DFFR_X1 \id_ex/imm32_q_reg[27]  ( .D(n2093), .CK(clk), .RN(net224659), .Q(
        n2928), .QN(n7728) );
  DFFR_X1 \id_ex/imm32_q_reg[28]  ( .D(n2092), .CK(clk), .RN(net224669), .Q(
        n2913), .QN(n7731) );
  DFFR_X1 \id_ex/imm32_q_reg[29]  ( .D(n2091), .CK(clk), .RN(net224659), .Q(
        n2898), .QN(n7732) );
  DFFR_X1 \id_ex/imm32_q_reg[30]  ( .D(n2090), .CK(clk), .RN(net224659), .Q(
        n2905), .QN(n7730) );
  DFFR_X1 \id_ex/imm32_q_reg[31]  ( .D(n2089), .CK(clk), .RN(net224669), .Q(
        n2923), .QN(n7723) );
  DFFR_X1 \id_ex/rd_q_reg[1]  ( .D(n2088), .CK(clk), .RN(net224611), .Q(
        rd_2[1]), .QN(n2851) );
  DFFR_X1 \id_ex/rd_q_reg[2]  ( .D(n2086), .CK(clk), .RN(net224655), .Q(
        rd_2[2]), .QN(n2850) );
  DFFR_X1 \id_ex/rd_q_reg[3]  ( .D(n2084), .CK(clk), .RN(net224671), .Q(
        rd_2[3]), .QN(n2854) );
  DFFR_X1 \id_ex/rd_q_reg[4]  ( .D(n2083), .CK(clk), .RN(net224655), .Q(
        rd_2[4]), .QN(n2852) );
  DFFR_X1 \id_ex/busA_q_reg[0]  ( .D(n7812), .CK(clk), .RN(net224619), .Q(
        n2755) );
  DFFR_X1 \id_ex/busA_q_reg[1]  ( .D(n7811), .CK(clk), .RN(net224675), .Q(
        n2754) );
  DFFR_X1 \id_ex/busA_q_reg[6]  ( .D(n7806), .CK(clk), .RN(net224635), .Q(
        n2753) );
  DFFR_X1 \id_ex/busA_q_reg[7]  ( .D(n7805), .CK(clk), .RN(net224673), .QN(
        n7688) );
  DFFR_X1 \id_ex/busA_q_reg[18]  ( .D(n7794), .CK(clk), .RN(net224675), .Q(
        n2752) );
  DFFR_X1 \id_ex/busA_q_reg[19]  ( .D(n7793), .CK(clk), .RN(net224679), .Q(
        n2718) );
  DFFR_X1 \id_ex/busA_q_reg[20]  ( .D(n7792), .CK(clk), .RN(net224679), .Q(
        n2717) );
  DFFR_X1 \id_ex/busA_q_reg[21]  ( .D(n7791), .CK(clk), .RN(net224675), .Q(
        n7603), .QN(n7698) );
  DFFR_X1 \id_ex/busA_q_reg[22]  ( .D(n7790), .CK(clk), .RN(net224679), .Q(
        n2716) );
  DFFR_X1 \id_ex/busA_q_reg[23]  ( .D(n7789), .CK(clk), .RN(net224675), .Q(
        n2715) );
  DFFR_X1 \id_ex/busA_q_reg[25]  ( .D(n7787), .CK(clk), .RN(net224675), .Q(
        n2751) );
  DFFR_X1 \id_ex/busA_q_reg[29]  ( .D(n7783), .CK(clk), .RN(net224675), .Q(
        n2750) );
  DFFR_X1 \id_ex/busA_q_reg[31]  ( .D(n7781), .CK(clk), .RN(net224653), .Q(
        n2714) );
  DFFR_X1 \id_ex/busB_q_reg[1]  ( .D(n7843), .CK(clk), .RN(net224673), .Q(
        n2749) );
  DFFR_X1 \id_ex/busB_q_reg[2]  ( .D(n7842), .CK(clk), .RN(net224661), .Q(
        n2748) );
  DFFR_X1 \id_ex/busB_q_reg[4]  ( .D(n7840), .CK(clk), .RN(net224661), .Q(
        n2747) );
  DFFR_X1 \id_ex/busB_q_reg[5]  ( .D(n7839), .CK(clk), .RN(net224671), .Q(
        n2745), .QN(n7956) );
  DFFR_X1 \id_ex/busB_q_reg[9]  ( .D(n7835), .CK(clk), .RN(net224671), .Q(
        n2845) );
  DFFR_X1 \id_ex/busB_q_reg[12]  ( .D(n7832), .CK(clk), .RN(net224673), .Q(
        n2746) );
  DFFR_X1 \id_ex/busB_q_reg[14]  ( .D(n7830), .CK(clk), .RN(net224673), .Q(
        n2713) );
  DFFR_X1 \id_ex/busB_q_reg[17]  ( .D(n7827), .CK(clk), .RN(net224663), .Q(
        n2844) );
  DFFR_X1 \id_ex/busB_q_reg[24]  ( .D(n7820), .CK(clk), .RN(net224663), .Q(
        n2712) );
  DFFR_X1 \id_ex/busB_q_reg[28]  ( .D(n7816), .CK(clk), .RN(net224663), .Q(
        n2709) );
  DFFR_X1 \id_ex/busB_q_reg[29]  ( .D(n7815), .CK(clk), .RN(net224671), .Q(
        n2708) );
  DFFR_X1 \id_ex/aluCtrl_q_reg[2]  ( .D(n2016), .CK(clk), .RN(net224641), .Q(
        n2786), .QN(n7719) );
  DFFR_X1 \if_id/incPC_q_reg[0]  ( .D(n7863), .CK(clk), .RN(net224655), .Q(
        n2828) );
  DFFR_X1 \id_ex/incPC_q_reg[0]  ( .D(n7874), .CK(clk), .RN(net224661), .Q(
        n3034), .QN(n7715) );
  DFFR_X1 \if_id/incPC_q_reg[1]  ( .D(n7862), .CK(clk), .RN(net224627), .Q(
        n3017) );
  DFFR_X1 \id_ex/incPC_q_reg[1]  ( .D(n7873), .CK(clk), .RN(net224657), .Q(
        n2807), .QN(n7714) );
  DFFR_X1 \if_id/incPC_q_reg[2]  ( .D(n1981), .CK(clk), .RN(net224653), .Q(
        n2827) );
  DFFR_X1 \id_ex/incPC_q_reg[2]  ( .D(n1980), .CK(clk), .RN(net224639), .Q(
        n3033), .QN(n7639) );
  DFFR_X1 \if_id/incPC_q_reg[3]  ( .D(n1977), .CK(clk), .RN(net224627), .Q(
        n2705) );
  DFFR_X1 \id_ex/incPC_q_reg[3]  ( .D(n1976), .CK(clk), .RN(net224657), .Q(
        n2834), .QN(n7638) );
  DFFR_X1 \if_id/incPC_q_reg[4]  ( .D(n1973), .CK(clk), .RN(net224653), .Q(
        n2722) );
  DFFR_X1 \id_ex/incPC_q_reg[4]  ( .D(n1972), .CK(clk), .RN(net224641), .Q(
        n2806), .QN(n7637) );
  DFFR_X1 \if_id/incPC_q_reg[6]  ( .D(n1969), .CK(clk), .RN(net224653), .Q(
        n3016) );
  DFFR_X1 \id_ex/incPC_q_reg[6]  ( .D(n1968), .CK(clk), .RN(net224671), .Q(
        n2805), .QN(n7636) );
  DFFR_X1 \if_id/incPC_q_reg[7]  ( .D(n1966), .CK(clk), .RN(net224627), .Q(
        n3015) );
  DFFR_X1 \if_id/incPC_q_reg[8]  ( .D(n1963), .CK(clk), .RN(net224653), .Q(
        n3014) );
  DFFR_X1 \if_id/incPC_q_reg[9]  ( .D(n1960), .CK(clk), .RN(net224627), .Q(
        n2826) );
  DFFR_X1 \id_ex/incPC_q_reg[9]  ( .D(n1959), .CK(clk), .RN(net224655), .Q(
        n3032), .QN(n7633) );
  DFFR_X1 \if_id/incPC_q_reg[12]  ( .D(n1957), .CK(clk), .RN(net224629), .Q(
        n3013) );
  DFFR_X1 \if_id/incPC_q_reg[5]  ( .D(n1946), .CK(clk), .RN(net224627), .Q(
        n2721) );
  DFFR_X1 \if_id/incPC_q_reg[31]  ( .D(n1917), .CK(clk), .RN(net224653), .Q(
        n3012) );
  DFFR_X1 \id_ex/incPC_q_reg[31]  ( .D(n1916), .CK(clk), .RN(net224643), .Q(
        n2800), .QN(n7629) );
  DFFS_X2 \id_ex/instr_q_reg[4]  ( .D(n7884), .CK(clk), .SN(net224681), .Q(
        instr_2[4]) );
  DFFS_X2 \id_ex/instr_q_reg[2]  ( .D(n7886), .CK(clk), .SN(net224681), .Q(
        instr_2[2]) );
  DFFS_X2 \id_ex/not_trap_q_reg  ( .D(\id_ex/N45 ), .CK(clk), .SN(net224681), 
        .QN(n7579) );
  DFFS_X2 \ex_mem/not_trap_q_reg  ( .D(\ex_mem/N242 ), .CK(clk), .SN(net224681), .QN(n3040) );
  DFFS_X2 \id_ex/instr_q_reg[0]  ( .D(\id_ex/N4 ), .CK(clk), .SN(net224679), 
        .Q(instr_2[0]) );
  DFF_X2 \mem_wb/memRdData_q_reg[0]  ( .D(n2267), .CK(clk), .Q(
        \wb/dsize_reg/z2 [0]), .QN(n2727) );
  DFF_X2 \mem_wb/memRdData_q_reg[1]  ( .D(n2266), .CK(clk), .Q(
        \wb/dsize_reg/z2 [1]), .QN(n2785) );
  DFF_X2 \mem_wb/memRdData_q_reg[2]  ( .D(n2265), .CK(clk), .Q(
        \wb/dsize_reg/z2 [2]), .QN(n2780) );
  DFF_X2 \mem_wb/memRdData_q_reg[3]  ( .D(n2264), .CK(clk), .Q(
        \wb/dsize_reg/z2 [3]), .QN(n3772) );
  DFF_X2 \mem_wb/memRdData_q_reg[4]  ( .D(n2263), .CK(clk), .Q(
        \wb/dsize_reg/z2 [4]), .QN(n2777) );
  DFF_X2 \mem_wb/memRdData_q_reg[5]  ( .D(n2262), .CK(clk), .Q(
        \wb/dsize_reg/z2 [5]), .QN(n2779) );
  DFF_X2 \mem_wb/memRdData_q_reg[6]  ( .D(n2261), .CK(clk), .Q(
        \wb/dsize_reg/z2 [6]), .QN(n3010) );
  DFF_X2 \mem_wb/memRdData_q_reg[7]  ( .D(n2260), .CK(clk), .Q(
        \wb/dsize_reg/z2 [7]), .QN(n2783) );
  DFF_X2 \mem_wb/memRdData_q_reg[8]  ( .D(n2259), .CK(clk), .Q(
        \wb/dsize_reg/z2 [8]), .QN(n2949) );
  DFF_X2 \mem_wb/memRdData_q_reg[9]  ( .D(n2258), .CK(clk), .Q(
        \wb/dsize_reg/z2 [9]), .QN(n2927) );
  DFF_X2 \mem_wb/memRdData_q_reg[10]  ( .D(n2257), .CK(clk), .Q(
        \wb/dsize_reg/z2 [10]), .QN(n2964) );
  DFF_X2 \mem_wb/memRdData_q_reg[11]  ( .D(n2256), .CK(clk), .Q(
        \wb/dsize_reg/z2 [11]), .QN(n2947) );
  DFF_X2 \mem_wb/memRdData_q_reg[12]  ( .D(n2255), .CK(clk), .Q(
        \wb/dsize_reg/z2 [12]), .QN(n2948) );
  DFF_X2 \mem_wb/memRdData_q_reg[13]  ( .D(n2254), .CK(clk), .Q(
        \wb/dsize_reg/z2 [13]), .QN(n3078) );
  DFF_X2 \mem_wb/memRdData_q_reg[14]  ( .D(n2253), .CK(clk), .Q(
        \wb/dsize_reg/z2 [14]), .QN(n2782) );
  DFF_X2 \mem_wb/memRdData_q_reg[15]  ( .D(n2252), .CK(clk), .Q(
        \wb/dsize_reg/z2 [15]), .QN(n2967) );
  DFF_X2 \mem_wb/memRdData_q_reg[16]  ( .D(n2251), .CK(clk), .Q(
        \wb/dsize_reg/z2 [16]), .QN(n2737) );
  DFF_X2 \mem_wb/memRdData_q_reg[17]  ( .D(n2250), .CK(clk), .Q(
        \wb/dsize_reg/z2 [17]), .QN(n2726) );
  DFF_X2 \mem_wb/memRdData_q_reg[18]  ( .D(n2249), .CK(clk), .Q(
        \wb/dsize_reg/z2 [18]), .QN(n2734) );
  DFF_X2 \mem_wb/memRdData_q_reg[19]  ( .D(n2248), .CK(clk), .Q(
        \wb/dsize_reg/z2 [19]), .QN(n2735) );
  DFF_X2 \mem_wb/memRdData_q_reg[20]  ( .D(n2247), .CK(clk), .Q(
        \wb/dsize_reg/z2 [20]), .QN(n2728) );
  DFF_X2 \mem_wb/memRdData_q_reg[21]  ( .D(n2246), .CK(clk), .Q(
        \wb/dsize_reg/z2 [21]), .QN(n2736) );
  DFF_X2 \mem_wb/memRdData_q_reg[22]  ( .D(n2245), .CK(clk), .Q(
        \wb/dsize_reg/z2 [22]), .QN(n2732) );
  DFF_X2 \mem_wb/memRdData_q_reg[23]  ( .D(n2244), .CK(clk), .Q(
        \wb/dsize_reg/z2 [23]), .QN(n2729) );
  DFF_X2 \mem_wb/memRdData_q_reg[24]  ( .D(n2243), .CK(clk), .Q(
        \wb/dsize_reg/z2 [24]), .QN(n2730) );
  DFF_X2 \mem_wb/memRdData_q_reg[25]  ( .D(n2242), .CK(clk), .Q(
        \wb/dsize_reg/z2 [25]), .QN(n2733) );
  DFF_X2 \mem_wb/memRdData_q_reg[26]  ( .D(n2241), .CK(clk), .Q(
        \wb/dsize_reg/z2 [26]), .QN(n2719) );
  DFF_X2 \mem_wb/memRdData_q_reg[27]  ( .D(n2240), .CK(clk), .Q(
        \wb/dsize_reg/z2 [27]), .QN(n2784) );
  DFF_X2 \mem_wb/memRdData_q_reg[28]  ( .D(n2239), .CK(clk), .Q(
        \wb/dsize_reg/z2 [28]), .QN(n2787) );
  DFF_X2 \mem_wb/memRdData_q_reg[29]  ( .D(n2238), .CK(clk), .Q(
        \wb/dsize_reg/z2 [29]), .QN(n2791) );
  DFF_X2 \mem_wb/memRdData_q_reg[30]  ( .D(n2237), .CK(clk), .Q(
        \wb/dsize_reg/z2 [30]), .QN(n2781) );
  DFF_X2 \mem_wb/memRdData_q_reg[31]  ( .D(n2236), .CK(clk), .Q(
        \wb/dsize_reg/z2 [31]), .QN(n2731) );
  DFF_X2 \mem_wb/aluRes_q_reg[0]  ( .D(n2235), .CK(clk), .QN(n7578) );
  DFF_X2 \mem_wb/aluRes_q_reg[16]  ( .D(n7774), .CK(clk), .Q(n2992), .QN(n7577) );
  DFF_X2 \mem_wb/aluRes_q_reg[21]  ( .D(n7770), .CK(clk), .Q(n3077), .QN(n7576) );
  DFF_X2 \mem_wb/aluRes_q_reg[22]  ( .D(n7769), .CK(clk), .QN(n7575) );
  DFF_X2 \mem_wb/aluRes_q_reg[23]  ( .D(n7768), .CK(clk), .QN(n7574) );
  DFF_X2 \mem_wb/aluRes_q_reg[24]  ( .D(n7767), .CK(clk), .Q(n2977), .QN(n7573) );
  DFF_X2 \mem_wb/aluRes_q_reg[25]  ( .D(n7766), .CK(clk), .Q(n3090), .QN(n7572) );
  DFF_X2 \mem_wb/aluRes_q_reg[31]  ( .D(n7760), .CK(clk), .QN(n7571) );
  DFF_X2 \mem_wb/aluRes_q_reg[4]  ( .D(n2227), .CK(clk), .Q(n3122), .QN(n7570)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[9]  ( .D(n7758), .CK(clk), .QN(n7569) );
  DFF_X2 \mem_wb/aluRes_q_reg[2]  ( .D(n2225), .CK(clk), .Q(n2651), .QN(n7568)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[1]  ( .D(n2224), .CK(clk), .QN(n7567) );
  DFF_X2 \mem_wb/aluRes_q_reg[3]  ( .D(n2223), .CK(clk), .QN(n7566) );
  DFF_X2 \mem_wb/aluRes_q_reg[6]  ( .D(n2222), .CK(clk), .Q(n2966), .QN(n7565)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[11]  ( .D(n7779), .CK(clk), .QN(n7564) );
  DFF_X2 \mem_wb/aluRes_q_reg[7]  ( .D(n2220), .CK(clk), .Q(n3118), .QN(n7563)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[29]  ( .D(n7762), .CK(clk), .QN(n7562) );
  DFF_X2 \mem_wb/aluRes_q_reg[8]  ( .D(n7759), .CK(clk), .Q(n3096), .QN(n7561)
         );
  DFF_X2 \mem_wb/aluRes_q_reg[12]  ( .D(n7778), .CK(clk), .QN(n7560) );
  DFF_X2 \mem_wb/aluRes_q_reg[13]  ( .D(n7777), .CK(clk), .Q(n3086), .QN(n7559) );
  DFF_X2 \mem_wb/aluRes_q_reg[10]  ( .D(n7780), .CK(clk), .Q(n2979), .QN(n7558) );
  DFF_X2 \mem_wb/aluRes_q_reg[30]  ( .D(n7761), .CK(clk), .QN(n7557) );
  DFF_X2 \mem_wb/aluRes_q_reg[19]  ( .D(net33021), .CK(clk), .QN(net35052) );
  DFFS_X2 \if_id/instr_q_reg[4]  ( .D(n2143), .CK(clk), .SN(net224679), .Q(
        n2870), .QN(n7556) );
  DFFS_X2 \if_id/instr_q_reg[2]  ( .D(n2141), .CK(clk), .SN(net224679), .Q(
        n2765), .QN(n7555) );
  DFFS_X2 \if_id/instr_q_reg[0]  ( .D(n2139), .CK(clk), .SN(net224679), .Q(
        n2766), .QN(n7554) );
  DFF_X2 \mem_wb/fp_q_reg  ( .D(n2128), .CK(clk), .Q(net229988), .QN(net35047)
         );
  DFF_X2 \ex_mem/dSize_q_reg[0]  ( .D(n2125), .CK(clk), .Q(dSize[0]) );
  DFF_X2 \mem_wb/dSize_q_reg[0]  ( .D(n2124), .CK(clk), .QN(n7553) );
  DFF_X2 \ex_mem/dSize_q_reg[1]  ( .D(n2122), .CK(clk), .Q(dSize[1]) );
  DFF_X2 \mem_wb/dSize_q_reg[1]  ( .D(n2121), .CK(clk), .Q(n2843), .QN(n7552)
         );
  DFF_X2 \mem_wb/rd_q_reg[1]  ( .D(n7755), .CK(clk), .Q(rd[1]) );
  DFF_X2 \mem_wb/rd_q_reg[2]  ( .D(n7754), .CK(clk), .Q(rd[2]) );
  DFFRS_X2 \ifetch/dffa/q_reg[16]  ( .D(n2001), .CK(clk), .RN(n1886), .SN(
        n1885), .Q(n3129), .QN(n7671) );
  DFF_X2 \mem_wb/rd_q_reg[0]  ( .D(n7756), .CK(clk), .Q(rd[0]) );
  DFF_X2 \mem_wb/rd_q_reg[4]  ( .D(n7752), .CK(clk), .Q(rd[4]) );
  DFF_X2 \mem_wb/rd_q_reg[3]  ( .D(n7753), .CK(clk), .Q(rd[3]) );
  DFF_X2 \mem_wb/link_q_reg  ( .D(n1992), .CK(clk), .Q(net228233), .QN(
        net35037) );
  DFF_X2 \mem_wb/memRd_q_reg  ( .D(n7757), .CK(clk), .Q(n3127), .QN(net35036)
         );
  DFFRS_X2 \ifetch/dffa/q_reg[0]  ( .D(n1990), .CK(clk), .RN(n1874), .SN(n1873), .QN(n7641) );
  DFF_X2 \mem_wb/reg31Val_q_reg[0]  ( .D(n7751), .CK(clk), .Q(reg31Val_0[0])
         );
  DFFRS_X2 \ifetch/dffa/q_reg[1]  ( .D(n1986), .CK(clk), .RN(n1872), .SN(n1871), .QN(n7640) );
  DFF_X2 \mem_wb/reg31Val_q_reg[1]  ( .D(n7750), .CK(clk), .Q(reg31Val_0[1])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[2]  ( .D(n1979), .CK(clk), .Q(reg31Val_0[2])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[3]  ( .D(n1975), .CK(clk), .Q(reg31Val_0[3]), 
        .QN(n3087) );
  DFF_X2 \mem_wb/reg31Val_q_reg[4]  ( .D(n1971), .CK(clk), .Q(reg31Val_0[4])
         );
  DFFRS_X2 \ifetch/dffa/q_reg[8]  ( .D(n1964), .CK(clk), .RN(n1860), .SN(n1859), .Q(n3131), .QN(n7673) );
  DFF_X2 \mem_wb/reg31Val_q_reg[29]  ( .D(n1955), .CK(clk), .Q(reg31Val_0[29]), 
        .QN(n2981) );
  DFF_X2 \mem_wb/reg31Val_q_reg[28]  ( .D(n1954), .CK(clk), .Q(reg31Val_0[28]), 
        .QN(n3081) );
  DFF_X2 \mem_wb/aluRes_q_reg[28]  ( .D(n7763), .CK(clk), .QN(n7551) );
  DFF_X2 \mem_wb/reg31Val_q_reg[27]  ( .D(n1952), .CK(clk), .Q(reg31Val_0[27]), 
        .QN(n2916) );
  DFF_X2 \mem_wb/aluRes_q_reg[27]  ( .D(n7764), .CK(clk), .Q(n2925), .QN(n7550) );
  DFF_X2 \mem_wb/reg31Val_q_reg[26]  ( .D(n1950), .CK(clk), .Q(reg31Val_0[26]), 
        .QN(n2960) );
  DFF_X2 \mem_wb/aluRes_q_reg[26]  ( .D(n7765), .CK(clk), .Q(n2976), .QN(n7549) );
  DFF_X2 \mem_wb/aluRes_q_reg[5]  ( .D(n1948), .CK(clk), .Q(n3079), .QN(n7548)
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[6]  ( .D(n1944), .CK(clk), .Q(reg31Val_0[6])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[5]  ( .D(n1943), .CK(clk), .Q(reg31Val_0[5])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[8]  ( .D(n1942), .CK(clk), .Q(reg31Val_0[8]), 
        .QN(n2959) );
  DFF_X2 \mem_wb/reg31Val_q_reg[7]  ( .D(n1941), .CK(clk), .Q(reg31Val_0[7])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[9]  ( .D(n1940), .CK(clk), .Q(reg31Val_0[9])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[11]  ( .D(n1939), .CK(clk), .Q(reg31Val_0[11])
         );
  DFF_X2 \mem_wb/reg31Val_q_reg[10]  ( .D(n1938), .CK(clk), .Q(reg31Val_0[10]), 
        .QN(n3083) );
  DFF_X2 \mem_wb/reg31Val_q_reg[25]  ( .D(n1937), .CK(clk), .Q(reg31Val_0[25]), 
        .QN(n2983) );
  DFF_X2 \mem_wb/reg31Val_q_reg[24]  ( .D(n1936), .CK(clk), .Q(reg31Val_0[24]), 
        .QN(n2982) );
  DFF_X2 \mem_wb/reg31Val_q_reg[23]  ( .D(n1935), .CK(clk), .Q(reg31Val_0[23]), 
        .QN(n3080) );
  DFF_X2 \mem_wb/reg31Val_q_reg[22]  ( .D(n1934), .CK(clk), .Q(reg31Val_0[22]), 
        .QN(n2792) );
  DFF_X2 \mem_wb/reg31Val_q_reg[21]  ( .D(n1933), .CK(clk), .Q(reg31Val_0[21]), 
        .QN(n3075) );
  DFF_X2 \mem_wb/reg31Val_q_reg[20]  ( .D(n1932), .CK(clk), .Q(reg31Val_0[20]), 
        .QN(n2950) );
  DFF_X2 \mem_wb/reg31Val_q_reg[19]  ( .D(n1931), .CK(clk), .Q(reg31Val_0[19]), 
        .QN(n2937) );
  DFF_X2 \mem_wb/reg31Val_q_reg[18]  ( .D(n1930), .CK(clk), .Q(reg31Val_0[18]), 
        .QN(n2974) );
  DFF_X2 \mem_wb/reg31Val_q_reg[17]  ( .D(n1929), .CK(clk), .Q(reg31Val_0[17]), 
        .QN(n3082) );
  DFF_X2 \mem_wb/reg31Val_q_reg[16]  ( .D(n1928), .CK(clk), .Q(reg31Val_0[16]), 
        .QN(n3076) );
  DFF_X2 \mem_wb/reg31Val_q_reg[15]  ( .D(n1927), .CK(clk), .Q(reg31Val_0[15]), 
        .QN(n3126) );
  DFF_X2 \mem_wb/reg31Val_q_reg[14]  ( .D(n1926), .CK(clk), .Q(reg31Val_0[14])
         );
  DFF_X2 \mem_wb/aluRes_q_reg[14]  ( .D(n7776), .CK(clk), .Q(n2799), .QN(n7547) );
  DFF_X2 \mem_wb/aluRes_q_reg[20]  ( .D(n7771), .CK(clk), .QN(n7546) );
  DFF_X2 \mem_wb/aluRes_q_reg[15]  ( .D(n7775), .CK(clk), .QN(n7545) );
  DFF_X2 \mem_wb/aluRes_q_reg[18]  ( .D(n7772), .CK(clk), .Q(n3089), .QN(n7544) );
  DFF_X2 \mem_wb/aluRes_q_reg[17]  ( .D(n7773), .CK(clk), .Q(n3121), .QN(n7543) );
  DFF_X2 \mem_wb/reg31Val_q_reg[13]  ( .D(n1920), .CK(clk), .Q(reg31Val_0[13]), 
        .QN(n2837) );
  DFF_X2 \mem_wb/reg31Val_q_reg[12]  ( .D(n1919), .CK(clk), .Q(reg31Val_0[12])
         );
  DFFR_X2 \id_ex/busB_sel_q_reg[0]  ( .D(\id_ex/N40 ), .CK(clk), .RN(net224629), .Q(net229071), .QN(net34726) );
  DFFR_X2 \id_ex/busB_sel_q_reg[1]  ( .D(\id_ex/N41 ), .CK(clk), .RN(net224627), .Q(net225520), .QN(net34717) );
  DFFR_X2 \if_id/instr_q_reg[26]  ( .D(n2165), .CK(clk), .RN(net224669), .Q(
        op0_1), .QN(n2846) );
  DFFR_X2 \id_ex/aluCtrl_q_reg[1]  ( .D(n2017), .CK(clk), .RN(net224639), .Q(
        n2839), .QN(net33219) );
  DFFR_X2 \ex_mem/incPC_q_reg[2]  ( .D(\ex_mem/N37 ), .CK(clk), .RN(net224641), 
        .QN(n7433) );
  DFFR_X2 \ex_mem/incPC_q_reg[3]  ( .D(\ex_mem/N38 ), .CK(clk), .RN(net224639), 
        .Q(n3070), .QN(n7432) );
  DFFR_X2 \ex_mem/incPC_q_reg[9]  ( .D(\ex_mem/N44 ), .CK(clk), .RN(net224639), 
        .Q(n3173), .QN(n7426) );
  DFFR_X2 \ex_mem/incPC_q_reg[11]  ( .D(\ex_mem/N46 ), .CK(clk), .RN(net224619), .Q(n3723), .QN(n7519) );
  DFFR_X2 \id_ex/aluSrc_q_reg  ( .D(n2136), .CK(clk), .RN(net224643), .Q(
        net225434), .QN(net33207) );
  DFFR_X2 \id_ex/busA_sel_q_reg[1]  ( .D(n3125), .CK(clk), .RN(net224619), 
        .QN(n7476) );
  DFFR_X2 \id_ex/busA_sel_q_reg[0]  ( .D(\id_ex/N38 ), .CK(clk), .RN(net224615), .QN(n7496) );
  DFFR_X2 \ex_mem/incPC_q_reg[8]  ( .D(\ex_mem/N43 ), .CK(clk), .RN(net224639), 
        .Q(n2744), .QN(n7427) );
  DFFR_X2 \if_id/instr_q_reg[27]  ( .D(n2166), .CK(clk), .RN(net224625), .QN(
        n7709) );
  DFFR_X2 \ex_mem/imm32_q_reg[11]  ( .D(\ex_mem/N142 ), .CK(clk), .RN(
        net224643), .Q(n3149), .QN(n7447) );
  DFFR_X2 \ex_mem/incPC_q_reg[6]  ( .D(\ex_mem/N41 ), .CK(clk), .RN(net224639), 
        .Q(n2741), .QN(n7429) );
  DFFR_X2 \ex_mem/imm32_q_reg[6]  ( .D(\ex_mem/N137 ), .CK(clk), .RN(net224641), .Q(n2988), .QN(n7442) );
  DFFR_X2 \ex_mem/incPC_q_reg[17]  ( .D(\ex_mem/N52 ), .CK(clk), .RN(net224619), .Q(n3177), .QN(n7514) );
  DFFR_X2 \id_ex/aluCtrl_q_reg[0]  ( .D(n2018), .CK(clk), .RN(net224615), .Q(
        n2841), .QN(net33205) );
  DFFR_X2 \ex_mem/aluRes_q_reg[3]  ( .D(\ex_mem/N198 ), .CK(clk), .RN(
        net224621), .Q(memAddr[3]), .QN(n7530) );
  DFFR_X2 \ex_mem/incPC_q_reg[1]  ( .D(\ex_mem/N36 ), .CK(clk), .RN(net224641), 
        .Q(reg31Val_3[1]), .QN(n3385) );
  DFFR_X2 \id_ex/zeroExt_q_reg  ( .D(n2702), .CK(clk), .RN(net224615), .Q(
        zeroExt_2), .QN(n3133) );
  DFFR_X2 \ex_mem/incPC_q_reg[4]  ( .D(\ex_mem/N39 ), .CK(clk), .RN(net224639), 
        .Q(n2793), .QN(n7431) );
  DFF_X1 \mem_wb/reg31Val_q_reg[31]  ( .D(n1915), .CK(clk), .Q(reg31Val_0[31]), 
        .QN(n2951) );
  DFFR_X2 \id_ex/busB_q_reg[15]  ( .D(n7829), .CK(clk), .RN(net224663), .QN(
        net33276) );
  DFFR_X2 \ex_mem/aluRes_q_reg[19]  ( .D(\ex_mem/N215 ), .CK(clk), .RN(
        net224615), .Q(memAddr[19]), .QN(net34763) );
  DFFR_X2 \mem_wb/regWr_q_reg  ( .D(\mem_wb/N36 ), .CK(clk), .RN(net224625), 
        .Q(net230040), .QN(net225580) );
  DFFR_X2 \ex_mem/imm32_q_reg[18]  ( .D(\ex_mem/N149 ), .CK(clk), .RN(
        net224643), .QN(n7454) );
  DFFR_X2 \ex_mem/incPC_q_reg[18]  ( .D(\ex_mem/N53 ), .CK(clk), .RN(net224619), .QN(n7513) );
  DFFR_X2 \if_id/instr_q_reg[28]  ( .D(n2167), .CK(clk), .RN(net224675), .Q(
        n2855), .QN(n7707) );
  DFFR_X2 \ex_mem/incPC_q_reg[19]  ( .D(\ex_mem/N54 ), .CK(clk), .RN(net224619), .Q(n2778), .QN(n7512) );
  DFFR_X2 \ex_mem/imm32_q_reg[17]  ( .D(\ex_mem/N148 ), .CK(clk), .RN(
        net224643), .QN(n7453) );
  DFFR_X2 \ex_mem/incPC_q_reg[10]  ( .D(\ex_mem/N45 ), .CK(clk), .RN(net224619), .Q(n2921), .QN(n7520) );
  DFFR_X2 \ex_mem/incPC_q_reg[16]  ( .D(\ex_mem/N51 ), .CK(clk), .RN(net224619), .QN(n7515) );
  DFFR_X2 \ex_mem/imm32_q_reg[9]  ( .D(\ex_mem/N140 ), .CK(clk), .RN(net224643), .QN(n7445) );
  DFFR_X2 \ex_mem/incPC_q_reg[20]  ( .D(\ex_mem/N55 ), .CK(clk), .RN(net224617), .Q(n2762), .QN(n7511) );
  DFFR_X2 \if_id/instr_q_reg[31]  ( .D(n2170), .CK(clk), .RN(net224655), .Q(
        n2849), .QN(n7708) );
  DFFR_X2 \ex_mem/imm32_q_reg[10]  ( .D(\ex_mem/N141 ), .CK(clk), .RN(
        net224643), .QN(n7446) );
  DFFR_X2 \ex_mem/imm32_q_reg[16]  ( .D(\ex_mem/N147 ), .CK(clk), .RN(
        net224643), .QN(n7452) );
  DFFR_X2 \ex_mem/incPC_q_reg[22]  ( .D(\ex_mem/N57 ), .CK(clk), .RN(net224617), .Q(n3162), .QN(n7509) );
  DFFR_X2 \ex_mem/isZero_q_reg  ( .D(\ex_mem/N232 ), .CK(clk), .RN(net224615), 
        .QN(n7499) );
  DFFRS_X1 \ifetch/dffa/q_reg[27]  ( .D(n2012), .CK(clk), .RN(n1908), .SN(
        n1907), .Q(n3050) );
  DFF_X1 \mem_wb/reg31Val_q_reg[30]  ( .D(n2174), .CK(clk), .Q(reg31Val_0[30])
         );
  DFFRS_X1 \ifetch/dffa/q_reg[25]  ( .D(n2010), .CK(clk), .RN(n1904), .SN(
        n1903), .Q(n3045) );
  DFFRS_X1 \ifetch/dffa/q_reg[29]  ( .D(n2014), .CK(clk), .RN(n1912), .SN(
        n1911), .Q(n3048) );
  DFFRS_X1 \ifetch/dffa/q_reg[31]  ( .D(n1918), .CK(clk), .RN(n1852), .SN(
        n1851), .Q(n2985), .QN(n7630) );
  DFFR_X2 \ex_mem/imm32_q_reg[1]  ( .D(\ex_mem/N132 ), .CK(clk), .RN(net224641), .Q(n3093), .QN(n7437) );
  DFFR_X2 \ex_mem/imm32_q_reg[20]  ( .D(\ex_mem/N151 ), .CK(clk), .RN(
        net224645), .Q(n3097), .QN(n7456) );
  DFFR_X2 \ex_mem/incPC_q_reg[23]  ( .D(\ex_mem/N58 ), .CK(clk), .RN(net224617), .Q(n2965), .QN(n7508) );
  DFFR_X2 \ex_mem/incPC_q_reg[0]  ( .D(\ex_mem/N35 ), .CK(clk), .RN(net224641), 
        .Q(reg31Val_3[0]) );
  DFFRS_X1 \ifetch/dffa/q_reg[30]  ( .D(n2015), .CK(clk), .RN(n1914), .SN(
        n1913), .Q(n3047) );
  DFFR_X2 \if_id/instr_q_reg[29]  ( .D(n2168), .CK(clk), .RN(net224625), .Q(
        n2868), .QN(n7710) );
  DFFRS_X1 \ifetch/dffa/q_reg[23]  ( .D(n2008), .CK(clk), .RN(n1900), .SN(
        n1899), .Q(n3046) );
  DFFRS_X1 \ifetch/dffa/q_reg[20]  ( .D(n2005), .CK(clk), .RN(n1894), .SN(
        n1893), .Q(n3009), .QN(n7670) );
  DFFRS_X1 \ifetch/dffa/q_reg[14]  ( .D(n1999), .CK(clk), .RN(n1882), .SN(
        n1881), .Q(n3043) );
  DFFRS_X1 \ifetch/dffa/q_reg[22]  ( .D(n2007), .CK(clk), .RN(n1898), .SN(
        n1897), .Q(n3051) );
  DFFRS_X1 \ifetch/dffa/q_reg[15]  ( .D(n2000), .CK(clk), .RN(n1884), .SN(
        n1883), .Q(n2984), .QN(n7672) );
  DFFRS_X1 \ifetch/dffa/q_reg[28]  ( .D(n2013), .CK(clk), .RN(n1910), .SN(
        n1909), .Q(n3049) );
  DFFRS_X1 \ifetch/dffa/q_reg[19]  ( .D(n2004), .CK(clk), .RN(n1892), .SN(
        n1891), .Q(n3044) );
  DFFR_X2 \id_ex/busB_q_reg[8]  ( .D(n7836), .CK(clk), .RN(net224661), .QN(
        n7674) );
  DFFR_X2 \ex_mem/imm32_q_reg[19]  ( .D(\ex_mem/N150 ), .CK(clk), .RN(
        net224645), .Q(n3002), .QN(n7455) );
  DFFR_X2 \id_ex/busB_q_reg[3]  ( .D(n7841), .CK(clk), .RN(net224671), .Q(
        n2924), .QN(n7675) );
  DFFR_X2 \id_ex/imm32_q_reg[10]  ( .D(n7880), .CK(clk), .RN(net224661), .Q(
        n2902), .QN(net33193) );
  DFFR_X2 \id_ex/busB_q_reg[7]  ( .D(n7837), .CK(clk), .RN(net224671), .Q(
        n2869) );
  DFFR_X2 \id_ex/busB_q_reg[6]  ( .D(n7838), .CK(clk), .RN(net224661), .Q(
        n2760) );
  DFFR_X2 \id_ex/busB_q_reg[11]  ( .D(n7833), .CK(clk), .RN(net224663), .Q(
        n2743) );
  DFFR_X2 \id_ex/busB_q_reg[13]  ( .D(n7831), .CK(clk), .RN(net224663), .Q(
        n2742) );
  DFFR_X2 \id_ex/busB_q_reg[10]  ( .D(n7834), .CK(clk), .RN(net224673), .Q(
        n2711) );
  DFFR_X2 \id_ex/busB_q_reg[23]  ( .D(n7821), .CK(clk), .RN(net224673), .Q(
        n2710) );
  DFFR_X2 \id_ex/busB_q_reg[30]  ( .D(n7814), .CK(clk), .RN(net224671), .Q(
        n2707) );
  DFFR_X2 \id_ex/aluCtrl_q_reg[3]  ( .D(n2137), .CK(clk), .RN(net224671), .Q(
        n2704), .QN(net33204) );
  NOR2_X2 U2578 ( .A1(n4764), .A2(n4763), .ZN(n5115) );
  CLKBUF_X2 U2579 ( .A(n3250), .Z(n2576) );
  NOR2_X2 U2580 ( .A1(n3495), .A2(n5217), .ZN(n5221) );
  NAND3_X1 U2582 ( .A1(n3540), .A2(n6402), .A3(n6403), .ZN(n2577) );
  INV_X1 U2583 ( .A(n5710), .ZN(n2578) );
  AND3_X4 U2584 ( .A1(n5010), .A2(n5015), .A3(net224993), .ZN(n3495) );
  AOI21_X2 U2585 ( .B1(n3295), .B2(net220885), .A(net228940), .ZN(net221892)
         );
  NAND2_X2 U2586 ( .A1(n6883), .A2(net228941), .ZN(n6899) );
  NOR2_X4 U2587 ( .A1(net220753), .A2(n6983), .ZN(n6987) );
  CLKBUF_X2 U2588 ( .A(n5187), .Z(n2579) );
  NAND2_X2 U2589 ( .A1(n3708), .A2(n4927), .ZN(n2580) );
  NAND2_X1 U2591 ( .A1(n5948), .A2(n5967), .ZN(n5956) );
  NAND2_X2 U2593 ( .A1(n5095), .A2(net224995), .ZN(n2581) );
  NAND3_X1 U2596 ( .A1(n5499), .A2(n3133), .A3(n3944), .ZN(n5501) );
  NAND3_X1 U2597 ( .A1(regWrData[2]), .A2(n3133), .A3(n3945), .ZN(n5572) );
  INV_X4 U2598 ( .A(n6955), .ZN(n6957) );
  INV_X4 U2600 ( .A(net220882), .ZN(net228816) );
  AND3_X4 U2601 ( .A1(reg31Val_0[16]), .A2(net224781), .A3(n3898), .ZN(n4727)
         );
  NOR2_X2 U2602 ( .A1(n4773), .A2(net225051), .ZN(n4775) );
  INV_X1 U2603 ( .A(n4892), .ZN(n5155) );
  MUX2_X2 U2604 ( .A(n2897), .B(n5071), .S(net224735), .Z(n2582) );
  INV_X8 U2605 ( .A(n3675), .ZN(n5048) );
  OAI211_X4 U2606 ( .C1(n3676), .C2(n3291), .A(n3677), .B(n3678), .ZN(n3675)
         );
  OAI21_X4 U2607 ( .B1(n6925), .B2(n6924), .A(n6923), .ZN(n2583) );
  AOI21_X4 U2608 ( .B1(n6922), .B2(n3358), .A(n3254), .ZN(n6923) );
  NAND2_X4 U2609 ( .A1(n5554), .A2(n3383), .ZN(n3503) );
  NAND2_X2 U2610 ( .A1(n5415), .A2(n5414), .ZN(n2584) );
  AOI21_X2 U2612 ( .B1(n5601), .B2(n5605), .A(net224745), .ZN(n5604) );
  OAI21_X1 U2613 ( .B1(n5681), .B2(n3940), .A(n5680), .ZN(n2585) );
  INV_X8 U2615 ( .A(n6798), .ZN(n6751) );
  NAND2_X1 U2616 ( .A1(n5344), .A2(n5120), .ZN(n5122) );
  MUX2_X2 U2617 ( .A(n5372), .B(n7746), .S(net225434), .Z(n2586) );
  XNOR2_X2 U2618 ( .A(n7029), .B(n2642), .ZN(n6067) );
  INV_X8 U2619 ( .A(n6066), .ZN(n7029) );
  NAND2_X4 U2621 ( .A1(n6349), .A2(net225029), .ZN(n5675) );
  NOR2_X4 U2623 ( .A1(n2590), .A2(n2589), .ZN(n2588) );
  INV_X32 U2624 ( .A(n2641), .ZN(n2589) );
  AND2_X2 U2626 ( .A1(n5401), .A2(n5400), .ZN(n2591) );
  AND2_X2 U2627 ( .A1(net225242), .A2(net35542), .ZN(net223300) );
  XNOR2_X1 U2628 ( .A(n3833), .B(n6685), .ZN(n6680) );
  INV_X2 U2629 ( .A(n3745), .ZN(n2592) );
  INV_X2 U2630 ( .A(n3241), .ZN(n3745) );
  NOR2_X2 U2631 ( .A1(n6525), .A2(n3662), .ZN(n6529) );
  INV_X8 U2632 ( .A(net228495), .ZN(net230097) );
  NAND2_X1 U2633 ( .A1(net225237), .A2(n3089), .ZN(n4897) );
  OAI221_X1 U2634 ( .B1(n7702), .B2(n2578), .C1(n3942), .C2(n5110), .A(n5109), 
        .ZN(n2593) );
  NAND2_X1 U2635 ( .A1(n7998), .A2(net225047), .ZN(n2594) );
  INV_X4 U2637 ( .A(n6164), .ZN(n4935) );
  INV_X4 U2638 ( .A(net225047), .ZN(n2618) );
  INV_X8 U2639 ( .A(n3787), .ZN(n2595) );
  INV_X4 U2640 ( .A(n6075), .ZN(n3787) );
  INV_X16 U2641 ( .A(net230144), .ZN(n3252) );
  INV_X8 U2642 ( .A(n7117), .ZN(n7325) );
  NOR2_X1 U2643 ( .A1(n5311), .A2(net228087), .ZN(n5312) );
  INV_X2 U2644 ( .A(n5312), .ZN(n5315) );
  NAND2_X4 U2645 ( .A1(n3213), .A2(n3214), .ZN(n5185) );
  AOI21_X2 U2646 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7024) );
  AOI21_X4 U2647 ( .B1(n5306), .B2(n5305), .A(n5304), .ZN(n2607) );
  BUF_X16 U2648 ( .A(net220851), .Z(net230611) );
  NAND2_X4 U2649 ( .A1(n7106), .A2(net224861), .ZN(n3604) );
  NAND3_X2 U2651 ( .A1(n4804), .A2(n4803), .A3(net225251), .ZN(n2596) );
  AOI22_X4 U2652 ( .A1(n8096), .A2(n2713), .B1(n3643), .B2(memAddr[14]), .ZN(
        n4878) );
  NAND3_X2 U2653 ( .A1(n6917), .A2(n3254), .A3(n6914), .ZN(n2597) );
  NAND2_X4 U2654 ( .A1(n6916), .A2(n6915), .ZN(n6917) );
  INV_X4 U2656 ( .A(net229291), .ZN(net225600) );
  INV_X2 U2657 ( .A(n3866), .ZN(n2598) );
  NOR2_X1 U2658 ( .A1(n7331), .A2(n3950), .ZN(n6996) );
  OAI22_X4 U2659 ( .A1(n7539), .A2(n2623), .B1(n7680), .B2(net225243), .ZN(
        n4736) );
  INV_X2 U2660 ( .A(n5644), .ZN(n2599) );
  INV_X8 U2661 ( .A(n6678), .ZN(n5644) );
  NOR3_X4 U2662 ( .A1(n5382), .A2(n5377), .A3(net222515), .ZN(n5381) );
  INV_X4 U2663 ( .A(n6917), .ZN(n6924) );
  NAND2_X2 U2664 ( .A1(n5155), .A2(n5156), .ZN(n3461) );
  BUF_X32 U2665 ( .A(n5467), .Z(n2600) );
  NAND2_X1 U2666 ( .A1(n4930), .A2(n4856), .ZN(n4933) );
  NAND2_X1 U2667 ( .A1(n4856), .A2(n3840), .ZN(n3676) );
  NAND2_X4 U2668 ( .A1(n3527), .A2(n3526), .ZN(n5401) );
  MUX2_X2 U2669 ( .A(n5116), .B(n2923), .S(n2601), .Z(net220921) );
  INV_X32 U2670 ( .A(net224735), .ZN(n2601) );
  INV_X8 U2671 ( .A(n6466), .ZN(n5989) );
  OAI22_X2 U2673 ( .A1(n7993), .A2(net222515), .B1(n3200), .B2(n3920), .ZN(
        n5538) );
  NAND2_X1 U2674 ( .A1(n3572), .A2(n2597), .ZN(n2602) );
  NAND2_X2 U2675 ( .A1(n3572), .A2(n6907), .ZN(n7342) );
  INV_X2 U2676 ( .A(n3903), .ZN(n4924) );
  AOI22_X2 U2677 ( .A1(net223245), .A2(n2710), .B1(n4812), .B2(memAddr[23]), 
        .ZN(n4741) );
  INV_X1 U2678 ( .A(n2577), .ZN(n6408) );
  NAND3_X2 U2679 ( .A1(n4986), .A2(n4987), .A3(n3206), .ZN(n2603) );
  NAND3_X2 U2680 ( .A1(n4986), .A2(n4987), .A3(n3206), .ZN(n4990) );
  INV_X8 U2681 ( .A(n3283), .ZN(net224781) );
  NOR2_X2 U2682 ( .A1(n7986), .A2(n6755), .ZN(n6186) );
  NAND2_X4 U2683 ( .A1(n3307), .A2(n3308), .ZN(n3306) );
  INV_X4 U2684 ( .A(net223242), .ZN(n3308) );
  NAND2_X4 U2685 ( .A1(net221477), .A2(net220851), .ZN(n2604) );
  NAND2_X2 U2686 ( .A1(net221477), .A2(net220851), .ZN(net220638) );
  NAND2_X4 U2687 ( .A1(n5360), .A2(net225047), .ZN(n5361) );
  NAND2_X2 U2689 ( .A1(n5768), .A2(net224737), .ZN(n5769) );
  INV_X8 U2690 ( .A(n3290), .ZN(n2605) );
  INV_X8 U2691 ( .A(n2605), .ZN(n2606) );
  INV_X4 U2693 ( .A(net225238), .ZN(n3304) );
  NAND2_X1 U2695 ( .A1(n6058), .A2(n3212), .ZN(n3419) );
  NOR2_X4 U2696 ( .A1(n5323), .A2(n5303), .ZN(n5306) );
  XNOR2_X2 U2697 ( .A(n7974), .B(net224865), .ZN(n2608) );
  NOR3_X4 U2698 ( .A1(net225226), .A2(n3899), .A3(n2719), .ZN(n4911) );
  AOI21_X4 U2699 ( .B1(n6372), .B2(n2611), .A(n2610), .ZN(n2609) );
  INV_X4 U2700 ( .A(n2609), .ZN(n6376) );
  INV_X32 U2701 ( .A(n6375), .ZN(n2610) );
  AND2_X2 U2702 ( .A1(n6374), .A2(net221479), .ZN(n2611) );
  INV_X1 U2703 ( .A(n3785), .ZN(n2612) );
  NAND2_X2 U2704 ( .A1(net229628), .A2(net225601), .ZN(n2645) );
  INV_X2 U2705 ( .A(n2646), .ZN(net220757) );
  NOR3_X2 U2706 ( .A1(net225226), .A2(n2728), .A3(n3860), .ZN(n4903) );
  NOR2_X2 U2707 ( .A1(n3860), .A2(n2726), .ZN(n3840) );
  NAND2_X2 U2708 ( .A1(net223346), .A2(net225091), .ZN(n3860) );
  NAND2_X4 U2710 ( .A1(net221770), .A2(net221165), .ZN(n2613) );
  INV_X8 U2711 ( .A(net221432), .ZN(net221770) );
  NAND2_X2 U2712 ( .A1(net221770), .A2(net221165), .ZN(net220876) );
  NAND4_X2 U2713 ( .A1(n5031), .A2(n5028), .A3(n5030), .A4(n5029), .ZN(n2614)
         );
  INV_X8 U2714 ( .A(n5027), .ZN(n5028) );
  NOR2_X1 U2715 ( .A1(n3860), .A2(n2960), .ZN(n4908) );
  INV_X2 U2716 ( .A(net221757), .ZN(n3191) );
  NAND2_X1 U2717 ( .A1(net221757), .A2(net220651), .ZN(n3193) );
  INV_X1 U2718 ( .A(net220921), .ZN(net220310) );
  NAND2_X2 U2719 ( .A1(n5075), .A2(n5074), .ZN(n5076) );
  NAND2_X1 U2720 ( .A1(n6873), .A2(n2577), .ZN(n6413) );
  INV_X32 U2721 ( .A(net230142), .ZN(net230143) );
  OAI21_X4 U2722 ( .B1(n5607), .B2(n5606), .A(n2970), .ZN(n5608) );
  NAND2_X4 U2723 ( .A1(net223245), .A2(n2749), .ZN(n4974) );
  INV_X8 U2724 ( .A(n5593), .ZN(n5595) );
  AOI21_X4 U2726 ( .B1(n6561), .B2(n6560), .A(n3742), .ZN(n6562) );
  NAND3_X2 U2727 ( .A1(n6559), .A2(n6558), .A3(n6698), .ZN(n6560) );
  INV_X8 U2728 ( .A(n4812), .ZN(n2623) );
  INV_X2 U2729 ( .A(n6770), .ZN(n6772) );
  XOR2_X2 U2730 ( .A(net224865), .B(n7032), .Z(n6065) );
  INV_X4 U2731 ( .A(n7032), .ZN(n7027) );
  NAND3_X2 U2732 ( .A1(n6583), .A2(n5457), .A3(n5456), .ZN(n2615) );
  NOR2_X4 U2734 ( .A1(n6229), .A2(n6227), .ZN(n2617) );
  NAND2_X1 U2735 ( .A1(n5007), .A2(n2618), .ZN(n3845) );
  NAND2_X4 U2736 ( .A1(n3409), .A2(n3410), .ZN(n6404) );
  INV_X4 U2737 ( .A(net221819), .ZN(n3342) );
  AND2_X2 U2739 ( .A1(n3127), .A2(n4722), .ZN(n2619) );
  INV_X32 U2740 ( .A(n3863), .ZN(n3864) );
  INV_X2 U2741 ( .A(n6888), .ZN(n3496) );
  AOI22_X2 U2742 ( .A1(n6650), .A2(n6651), .B1(n6649), .B2(n6648), .ZN(n2620)
         );
  INV_X4 U2743 ( .A(n6168), .ZN(n3621) );
  NOR3_X4 U2744 ( .A1(n2675), .A2(n6161), .A3(n6645), .ZN(n6162) );
  NAND2_X4 U2745 ( .A1(n6586), .A2(n7297), .ZN(n2621) );
  INV_X1 U2746 ( .A(n6586), .ZN(n2622) );
  NAND2_X4 U2747 ( .A1(net230231), .A2(n7326), .ZN(n7280) );
  AOI21_X4 U2748 ( .B1(n5319), .B2(n3133), .A(net222745), .ZN(n5320) );
  INV_X2 U2749 ( .A(n5888), .ZN(n5889) );
  NOR2_X2 U2750 ( .A1(n3042), .A2(n3416), .ZN(n2675) );
  INV_X8 U2751 ( .A(n5093), .ZN(n4812) );
  AND2_X2 U2752 ( .A1(net225091), .A2(net228615), .ZN(n3248) );
  AOI211_X4 U2755 ( .C1(n4296), .C2(n4297), .A(n4295), .B(n4294), .ZN(n2625)
         );
  AOI211_X2 U2756 ( .C1(n4296), .C2(n4297), .A(n4295), .B(n4294), .ZN(n4301)
         );
  INV_X2 U2758 ( .A(n4513), .ZN(n4511) );
  INV_X2 U2761 ( .A(iAddr[26]), .ZN(n4533) );
  NAND2_X4 U2762 ( .A1(n7148), .A2(n7304), .ZN(n7149) );
  NOR2_X4 U2763 ( .A1(n7057), .A2(n3482), .ZN(n5814) );
  BUF_X4 U2764 ( .A(n6606), .Z(n3151) );
  XNOR2_X2 U2765 ( .A(n3544), .B(n5910), .ZN(n2627) );
  AOI21_X4 U2766 ( .B1(n5909), .B2(n6528), .A(n5908), .ZN(n5910) );
  NOR2_X2 U2767 ( .A1(n4865), .A2(n2787), .ZN(n4930) );
  NAND2_X1 U2768 ( .A1(n5731), .A2(n7169), .ZN(n5263) );
  BUF_X32 U2769 ( .A(n3784), .Z(n2628) );
  OAI211_X2 U2770 ( .C1(n6964), .C2(n7230), .A(n6480), .B(n6479), .ZN(n3166)
         );
  INV_X4 U2772 ( .A(n7126), .ZN(n6697) );
  BUF_X32 U2773 ( .A(net228087), .Z(n2629) );
  AND2_X2 U2774 ( .A1(n2627), .A2(n2630), .ZN(n5917) );
  INV_X32 U2775 ( .A(n3950), .ZN(n2630) );
  OAI211_X1 U2777 ( .C1(n6225), .C2(n3942), .A(n6224), .B(n6223), .ZN(n6350)
         );
  OAI211_X1 U2778 ( .C1(n4792), .C2(n3942), .A(n6210), .B(n6209), .ZN(n6783)
         );
  AOI22_X4 U2779 ( .A1(n7239), .A2(n6514), .B1(n7176), .B2(n6620), .ZN(n6515)
         );
  NAND2_X2 U2780 ( .A1(n5967), .A2(n5960), .ZN(n5240) );
  NAND2_X4 U2782 ( .A1(n6462), .A2(n6840), .ZN(n6193) );
  INV_X8 U2783 ( .A(n5409), .ZN(n4843) );
  NAND2_X4 U2785 ( .A1(n4746), .A2(n4745), .ZN(n5203) );
  NOR2_X2 U2786 ( .A1(n7684), .A2(net225243), .ZN(n4724) );
  INV_X1 U2787 ( .A(n6685), .ZN(n2631) );
  INV_X4 U2788 ( .A(n2631), .ZN(n2632) );
  BUF_X32 U2789 ( .A(n6038), .Z(n2633) );
  OAI21_X1 U2790 ( .B1(n6742), .B2(n7933), .A(n6740), .ZN(n6743) );
  NAND2_X4 U2792 ( .A1(n3517), .A2(n3257), .ZN(n3497) );
  NOR2_X2 U2793 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  AND3_X2 U2794 ( .A1(net225237), .A2(n3904), .A3(n2992), .ZN(n2634) );
  INV_X16 U2795 ( .A(n6842), .ZN(n3915) );
  NAND3_X2 U2796 ( .A1(n4815), .A2(net225237), .A3(net225045), .ZN(n5036) );
  INV_X8 U2797 ( .A(n3263), .ZN(n5120) );
  NAND2_X4 U2798 ( .A1(n5119), .A2(net224737), .ZN(n3263) );
  INV_X16 U2799 ( .A(n3902), .ZN(n3903) );
  AND3_X4 U2800 ( .A1(reg31Val_0[23]), .A2(n3898), .A3(net228359), .ZN(n2635)
         );
  INV_X8 U2801 ( .A(n5751), .ZN(n3267) );
  INV_X8 U2802 ( .A(n6721), .ZN(n3525) );
  NAND2_X2 U2803 ( .A1(n4755), .A2(n4754), .ZN(n3517) );
  INV_X8 U2805 ( .A(n6530), .ZN(n5902) );
  NAND2_X1 U2806 ( .A1(n3916), .A2(n7044), .ZN(n2636) );
  NAND2_X4 U2807 ( .A1(n3419), .A2(n3420), .ZN(n2692) );
  NAND2_X4 U2808 ( .A1(n5298), .A2(n3907), .ZN(n5605) );
  INV_X16 U2809 ( .A(n2701), .ZN(n3921) );
  NOR2_X4 U2810 ( .A1(n7260), .A2(n7259), .ZN(n7196) );
  INV_X2 U2811 ( .A(n6120), .ZN(n6121) );
  NAND2_X2 U2812 ( .A1(net220882), .A2(net225601), .ZN(n6120) );
  NAND2_X4 U2813 ( .A1(n5052), .A2(net230683), .ZN(n3378) );
  AND2_X2 U2814 ( .A1(n5777), .A2(n7997), .ZN(n2637) );
  INV_X8 U2815 ( .A(n7140), .ZN(n3652) );
  INV_X4 U2816 ( .A(n5205), .ZN(n5648) );
  NAND2_X4 U2817 ( .A1(n3461), .A2(net229596), .ZN(n3601) );
  AND2_X2 U2818 ( .A1(n7217), .A2(n7939), .ZN(n2638) );
  INV_X8 U2819 ( .A(n5972), .ZN(n3815) );
  INV_X8 U2821 ( .A(n6835), .ZN(n6836) );
  NAND3_X4 U2823 ( .A1(n5289), .A2(n3947), .A3(n5288), .ZN(n7168) );
  NAND2_X4 U2824 ( .A1(n5453), .A2(n7967), .ZN(n3473) );
  AND3_X4 U2825 ( .A1(n2924), .A2(n3297), .A3(n3298), .ZN(n2639) );
  NAND2_X4 U2826 ( .A1(n2928), .A2(net229061), .ZN(n2641) );
  INV_X4 U2827 ( .A(net229061), .ZN(n2640) );
  NOR2_X1 U2828 ( .A1(n6557), .A2(n6556), .ZN(n6559) );
  AND3_X4 U2829 ( .A1(n6936), .A2(n3722), .A3(n6935), .ZN(n6127) );
  NOR2_X4 U2830 ( .A1(net221761), .A2(n6144), .ZN(n6163) );
  NAND2_X1 U2832 ( .A1(n5205), .A2(n3272), .ZN(n2643) );
  NAND2_X2 U2833 ( .A1(n5648), .A2(n2642), .ZN(n2644) );
  NAND2_X2 U2834 ( .A1(n2644), .A2(n2643), .ZN(n5649) );
  INV_X1 U2835 ( .A(n3272), .ZN(n2642) );
  INV_X8 U2836 ( .A(net224861), .ZN(n3272) );
  NAND2_X2 U2837 ( .A1(n3092), .A2(n3450), .ZN(n3451) );
  NAND2_X4 U2838 ( .A1(net229628), .A2(net225601), .ZN(n2646) );
  INV_X1 U2839 ( .A(n6035), .ZN(n3821) );
  NAND2_X4 U2840 ( .A1(net221863), .A2(n2658), .ZN(net229736) );
  INV_X1 U2841 ( .A(n6175), .ZN(n6362) );
  INV_X1 U2842 ( .A(n5298), .ZN(n2647) );
  INV_X1 U2846 ( .A(n5071), .ZN(n4845) );
  NAND2_X2 U2847 ( .A1(net220894), .A2(n6881), .ZN(n3394) );
  NAND3_X1 U2848 ( .A1(n3904), .A2(n2651), .A3(net224749), .ZN(n2650) );
  NOR3_X4 U2849 ( .A1(n2780), .A2(n3864), .A3(net224997), .ZN(n2652) );
  INV_X4 U2850 ( .A(n2652), .ZN(n5613) );
  INV_X4 U2851 ( .A(n3824), .ZN(n6157) );
  NAND2_X4 U2852 ( .A1(n5612), .A2(n6780), .ZN(n2653) );
  NAND2_X1 U2854 ( .A1(n5611), .A2(n6965), .ZN(n3693) );
  INV_X2 U2855 ( .A(n5611), .ZN(n3691) );
  NAND2_X2 U2856 ( .A1(n3639), .A2(net228942), .ZN(n3359) );
  AOI211_X2 U2858 ( .C1(n4726), .C2(net225045), .A(n4724), .B(n4725), .ZN(
        n5153) );
  NAND2_X1 U2859 ( .A1(n2621), .A2(n3615), .ZN(n6556) );
  NOR2_X2 U2860 ( .A1(n6837), .A2(n6591), .ZN(n3241) );
  NOR2_X4 U2861 ( .A1(n4995), .A2(n4994), .ZN(n5001) );
  OAI21_X2 U2862 ( .B1(n7096), .B2(n5845), .A(n5844), .ZN(n5848) );
  INV_X8 U2863 ( .A(n6873), .ZN(n6875) );
  OAI22_X1 U2864 ( .A1(net225243), .A2(n7676), .B1(n3901), .B2(n7535), .ZN(
        n4763) );
  AND2_X2 U2865 ( .A1(net224731), .A2(net224859), .ZN(n3120) );
  INV_X8 U2866 ( .A(net221922), .ZN(net229628) );
  OAI221_X4 U2868 ( .B1(n7569), .B2(n4925), .C1(net225226), .C2(n2927), .A(
        n5358), .ZN(n5360) );
  INV_X8 U2869 ( .A(n6909), .ZN(n6373) );
  NOR2_X2 U2871 ( .A1(n5123), .A2(n3384), .ZN(n5138) );
  XNOR2_X2 U2872 ( .A(n5775), .B(net227884), .ZN(n2654) );
  NAND2_X2 U2874 ( .A1(n6500), .A2(n2655), .ZN(n2656) );
  NAND2_X1 U2875 ( .A1(n2902), .A2(net230157), .ZN(n2657) );
  NAND2_X2 U2876 ( .A1(n2656), .A2(n2657), .ZN(n5103) );
  INV_X4 U2877 ( .A(net230157), .ZN(n2655) );
  NAND2_X2 U2878 ( .A1(n5131), .A2(n5132), .ZN(n6500) );
  NAND2_X4 U2879 ( .A1(net223245), .A2(n2747), .ZN(n5004) );
  INV_X4 U2880 ( .A(n5004), .ZN(n4998) );
  INV_X4 U2881 ( .A(n5373), .ZN(n6739) );
  AND2_X2 U2882 ( .A1(n6413), .A2(net228941), .ZN(n2910) );
  INV_X8 U2884 ( .A(n3414), .ZN(n3415) );
  OAI21_X2 U2885 ( .B1(n7943), .B2(n5340), .A(n5339), .ZN(n5350) );
  INV_X4 U2886 ( .A(net228940), .ZN(net228941) );
  NAND2_X2 U2887 ( .A1(n5820), .A2(n5484), .ZN(n3364) );
  INV_X1 U2888 ( .A(net220875), .ZN(n2658) );
  NAND2_X4 U2889 ( .A1(n3368), .A2(n3369), .ZN(n6112) );
  NAND2_X4 U2890 ( .A1(net221165), .A2(n6141), .ZN(n6142) );
  INV_X8 U2891 ( .A(n5244), .ZN(n3857) );
  NAND2_X2 U2893 ( .A1(n5116), .A2(n2659), .ZN(n2660) );
  NAND2_X2 U2894 ( .A1(n2923), .A2(n3312), .ZN(n2661) );
  NAND2_X4 U2895 ( .A1(n2660), .A2(n2661), .ZN(n5117) );
  INV_X1 U2896 ( .A(n3312), .ZN(n2659) );
  NAND2_X2 U2897 ( .A1(n2859), .A2(net229656), .ZN(n2662) );
  NAND2_X2 U2898 ( .A1(n3601), .A2(n2662), .ZN(n5171) );
  NOR2_X2 U2899 ( .A1(n5171), .A2(n5045), .ZN(n3802) );
  OAI21_X4 U2900 ( .B1(n7986), .B2(n3196), .A(n3722), .ZN(n6948) );
  INV_X4 U2901 ( .A(net222840), .ZN(n3350) );
  INV_X2 U2902 ( .A(n3134), .ZN(n4431) );
  XNOR2_X1 U2903 ( .A(n7502), .B(n4433), .ZN(n4434) );
  AOI22_X4 U2904 ( .A1(n4584), .A2(n2846), .B1(n4583), .B2(n7554), .ZN(n4682)
         );
  NAND2_X4 U2905 ( .A1(n4305), .A2(n4304), .ZN(n4306) );
  NAND4_X2 U2908 ( .A1(n5788), .A2(n5789), .A3(n5790), .A4(n5791), .ZN(n2664)
         );
  NAND4_X2 U2909 ( .A1(n5788), .A2(n5789), .A3(n5791), .A4(n5790), .ZN(n7160)
         );
  OAI21_X4 U2910 ( .B1(n7154), .B2(n3950), .A(n7153), .ZN(n7159) );
  NAND3_X4 U2911 ( .A1(n4469), .A2(iAddr[12]), .A3(iAddr[11]), .ZN(n4473) );
  NOR3_X4 U2912 ( .A1(n4360), .A2(n4345), .A3(n3399), .ZN(n2665) );
  INV_X4 U2913 ( .A(n2665), .ZN(n4537) );
  INV_X1 U2914 ( .A(n4500), .ZN(n2666) );
  INV_X4 U2915 ( .A(n4491), .ZN(iAddr[19]) );
  NOR2_X1 U2916 ( .A1(n4692), .A2(n7925), .ZN(n4678) );
  NAND2_X1 U2917 ( .A1(op0_1), .A2(n7707), .ZN(n4676) );
  NOR2_X1 U2918 ( .A1(op0_1), .A2(n7707), .ZN(n4660) );
  NAND2_X1 U2919 ( .A1(n4617), .A2(n7707), .ZN(n6319) );
  NOR2_X1 U2920 ( .A1(n7707), .A2(n2849), .ZN(n4565) );
  NAND2_X4 U2921 ( .A1(n7707), .A2(n4692), .ZN(n4581) );
  AOI211_X4 U2922 ( .C1(n2664), .C2(n5825), .A(n5823), .B(n5824), .ZN(n5826)
         );
  INV_X8 U2923 ( .A(n3963), .ZN(n4389) );
  NAND2_X4 U2924 ( .A1(n3962), .A2(n2768), .ZN(n3963) );
  NOR2_X4 U2925 ( .A1(n3970), .A2(n7504), .ZN(n3134) );
  INV_X1 U2926 ( .A(n3970), .ZN(n4429) );
  BUF_X8 U2927 ( .A(n4045), .Z(n2668) );
  NAND2_X4 U2928 ( .A1(n4530), .A2(iAddr[26]), .ZN(n3687) );
  NAND2_X4 U2929 ( .A1(n4315), .A2(iAddr[26]), .ZN(n4317) );
  OAI21_X4 U2930 ( .B1(n7139), .B2(n7138), .A(n7141), .ZN(n5815) );
  XNOR2_X1 U2932 ( .A(n4362), .B(iAddr[31]), .ZN(n4552) );
  OAI21_X4 U2933 ( .B1(n3896), .B2(n4035), .A(n4034), .ZN(iAddr[31]) );
  INV_X4 U2934 ( .A(n2677), .ZN(n3502) );
  AOI22_X2 U2935 ( .A1(n6661), .A2(n6495), .B1(n5835), .B2(n3955), .ZN(n5836)
         );
  XNOR2_X2 U2936 ( .A(n4547), .B(n2669), .ZN(n4548) );
  MUX2_X2 U2938 ( .A(n4548), .B(reg31Val_0[30]), .S(net224691), .Z(n2174) );
  NAND3_X4 U2939 ( .A1(n3552), .A2(n2857), .A3(n3966), .ZN(n4404) );
  NOR2_X4 U2940 ( .A1(n7501), .A2(n4547), .ZN(n3972) );
  INV_X4 U2941 ( .A(net228615), .ZN(n2670) );
  INV_X16 U2942 ( .A(net225096), .ZN(net228615) );
  NAND2_X2 U2944 ( .A1(n6852), .A2(n3924), .ZN(n6855) );
  NAND2_X2 U2945 ( .A1(n7645), .A2(n4666), .ZN(\hazard_detect/eq_83/A[0] ) );
  INV_X1 U2946 ( .A(n4666), .ZN(n6311) );
  NAND2_X4 U2947 ( .A1(n7647), .A2(n4666), .ZN(\hazard_detect/eq_83/A[2] ) );
  NAND2_X4 U2948 ( .A1(op0_1), .A2(n4311), .ZN(n4666) );
  NAND2_X4 U2949 ( .A1(n4578), .A2(n7711), .ZN(n4592) );
  NAND3_X1 U2950 ( .A1(n4578), .A2(n2847), .A3(n2765), .ZN(n4579) );
  NOR3_X4 U2951 ( .A1(n7884), .A2(n2761), .A3(n6319), .ZN(n4578) );
  INV_X4 U2952 ( .A(n6608), .ZN(n6609) );
  INV_X4 U2953 ( .A(n4723), .ZN(n2671) );
  INV_X4 U2954 ( .A(n3158), .ZN(n6696) );
  NAND2_X1 U2955 ( .A1(n3924), .A2(n3158), .ZN(n7131) );
  INV_X1 U2956 ( .A(n5801), .ZN(n2672) );
  INV_X8 U2957 ( .A(n6570), .ZN(n3796) );
  AOI22_X2 U2958 ( .A1(n6852), .A2(n3921), .B1(n6853), .B2(n7127), .ZN(n6134)
         );
  INV_X8 U2959 ( .A(n6851), .ZN(n6100) );
  AOI211_X2 U2960 ( .C1(n6371), .C2(n6370), .A(net221487), .B(n6369), .ZN(
        n6380) );
  INV_X2 U2961 ( .A(n6058), .ZN(n5178) );
  NAND2_X2 U2962 ( .A1(n5182), .A2(n6685), .ZN(n3663) );
  OAI21_X2 U2963 ( .B1(n5180), .B2(n5181), .A(n5179), .ZN(n5182) );
  OAI22_X4 U2964 ( .A1(n6672), .A2(n6610), .B1(n6607), .B2(n2703), .ZN(n6497)
         );
  OAI22_X4 U2966 ( .A1(n2700), .A2(n4876), .B1(n3253), .B2(n4875), .ZN(n5474)
         );
  INV_X4 U2967 ( .A(net230144), .ZN(n3253) );
  INV_X1 U2968 ( .A(n5172), .ZN(n5177) );
  INV_X8 U2969 ( .A(n5098), .ZN(n5368) );
  NAND2_X4 U2970 ( .A1(n7245), .A2(n7247), .ZN(n6429) );
  INV_X8 U2971 ( .A(n6428), .ZN(n7247) );
  INV_X4 U2972 ( .A(n3847), .ZN(n3848) );
  BUF_X32 U2973 ( .A(n2596), .Z(n2673) );
  INV_X8 U2974 ( .A(n6061), .ZN(n4745) );
  NAND2_X4 U2975 ( .A1(n3969), .A2(n2771), .ZN(n3970) );
  NAND2_X4 U2976 ( .A1(n4433), .A2(n2887), .ZN(n4547) );
  BUF_X32 U2977 ( .A(n5116), .Z(n2674) );
  NAND2_X4 U2978 ( .A1(n5134), .A2(n5133), .ZN(n5194) );
  NAND3_X2 U2979 ( .A1(n5132), .A2(net224731), .A3(n5131), .ZN(n5134) );
  OAI211_X4 U2980 ( .C1(n5983), .C2(n7201), .A(n5982), .B(n7170), .ZN(n2681)
         );
  NAND3_X2 U2981 ( .A1(n6583), .A2(n5457), .A3(n5456), .ZN(n5451) );
  INV_X2 U2982 ( .A(n3300), .ZN(n7287) );
  INV_X4 U2983 ( .A(n3938), .ZN(n3944) );
  INV_X8 U2985 ( .A(n6753), .ZN(n5633) );
  NAND2_X2 U2986 ( .A1(n5309), .A2(n5310), .ZN(n4717) );
  NAND2_X4 U2987 ( .A1(n5308), .A2(n5310), .ZN(n5303) );
  AND2_X4 U2988 ( .A1(n4822), .A2(net225214), .ZN(n2676) );
  AND2_X2 U2989 ( .A1(n4822), .A2(net225214), .ZN(n3551) );
  NOR3_X4 U2990 ( .A1(n5617), .A2(n5616), .A3(n5615), .ZN(n5629) );
  NAND2_X2 U2992 ( .A1(net220851), .A2(n3205), .ZN(n7084) );
  INV_X4 U2993 ( .A(n7019), .ZN(n7007) );
  NAND2_X4 U2994 ( .A1(n5972), .A2(n2759), .ZN(n2678) );
  NAND2_X1 U2995 ( .A1(n2759), .A2(n5972), .ZN(n5716) );
  NOR2_X2 U2997 ( .A1(n2784), .A2(n3933), .ZN(n5264) );
  NOR2_X2 U2999 ( .A1(n7550), .A2(n2606), .ZN(n6088) );
  NOR2_X2 U3000 ( .A1(n7567), .A2(n3290), .ZN(n4789) );
  INV_X2 U3001 ( .A(n5216), .ZN(n5217) );
  NAND3_X2 U3002 ( .A1(n3845), .A2(n5015), .A3(n3844), .ZN(n5219) );
  NAND2_X2 U3003 ( .A1(n5015), .A2(n3510), .ZN(n5216) );
  NAND2_X1 U3004 ( .A1(n7007), .A2(n8005), .ZN(n7016) );
  INV_X4 U3005 ( .A(net221806), .ZN(net221888) );
  NAND2_X4 U3006 ( .A1(n4931), .A2(memAddr[5]), .ZN(n2679) );
  NAND2_X1 U3007 ( .A1(n4812), .A2(memAddr[5]), .ZN(n5056) );
  NOR2_X2 U3008 ( .A1(net35052), .A2(net223348), .ZN(n3335) );
  NOR2_X4 U3010 ( .A1(n4887), .A2(n3715), .ZN(n4917) );
  INV_X2 U3011 ( .A(n5458), .ZN(n5376) );
  OAI221_X2 U3012 ( .B1(n5473), .B2(n5474), .C1(n5472), .C2(n5471), .A(n5470), 
        .ZN(n2680) );
  OAI221_X2 U3013 ( .B1(n5473), .B2(n5474), .C1(n5472), .C2(n5471), .A(n5470), 
        .ZN(n5508) );
  INV_X8 U3016 ( .A(n5853), .ZN(n7227) );
  NAND2_X4 U3017 ( .A1(n4901), .A2(net224995), .ZN(n4905) );
  NAND2_X4 U3018 ( .A1(net221806), .A2(net221805), .ZN(net230730) );
  NAND2_X4 U3019 ( .A1(n7168), .A2(n7169), .ZN(n7170) );
  NOR2_X4 U3020 ( .A1(n6646), .A2(n3642), .ZN(n6649) );
  NAND2_X4 U3023 ( .A1(n6597), .A2(n6596), .ZN(n6599) );
  NAND3_X4 U3024 ( .A1(n5388), .A2(net224737), .A3(net224871), .ZN(n5389) );
  NAND4_X2 U3025 ( .A1(n7303), .A2(n3300), .A3(n7302), .A4(n7304), .ZN(n7309)
         );
  INV_X2 U3026 ( .A(n5193), .ZN(n3201) );
  NOR2_X2 U3027 ( .A1(net225230), .A2(n7550), .ZN(n3714) );
  NAND3_X2 U3028 ( .A1(n5648), .A2(n5366), .A3(n7997), .ZN(n5209) );
  NAND2_X4 U3029 ( .A1(net221799), .A2(net228495), .ZN(n3338) );
  NAND2_X1 U3030 ( .A1(n4955), .A2(n4954), .ZN(n5498) );
  INV_X32 U3032 ( .A(net225001), .ZN(net224997) );
  INV_X32 U3033 ( .A(net225003), .ZN(net225001) );
  NAND3_X2 U3034 ( .A1(n4883), .A2(n3455), .A3(net224993), .ZN(n4884) );
  NOR2_X4 U3035 ( .A1(n6165), .A2(n2580), .ZN(n6166) );
  AOI21_X4 U3036 ( .B1(n5423), .B2(net224745), .A(n5422), .ZN(n5424) );
  NOR3_X4 U3037 ( .A1(n3920), .A2(n3933), .A3(n7938), .ZN(n5422) );
  INV_X4 U3038 ( .A(n6631), .ZN(n3428) );
  NOR2_X4 U3039 ( .A1(n4715), .A2(net228359), .ZN(n2683) );
  INV_X2 U3040 ( .A(net220405), .ZN(net221791) );
  AOI21_X1 U3041 ( .B1(net225251), .B2(net223341), .A(net223342), .ZN(
        net223340) );
  NAND2_X4 U3043 ( .A1(n5540), .A2(n5551), .ZN(n6705) );
  BUF_X4 U3044 ( .A(n6249), .Z(n3542) );
  OAI22_X4 U3045 ( .A1(n7562), .A2(net225015), .B1(n2791), .B2(n2699), .ZN(
        n6249) );
  INV_X8 U3046 ( .A(n3350), .ZN(net225226) );
  NAND4_X4 U3047 ( .A1(n6133), .A2(n6132), .A3(n6130), .A4(n6131), .ZN(n6852)
         );
  INV_X8 U3049 ( .A(n4864), .ZN(n5190) );
  NAND2_X4 U3051 ( .A1(n6394), .A2(n5937), .ZN(n6192) );
  INV_X2 U3052 ( .A(n6382), .ZN(n6390) );
  NOR4_X1 U3054 ( .A1(n6296), .A2(n6295), .A3(net224957), .A4(n6294), .ZN(
        \id_ex/N41 ) );
  INV_X16 U3055 ( .A(net224753), .ZN(net224751) );
  INV_X8 U3056 ( .A(net33207), .ZN(net224753) );
  INV_X16 U3057 ( .A(net222698), .ZN(net225229) );
  INV_X8 U3058 ( .A(n5092), .ZN(n5130) );
  AOI21_X4 U3060 ( .B1(n5974), .B2(n6114), .A(n5973), .ZN(n5981) );
  NAND2_X4 U3061 ( .A1(n3722), .A2(n6935), .ZN(n3414) );
  INV_X4 U3062 ( .A(net230622), .ZN(n3455) );
  OAI21_X4 U3063 ( .B1(n7114), .B2(n7113), .A(net229482), .ZN(n7116) );
  NOR2_X4 U3064 ( .A1(n3933), .A2(n7938), .ZN(n5407) );
  NOR2_X2 U3065 ( .A1(n3936), .A2(n4757), .ZN(n5064) );
  NOR2_X2 U3066 ( .A1(net223345), .A2(net222840), .ZN(net223341) );
  OAI21_X2 U3067 ( .B1(n5093), .B2(n7525), .A(n4827), .ZN(n4828) );
  NAND3_X1 U3068 ( .A1(net228018), .A2(n7606), .A3(net228029), .ZN(n4827) );
  NAND2_X1 U3069 ( .A1(n3934), .A2(\wb/dsize_reg/z2 [16]), .ZN(n5560) );
  NAND2_X1 U3070 ( .A1(n3934), .A2(\wb/dsize_reg/z2 [21]), .ZN(n6049) );
  NAND2_X1 U3071 ( .A1(\wb/dsize_reg/z2 [14]), .A2(n3934), .ZN(n4948) );
  NAND2_X2 U3072 ( .A1(n3812), .A2(n6705), .ZN(n5542) );
  NAND3_X4 U3073 ( .A1(n4916), .A2(net224783), .A3(net225214), .ZN(n4922) );
  NOR2_X2 U3074 ( .A1(n6945), .A2(n3815), .ZN(n6949) );
  OAI22_X4 U3075 ( .A1(n5093), .A2(n7421), .B1(net225243), .B2(n7678), .ZN(
        n4910) );
  NAND2_X4 U3076 ( .A1(net223348), .A2(n2670), .ZN(n5093) );
  NAND2_X4 U3077 ( .A1(n5972), .A2(n5886), .ZN(n5214) );
  NAND2_X4 U3078 ( .A1(n4413), .A2(n3723), .ZN(n4383) );
  OAI21_X1 U3079 ( .B1(n3944), .B2(n5578), .A(n3133), .ZN(n5579) );
  INV_X4 U3080 ( .A(n4967), .ZN(n7254) );
  NAND2_X2 U3081 ( .A1(n7718), .A2(net224929), .ZN(n4967) );
  INV_X8 U3082 ( .A(n2638), .ZN(n3922) );
  OAI21_X1 U3084 ( .B1(n6207), .B2(n3940), .A(n6206), .ZN(n6356) );
  OAI21_X1 U3085 ( .B1(n5715), .B2(n3940), .A(n5714), .ZN(n6358) );
  OAI21_X1 U3086 ( .B1(n6536), .B2(n6535), .A(n6534), .ZN(n6537) );
  AOI21_X2 U3087 ( .B1(net224843), .B2(n6532), .A(net224835), .ZN(n6536) );
  OAI21_X2 U3088 ( .B1(n6735), .B2(net224851), .A(n2838), .ZN(n6738) );
  INV_X4 U3090 ( .A(net224855), .ZN(net224851) );
  NAND3_X2 U3091 ( .A1(n7254), .A2(n2704), .A3(n2756), .ZN(n3913) );
  INV_X8 U3092 ( .A(n3914), .ZN(n6661) );
  INV_X4 U3093 ( .A(n2838), .ZN(net224835) );
  NOR3_X2 U3094 ( .A1(n4192), .A2(n4188), .A3(n3895), .ZN(n4190) );
  INV_X4 U3095 ( .A(n4326), .ZN(n4524) );
  OAI21_X1 U3096 ( .B1(n5691), .B2(n3940), .A(n5690), .ZN(n6341) );
  OAI21_X2 U3097 ( .B1(n5284), .B2(n3941), .A(n5620), .ZN(n6791) );
  INV_X4 U3098 ( .A(n7182), .ZN(n7151) );
  OAI21_X1 U3099 ( .B1(n3944), .B2(n5563), .A(n3133), .ZN(n5564) );
  NAND2_X2 U3100 ( .A1(n7086), .A2(n7084), .ZN(n7090) );
  NAND2_X2 U3102 ( .A1(n5054), .A2(net224995), .ZN(n5518) );
  INV_X4 U3103 ( .A(n5243), .ZN(n5245) );
  INV_X4 U3104 ( .A(n6882), .ZN(n6147) );
  INV_X4 U3105 ( .A(n6373), .ZN(n3205) );
  INV_X4 U3106 ( .A(n5503), .ZN(n3477) );
  AOI21_X2 U3107 ( .B1(n6242), .B2(n3942), .A(net225083), .ZN(n5364) );
  NAND3_X2 U3108 ( .A1(n5362), .A2(n5361), .A3(n6242), .ZN(n5363) );
  OAI21_X2 U3109 ( .B1(n6472), .B2(n6471), .A(n3862), .ZN(n6473) );
  INV_X4 U3110 ( .A(n7097), .ZN(n3737) );
  NOR2_X2 U3111 ( .A1(n3921), .A2(n2914), .ZN(n7261) );
  NOR2_X2 U3112 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  AOI21_X2 U3113 ( .B1(n7185), .B2(n2838), .A(n7184), .ZN(n7186) );
  NAND2_X2 U3114 ( .A1(n3492), .A2(n3493), .ZN(n3606) );
  INV_X4 U3115 ( .A(n4127), .ZN(n3995) );
  NOR2_X2 U3116 ( .A1(n4023), .A2(n4024), .ZN(n3466) );
  AOI21_X2 U3117 ( .B1(n4287), .B2(n4293), .A(n4292), .ZN(n4279) );
  INV_X2 U3118 ( .A(n5653), .ZN(n5655) );
  INV_X4 U3119 ( .A(net224743), .ZN(net224733) );
  INV_X4 U3120 ( .A(n6984), .ZN(n6989) );
  NAND2_X2 U3121 ( .A1(net221798), .A2(net229037), .ZN(net220319) );
  INV_X4 U3122 ( .A(net220601), .ZN(net229481) );
  INV_X4 U3123 ( .A(n4117), .ZN(n4110) );
  OAI21_X2 U3125 ( .B1(n4210), .B2(n4318), .A(n4209), .ZN(n4211) );
  NOR2_X2 U3126 ( .A1(n7670), .A2(net224897), .ZN(n4203) );
  NAND2_X2 U3127 ( .A1(net220320), .A2(n3338), .ZN(net220405) );
  AOI21_X1 U3128 ( .B1(n6759), .B2(n2838), .A(n7201), .ZN(n6760) );
  NOR2_X1 U3129 ( .A1(n6756), .A2(n6755), .ZN(n6762) );
  AOI21_X1 U3130 ( .B1(net224843), .B2(n7201), .A(net224835), .ZN(n6756) );
  NOR3_X2 U3131 ( .A1(n4665), .A2(n2761), .A3(n2870), .ZN(n4591) );
  NAND3_X2 U3132 ( .A1(n2724), .A2(n4566), .A3(n4565), .ZN(n4657) );
  NOR2_X2 U3133 ( .A1(net225238), .A2(n2916), .ZN(n4916) );
  AOI21_X2 U3134 ( .B1(n3944), .B2(n7351), .A(n5226), .ZN(n5227) );
  AOI21_X2 U3136 ( .B1(net224843), .B2(n3876), .A(net224835), .ZN(n6177) );
  INV_X4 U3137 ( .A(n5635), .ZN(n5636) );
  OAI21_X1 U3138 ( .B1(n6235), .B2(n3940), .A(n6234), .ZN(n6334) );
  NOR2_X2 U3139 ( .A1(n2849), .A2(n4572), .ZN(n4617) );
  AOI21_X2 U3140 ( .B1(net224843), .B2(n6505), .A(net224835), .ZN(n6503) );
  NOR2_X2 U3141 ( .A1(n6565), .A2(n2840), .ZN(n6566) );
  NOR2_X2 U3142 ( .A1(net224833), .A2(n6564), .ZN(n6571) );
  NOR2_X2 U3143 ( .A1(net224833), .A2(n6716), .ZN(n6722) );
  NOR2_X2 U3145 ( .A1(n6717), .A2(n2840), .ZN(n6718) );
  NOR2_X2 U3146 ( .A1(n6736), .A2(n2840), .ZN(n6737) );
  OAI211_X2 U3147 ( .C1(n5101), .C2(n5445), .A(n5100), .B(net224737), .ZN(
        n5102) );
  NAND3_X2 U3148 ( .A1(n7254), .A2(n2704), .A3(n2756), .ZN(n7182) );
  NOR2_X2 U3149 ( .A1(net220307), .A2(n3011), .ZN(n3317) );
  NOR2_X2 U3150 ( .A1(n3318), .A2(n3319), .ZN(net220298) );
  NOR2_X2 U3151 ( .A1(setInv_2), .A2(n2841), .ZN(n3319) );
  NOR2_X2 U3153 ( .A1(n6236), .A2(n3075), .ZN(n6053) );
  NOR2_X2 U3154 ( .A1(n4168), .A2(n3896), .ZN(n4169) );
  NOR2_X1 U3155 ( .A1(n7418), .A2(n4465), .ZN(n4191) );
  NAND2_X2 U3156 ( .A1(n4029), .A2(n4266), .ZN(n4270) );
  NOR2_X2 U3157 ( .A1(n7630), .A2(net224909), .ZN(n4033) );
  NAND3_X2 U3158 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n6333) );
  NOR2_X2 U3159 ( .A1(n4374), .A2(n4373), .ZN(n4380) );
  NOR3_X2 U3160 ( .A1(n4377), .A2(n4376), .A3(n4375), .ZN(n4378) );
  NAND3_X2 U3161 ( .A1(n6267), .A2(n2856), .A3(n6266), .ZN(n6268) );
  NOR2_X2 U3162 ( .A1(rd_3[3]), .A2(rd_3[2]), .ZN(n6267) );
  NOR2_X2 U3163 ( .A1(rd_3[1]), .A2(rd_3[4]), .ZN(n6266) );
  INV_X4 U3164 ( .A(n3961), .ZN(n4385) );
  OAI21_X1 U3165 ( .B1(n7434), .B2(n4465), .A(n4460), .ZN(n4561) );
  OAI21_X1 U3166 ( .B1(n7435), .B2(n4465), .A(n4464), .ZN(n4563) );
  OAI21_X2 U3167 ( .B1(n4444), .B2(n4448), .A(n4443), .ZN(n4445) );
  AOI21_X2 U3168 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4559) );
  NOR2_X2 U3169 ( .A1(n4571), .A2(n4570), .ZN(n4687) );
  NOR2_X1 U3170 ( .A1(net224955), .A2(n4672), .ZN(n4570) );
  INV_X4 U3171 ( .A(n4657), .ZN(n4658) );
  NAND3_X2 U3172 ( .A1(n4604), .A2(n7556), .A3(n4569), .ZN(n4672) );
  NOR2_X2 U3173 ( .A1(net33230), .A2(n7711), .ZN(n4569) );
  INV_X4 U3174 ( .A(n4593), .ZN(n4583) );
  NOR2_X2 U3175 ( .A1(n4581), .A2(n7925), .ZN(n4584) );
  NOR2_X1 U3176 ( .A1(net224933), .A2(n2848), .ZN(net223657) );
  NAND3_X2 U3177 ( .A1(net33230), .A2(n7711), .A3(n7556), .ZN(n4603) );
  INV_X4 U3178 ( .A(n4496), .ZN(n3147) );
  INV_X4 U3179 ( .A(n5149), .ZN(n4755) );
  AOI22_X2 U3180 ( .A1(n6608), .A2(n7239), .B1(n6495), .B2(n7176), .ZN(n5729)
         );
  NOR2_X2 U3181 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  OAI21_X2 U3182 ( .B1(n6018), .B2(n6017), .A(n6016), .ZN(n6019) );
  NOR2_X2 U3183 ( .A1(n6100), .A2(n3918), .ZN(n6025) );
  NAND3_X2 U3184 ( .A1(n5689), .A2(n5688), .A3(n5687), .ZN(n6340) );
  AOI21_X2 U3185 ( .B1(n5686), .B2(n3945), .A(n6070), .ZN(n5687) );
  OAI21_X1 U3186 ( .B1(n5700), .B2(n3940), .A(n5699), .ZN(n6533) );
  NOR3_X2 U3187 ( .A1(n6273), .A2(n6272), .A3(n3008), .ZN(n6274) );
  NOR2_X2 U3188 ( .A1(n6331), .A2(n6308), .ZN(n6314) );
  NOR2_X1 U3189 ( .A1(n6312), .A2(net224955), .ZN(n6313) );
  NOR2_X2 U3190 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  NOR2_X2 U3191 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  NOR2_X2 U3192 ( .A1(n6670), .A2(n2703), .ZN(n6674) );
  NOR2_X1 U3193 ( .A1(n6774), .A2(n6965), .ZN(n6775) );
  OAI21_X2 U3194 ( .B1(n6772), .B2(net224851), .A(n2838), .ZN(n6773) );
  OAI21_X2 U3195 ( .B1(n6794), .B2(n6793), .A(n6792), .ZN(n6795) );
  AOI21_X2 U3196 ( .B1(n3725), .B2(net224843), .A(net224835), .ZN(n6794) );
  NOR2_X2 U3198 ( .A1(n7124), .A2(n2840), .ZN(n7125) );
  NOR2_X2 U3199 ( .A1(net224833), .A2(n7105), .ZN(n7111) );
  NAND4_X2 U3200 ( .A1(n5865), .A2(n5867), .A3(n5866), .A4(n5868), .ZN(n3158)
         );
  NAND3_X1 U3201 ( .A1(n4797), .A2(n5575), .A3(n5580), .ZN(regWrData[3]) );
  NAND3_X2 U3202 ( .A1(n4808), .A2(n2798), .A3(n4807), .ZN(regWrData[6]) );
  AOI21_X1 U3203 ( .B1(net225011), .B2(n2966), .A(n4801), .ZN(n4808) );
  NOR2_X2 U3204 ( .A1(n4806), .A2(n4805), .ZN(n4807) );
  NOR2_X2 U3205 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  NOR2_X1 U3206 ( .A1(n7413), .A2(n4465), .ZN(n4063) );
  NOR2_X1 U3207 ( .A1(n4164), .A2(n4171), .ZN(n4040) );
  NOR2_X2 U3209 ( .A1(net225015), .A2(n7973), .ZN(n5408) );
  OAI21_X1 U3210 ( .B1(n3944), .B2(n5476), .A(n5634), .ZN(n5479) );
  NOR2_X1 U3211 ( .A1(n3942), .A2(net225084), .ZN(n5397) );
  NAND2_X2 U3212 ( .A1(n3187), .A2(n3188), .ZN(n3190) );
  INV_X4 U3214 ( .A(n5631), .ZN(n3755) );
  NOR2_X2 U3215 ( .A1(n5525), .A2(n5524), .ZN(n5532) );
  NAND2_X2 U3216 ( .A1(n6400), .A2(n5522), .ZN(n5521) );
  OAI22_X2 U3217 ( .A1(n3933), .A2(n5385), .B1(net222672), .B2(net224737), 
        .ZN(n5392) );
  OAI21_X2 U3218 ( .B1(net225083), .B2(n5636), .A(net224859), .ZN(n5637) );
  INV_X4 U3219 ( .A(n5009), .ZN(n5010) );
  INV_X4 U3220 ( .A(n6064), .ZN(n3654) );
  INV_X4 U3221 ( .A(n5564), .ZN(n3287) );
  NAND2_X2 U3222 ( .A1(n3499), .A2(n2588), .ZN(n5210) );
  NOR2_X2 U3223 ( .A1(n4047), .A2(n4000), .ZN(n4001) );
  NAND2_X2 U3224 ( .A1(net223245), .A2(n2742), .ZN(n5414) );
  BUF_X4 U3225 ( .A(n3294), .Z(n3629) );
  NAND3_X1 U3226 ( .A1(n5523), .A2(net224731), .A3(n5518), .ZN(n5062) );
  NOR3_X2 U3227 ( .A1(n3242), .A2(regWrData[26]), .A3(n6070), .ZN(n6078) );
  NAND2_X2 U3228 ( .A1(n7730), .A2(net228407), .ZN(n3633) );
  NOR2_X1 U3229 ( .A1(n7242), .A2(n6502), .ZN(n5938) );
  INV_X4 U3230 ( .A(n3697), .ZN(n3698) );
  INV_X8 U3231 ( .A(n6486), .ZN(n5455) );
  NOR2_X1 U3232 ( .A1(n7242), .A2(n5675), .ZN(n5676) );
  NAND4_X2 U3233 ( .A1(n5245), .A2(n6216), .A3(n6214), .A4(n6212), .ZN(n5247)
         );
  NAND2_X2 U3234 ( .A1(n5014), .A2(n2995), .ZN(n3793) );
  NAND2_X2 U3236 ( .A1(\wb/dsize_reg/z2 [28]), .A2(net224993), .ZN(n3468) );
  INV_X4 U3237 ( .A(n3427), .ZN(n3426) );
  NOR2_X2 U3238 ( .A1(n3725), .A2(n3862), .ZN(n6442) );
  INV_X4 U3239 ( .A(zeroExt_2), .ZN(net225082) );
  NAND2_X2 U3240 ( .A1(n5989), .A2(n6114), .ZN(n3706) );
  NAND2_X2 U3241 ( .A1(n4754), .A2(n4755), .ZN(n6048) );
  NAND2_X2 U3242 ( .A1(net228809), .A2(n3352), .ZN(net220769) );
  NOR2_X2 U3244 ( .A1(net220838), .A2(n6910), .ZN(n6887) );
  NAND2_X2 U3245 ( .A1(n7243), .A2(n7242), .ZN(n7246) );
  NAND2_X2 U3246 ( .A1(n7203), .A2(n6430), .ZN(n6425) );
  NOR2_X2 U3247 ( .A1(n7205), .A2(n3952), .ZN(n7206) );
  NAND2_X2 U3248 ( .A1(n7110), .A2(net229579), .ZN(n3605) );
  NAND2_X2 U3249 ( .A1(n3992), .A2(n4119), .ZN(n4072) );
  NOR2_X2 U3251 ( .A1(n4082), .A2(n4151), .ZN(n3985) );
  NAND4_X2 U3252 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4530)
         );
  NAND3_X2 U3253 ( .A1(n4524), .A2(n4521), .A3(n4520), .ZN(n4528) );
  NAND3_X2 U3254 ( .A1(n4524), .A2(n4523), .A3(n4522), .ZN(n4527) );
  OAI21_X2 U3255 ( .B1(n7473), .B2(n3974), .A(n7472), .ZN(net221340) );
  NAND2_X2 U3256 ( .A1(n2608), .A2(n3197), .ZN(n3199) );
  NOR2_X1 U3258 ( .A1(n7242), .A2(n5940), .ZN(n5941) );
  NOR2_X2 U3259 ( .A1(n3522), .A2(n6551), .ZN(n6554) );
  NOR2_X1 U3260 ( .A1(n6594), .A2(n6588), .ZN(n6589) );
  NOR2_X2 U3262 ( .A1(n3522), .A2(n6701), .ZN(n6703) );
  INV_X4 U3263 ( .A(n6700), .ZN(n6711) );
  NOR2_X2 U3264 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  NAND2_X2 U3265 ( .A1(n3389), .A2(n3502), .ZN(n3504) );
  NAND3_X2 U3266 ( .A1(n6989), .A2(n6988), .A3(net220757), .ZN(n6990) );
  NAND2_X2 U3267 ( .A1(n7141), .A2(n7143), .ZN(n7136) );
  NAND3_X2 U3268 ( .A1(n7263), .A2(n7262), .A3(n7261), .ZN(n7264) );
  NOR2_X1 U3269 ( .A1(n2914), .A2(n7255), .ZN(n7258) );
  OAI21_X2 U3270 ( .B1(n3995), .B2(n3994), .A(n4131), .ZN(n3224) );
  NOR2_X2 U3271 ( .A1(n7457), .A2(n7510), .ZN(n4020) );
  OAI21_X2 U3272 ( .B1(n4279), .B2(n4280), .A(n4026), .ZN(n4027) );
  NAND2_X2 U3273 ( .A1(n6376), .A2(net230488), .ZN(n3800) );
  NAND3_X2 U3274 ( .A1(n4364), .A2(n2850), .A3(n4363), .ZN(n4365) );
  NOR2_X2 U3275 ( .A1(rd_2[3]), .A2(rd_2[4]), .ZN(n4364) );
  NOR2_X2 U3276 ( .A1(rd_2[0]), .A2(rd_2[1]), .ZN(n4363) );
  NAND3_X2 U3277 ( .A1(n4582), .A2(n6303), .A3(n2720), .ZN(n4593) );
  INV_X4 U3278 ( .A(n4472), .ZN(n4469) );
  NOR2_X1 U3279 ( .A1(n7324), .A2(n3950), .ZN(n5849) );
  NOR2_X2 U3280 ( .A1(n5829), .A2(n2840), .ZN(n5830) );
  NAND3_X1 U3281 ( .A1(n3944), .A2(net225013), .A3(n2925), .ZN(n5266) );
  NOR2_X2 U3282 ( .A1(n7620), .A2(n7617), .ZN(n6269) );
  NAND3_X2 U3283 ( .A1(n7626), .A2(n7625), .A3(n7627), .ZN(n6272) );
  NOR3_X2 U3284 ( .A1(net221424), .A2(net221425), .A3(net221426), .ZN(
        net221411) );
  NAND2_X2 U3285 ( .A1(n6661), .A2(n5864), .ZN(n5748) );
  NOR2_X2 U3286 ( .A1(n6190), .A2(n5973), .ZN(n6198) );
  OAI21_X2 U3287 ( .B1(n6488), .B2(n3285), .A(n2615), .ZN(n6826) );
  NOR2_X2 U3288 ( .A1(n6588), .A2(n6593), .ZN(n6488) );
  INV_X8 U3289 ( .A(n7205), .ZN(n3955) );
  NOR2_X2 U3290 ( .A1(net220314), .A2(net220537), .ZN(net220536) );
  NOR2_X1 U3291 ( .A1(n6236), .A2(n3076), .ZN(n5561) );
  INV_X4 U3292 ( .A(n4683), .ZN(n4311) );
  NOR2_X1 U3293 ( .A1(n4110), .A2(n4109), .ZN(n4112) );
  INV_X4 U3294 ( .A(n4045), .ZN(n4105) );
  NOR2_X2 U3295 ( .A1(n7672), .A2(net224909), .ZN(n4064) );
  NOR3_X2 U3296 ( .A1(n4238), .A2(n4250), .A3(n3681), .ZN(n4215) );
  AOI21_X2 U3297 ( .B1(n3897), .B2(n2993), .A(n4203), .ZN(n4204) );
  NOR2_X2 U3298 ( .A1(n4249), .A2(n4201), .ZN(n4206) );
  AOI21_X2 U3300 ( .B1(net221791), .B2(n7275), .A(n3950), .ZN(n6122) );
  NOR2_X2 U3301 ( .A1(n6094), .A2(n2840), .ZN(n6095) );
  NOR2_X2 U3302 ( .A1(n6632), .A2(n6791), .ZN(n6345) );
  NOR2_X1 U3303 ( .A1(n6341), .A2(n6340), .ZN(n6347) );
  NOR2_X1 U3304 ( .A1(n6358), .A2(n6357), .ZN(n6361) );
  NOR2_X1 U3305 ( .A1(n6334), .A2(n7046), .ZN(n6337) );
  NOR2_X2 U3306 ( .A1(n6422), .A2(n6783), .ZN(n6354) );
  NAND2_X2 U3307 ( .A1(n6728), .A2(n3921), .ZN(n6378) );
  NOR3_X2 U3308 ( .A1(n6762), .A2(n6761), .A3(n6760), .ZN(n6763) );
  NOR2_X2 U3309 ( .A1(n6757), .A2(n2840), .ZN(n6761) );
  INV_X4 U3310 ( .A(n4581), .ZN(n4595) );
  NOR2_X2 U3311 ( .A1(n2846), .A2(n4674), .ZN(n4596) );
  AOI21_X2 U3312 ( .B1(n2788), .B2(n2720), .A(n4599), .ZN(n4600) );
  NOR2_X2 U3313 ( .A1(n2846), .A2(n4663), .ZN(n4597) );
  INV_X4 U3314 ( .A(net224749), .ZN(net224747) );
  INV_X4 U3315 ( .A(n4404), .ZN(n3163) );
  INV_X4 U3316 ( .A(n3959), .ZN(n4413) );
  NAND2_X2 U3317 ( .A1(n3958), .A2(n2921), .ZN(n3959) );
  INV_X4 U3318 ( .A(n4411), .ZN(n3958) );
  INV_X4 U3319 ( .A(net224693), .ZN(net224683) );
  INV_X4 U3320 ( .A(n3971), .ZN(n4433) );
  NAND2_X2 U3321 ( .A1(n3134), .A2(n2769), .ZN(n3971) );
  INV_X4 U3322 ( .A(\mem_wb/N41 ), .ZN(net224719) );
  INV_X4 U3323 ( .A(\mem_wb/N41 ), .ZN(net224725) );
  INV_X4 U3324 ( .A(\mem_wb/N41 ), .ZN(net224723) );
  INV_X4 U3325 ( .A(\mem_wb/N41 ), .ZN(net224721) );
  OAI21_X2 U3326 ( .B1(n4549), .B2(n6271), .A(net224919), .ZN(net221531) );
  INV_X4 U3327 ( .A(\mem_wb/N41 ), .ZN(net224693) );
  NOR2_X2 U3328 ( .A1(n4616), .A2(n4615), .ZN(n4619) );
  AOI21_X2 U3329 ( .B1(n2772), .B2(n4670), .A(n7554), .ZN(n4618) );
  NAND2_X2 U3330 ( .A1(n4604), .A2(n7378), .ZN(n4665) );
  NAND2_X2 U3331 ( .A1(n2911), .A2(n4595), .ZN(n4683) );
  NAND3_X2 U3332 ( .A1(net224933), .A2(n4690), .A3(n4605), .ZN(n4691) );
  NAND2_X2 U3333 ( .A1(n4538), .A2(n4540), .ZN(n4539) );
  NOR2_X2 U3334 ( .A1(n3240), .A2(n4511), .ZN(n4698) );
  NOR2_X2 U3335 ( .A1(n3238), .A2(n3239), .ZN(n3240) );
  INV_X4 U3336 ( .A(n3928), .ZN(n3930) );
  NOR3_X2 U3337 ( .A1(n3899), .A2(n3290), .A3(n7576), .ZN(n4732) );
  NAND2_X2 U3338 ( .A1(n5111), .A2(n5112), .ZN(n5071) );
  NOR2_X2 U3339 ( .A1(n4969), .A2(n2840), .ZN(n4970) );
  OAI21_X1 U3340 ( .B1(n5753), .B2(n5776), .A(n5752), .ZN(n5754) );
  NOR2_X1 U3341 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  AOI21_X1 U3342 ( .B1(net224843), .B2(n5820), .A(net224835), .ZN(n5822) );
  NOR2_X2 U3343 ( .A1(net221856), .A2(n6081), .ZN(n6082) );
  OAI21_X1 U3344 ( .B1(net221858), .B2(n6080), .A(n6079), .ZN(n6081) );
  NOR2_X2 U3345 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  AOI21_X1 U3346 ( .B1(n6173), .B2(n2838), .A(n3876), .ZN(n6179) );
  OAI21_X1 U3347 ( .B1(n6177), .B2(n6188), .A(n6176), .ZN(n6178) );
  NAND2_X2 U3348 ( .A1(net224933), .A2(n2858), .ZN(n4668) );
  NOR2_X2 U3349 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  NOR2_X2 U3350 ( .A1(n6503), .A2(n6502), .ZN(n6508) );
  AOI21_X1 U3351 ( .B1(n6506), .B2(n2838), .A(n6505), .ZN(n6507) );
  NOR2_X2 U3352 ( .A1(n7718), .A2(n6512), .ZN(n6513) );
  INV_X4 U3353 ( .A(n6537), .ZN(n3153) );
  AOI21_X2 U3354 ( .B1(n3951), .B2(n6573), .A(n6572), .ZN(n6574) );
  AOI21_X1 U3355 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(n6569) );
  NOR2_X2 U3356 ( .A1(n6580), .A2(n2840), .ZN(n6581) );
  OAI21_X1 U3357 ( .B1(n6584), .B2(net224851), .A(n2838), .ZN(n6582) );
  AOI21_X2 U3358 ( .B1(n3951), .B2(n7287), .A(n6723), .ZN(n6724) );
  AOI21_X1 U3359 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6740) );
  NOR2_X2 U3360 ( .A1(net224833), .A2(n6734), .ZN(n6742) );
  NOR2_X1 U3361 ( .A1(n7295), .A2(n3950), .ZN(n6849) );
  OAI21_X1 U3362 ( .B1(n6846), .B2(n6845), .A(n6844), .ZN(n6847) );
  AOI21_X1 U3363 ( .B1(net224843), .B2(n3916), .A(net224833), .ZN(n6846) );
  AOI21_X1 U3364 ( .B1(n6841), .B2(n2838), .A(n3916), .ZN(n6848) );
  NOR2_X1 U3365 ( .A1(net220310), .A2(n2838), .ZN(n6862) );
  NOR2_X2 U3366 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  NOR2_X2 U3367 ( .A1(n7051), .A2(n7050), .ZN(n7052) );
  OAI21_X1 U3368 ( .B1(n7049), .B2(n7048), .A(n7047), .ZN(n7050) );
  NOR2_X2 U3369 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  AOI21_X2 U3370 ( .B1(net224843), .B2(n7155), .A(net224835), .ZN(n7157) );
  NAND3_X2 U3371 ( .A1(n6241), .A2(n6240), .A3(n6239), .ZN(regWrData[9]) );
  NAND2_X2 U3372 ( .A1(n4960), .A2(n4959), .ZN(regWrData[11]) );
  NAND3_X1 U3373 ( .A1(net224991), .A2(n5356), .A3(\wb/dsize_reg/z2 [30]), 
        .ZN(n4949) );
  NAND3_X2 U3374 ( .A1(n4962), .A2(n6049), .A3(n6051), .ZN(regWrData[21]) );
  OAI21_X2 U3375 ( .B1(n7641), .B2(net224909), .A(n4564), .ZN(iAddr[0]) );
  OAI21_X2 U3376 ( .B1(n7640), .B2(net224909), .A(n4562), .ZN(iAddr[1]) );
  OAI211_X2 U3377 ( .C1(n4125), .C2(n3895), .A(n4124), .B(n4123), .ZN(iAddr[3]) );
  NAND3_X2 U3378 ( .A1(n4097), .A2(n4096), .A3(n4095), .ZN(iAddr[5]) );
  NAND3_X2 U3379 ( .A1(n4092), .A2(n4091), .A3(n2962), .ZN(iAddr[7]) );
  OAI211_X2 U3380 ( .C1(n4134), .C2(n3159), .A(n4524), .B(n3171), .ZN(n4136)
         );
  NAND3_X2 U3381 ( .A1(n4176), .A2(n4175), .A3(n4174), .ZN(iAddr[17]) );
  AOI21_X2 U3382 ( .B1(n2942), .B2(n4192), .A(n4191), .ZN(n4194) );
  NOR2_X2 U3383 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  NOR2_X2 U3384 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  NOR2_X2 U3385 ( .A1(n7468), .A2(n4465), .ZN(n4032) );
  NAND3_X2 U3386 ( .A1(n2855), .A2(n4684), .A3(n2757), .ZN(n4688) );
  NOR2_X2 U3387 ( .A1(net33197), .A2(net224897), .ZN(\ex_mem/N150 ) );
  NOR2_X2 U3388 ( .A1(n7720), .A2(net224899), .ZN(\ex_mem/N133 ) );
  NOR2_X2 U3389 ( .A1(n7739), .A2(net224897), .ZN(\ex_mem/N151 ) );
  NOR2_X2 U3390 ( .A1(n7749), .A2(net224899), .ZN(\ex_mem/N132 ) );
  NOR2_X2 U3391 ( .A1(net224909), .A2(n2945), .ZN(\ex_mem/N237 ) );
  NOR2_X2 U3392 ( .A1(n7658), .A2(net224893), .ZN(\ex_mem/N57 ) );
  NOR2_X2 U3393 ( .A1(n7742), .A2(net224897), .ZN(\ex_mem/N147 ) );
  NOR2_X2 U3394 ( .A1(n7748), .A2(net224899), .ZN(\ex_mem/N134 ) );
  NOR2_X2 U3395 ( .A1(n7631), .A2(net224903), .ZN(\ex_mem/N40 ) );
  NOR2_X2 U3396 ( .A1(n7660), .A2(net224893), .ZN(\ex_mem/N55 ) );
  NOR2_X2 U3397 ( .A1(n7664), .A2(net224895), .ZN(\ex_mem/N51 ) );
  NOR2_X2 U3398 ( .A1(n7669), .A2(net224899), .ZN(\ex_mem/N45 ) );
  NOR2_X2 U3399 ( .A1(n7741), .A2(net224897), .ZN(\ex_mem/N148 ) );
  NOR2_X2 U3400 ( .A1(n7661), .A2(net224895), .ZN(\ex_mem/N54 ) );
  NOR2_X2 U3401 ( .A1(n7740), .A2(net224897), .ZN(\ex_mem/N149 ) );
  NOR2_X2 U3402 ( .A1(n7637), .A2(net224901), .ZN(\ex_mem/N39 ) );
  NOR2_X2 U3403 ( .A1(n7714), .A2(net224899), .ZN(\ex_mem/N36 ) );
  NOR2_X2 U3404 ( .A1(n7746), .A2(net224899), .ZN(\ex_mem/N137 ) );
  NOR2_X2 U3405 ( .A1(n7636), .A2(net224901), .ZN(\ex_mem/N41 ) );
  NOR2_X2 U3406 ( .A1(n7635), .A2(net224901), .ZN(\ex_mem/N42 ) );
  NOR2_X2 U3407 ( .A1(n7634), .A2(net224901), .ZN(\ex_mem/N43 ) );
  NOR3_X2 U3408 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n6284) );
  NOR2_X2 U3409 ( .A1(n6280), .A2(n6279), .ZN(n6285) );
  OAI21_X2 U3410 ( .B1(n7640), .B2(n2789), .A(n4461), .ZN(n1986) );
  OAI21_X2 U3411 ( .B1(n7641), .B2(n2789), .A(n4466), .ZN(n1990) );
  NAND3_X2 U3412 ( .A1(n2919), .A2(net224933), .A3(n2772), .ZN(\id_ex/N45 ) );
  INV_X4 U3413 ( .A(net224693), .ZN(net224681) );
  NOR2_X2 U3414 ( .A1(n2702), .A2(n4568), .ZN(n4577) );
  NOR2_X2 U3415 ( .A1(n4574), .A2(n2788), .ZN(n4575) );
  OAI21_X2 U3416 ( .B1(n7717), .B2(net224933), .A(n6315), .ZN(n7882) );
  NAND3_X2 U3417 ( .A1(n7712), .A2(n6303), .A3(n4673), .ZN(n4680) );
  AOI21_X2 U3418 ( .B1(n4678), .B2(n4677), .A(net223657), .ZN(n4679) );
  NOR2_X2 U3419 ( .A1(n7554), .A2(n4672), .ZN(n4673) );
  NOR2_X2 U3420 ( .A1(n4721), .A2(net224893), .ZN(\ex_mem/N106 ) );
  NOR2_X2 U3421 ( .A1(n4728), .A2(net224909), .ZN(\ex_mem/N115 ) );
  NOR2_X2 U3422 ( .A1(n4756), .A2(net224903), .ZN(\ex_mem/N123 ) );
  NOR2_X2 U3423 ( .A1(n4767), .A2(net224895), .ZN(\ex_mem/N130 ) );
  NOR2_X2 U3424 ( .A1(n4771), .A2(net224903), .ZN(\ex_mem/N103 ) );
  NOR2_X2 U3425 ( .A1(n4788), .A2(net224903), .ZN(\ex_mem/N101 ) );
  NOR2_X2 U3426 ( .A1(n4795), .A2(net224903), .ZN(\ex_mem/N100 ) );
  AOI211_X1 U3427 ( .C1(n4924), .C2(regWrData[1]), .A(n4794), .B(n4793), .ZN(
        n4795) );
  AOI21_X1 U3428 ( .B1(n7919), .B2(regWrData[3]), .A(n2639), .ZN(n4799) );
  AOI21_X1 U3429 ( .B1(n7919), .B2(regWrData[6]), .A(n4809), .ZN(n4810) );
  NOR2_X2 U3430 ( .A1(n4833), .A2(net224891), .ZN(\ex_mem/N107 ) );
  OAI21_X2 U3431 ( .B1(n4839), .B2(n2975), .A(net224913), .ZN(n4840) );
  NOR2_X2 U3432 ( .A1(n4855), .A2(net224903), .ZN(\ex_mem/N109 ) );
  NOR2_X2 U3433 ( .A1(n7629), .A2(net224893), .ZN(\ex_mem/N66 ) );
  NOR2_X1 U3434 ( .A1(n6390), .A2(net224903), .ZN(\ex_mem/N129 ) );
  NOR2_X2 U3435 ( .A1(net223337), .A2(net224891), .ZN(\ex_mem/N118 ) );
  NOR2_X2 U3436 ( .A1(net223329), .A2(net224903), .ZN(n2552) );
  NOR2_X2 U3437 ( .A1(n4874), .A2(net224893), .ZN(\ex_mem/N104 ) );
  NOR2_X2 U3438 ( .A1(n3533), .A2(net224903), .ZN(\ex_mem/N114 ) );
  NOR2_X2 U3439 ( .A1(n4895), .A2(net224891), .ZN(\ex_mem/N116 ) );
  AOI21_X1 U3440 ( .B1(n5019), .B2(n5773), .A(net224909), .ZN(\ex_mem/N117 )
         );
  NOR2_X2 U3441 ( .A1(n4907), .A2(net224895), .ZN(\ex_mem/N119 ) );
  NOR2_X2 U3442 ( .A1(n4915), .A2(net224903), .ZN(\ex_mem/N125 ) );
  NOR2_X2 U3443 ( .A1(n4923), .A2(net224893), .ZN(\ex_mem/N126 ) );
  NOR2_X2 U3444 ( .A1(n3547), .A2(net224903), .ZN(\ex_mem/N127 ) );
  NOR2_X2 U3445 ( .A1(n4969), .A2(net224903), .ZN(n2537) );
  NOR2_X2 U3446 ( .A1(n5744), .A2(net224903), .ZN(n2532) );
  NOR2_X2 U3447 ( .A1(n5787), .A2(net224903), .ZN(n2547) );
  NOR2_X2 U3448 ( .A1(n5829), .A2(net224903), .ZN(n2555) );
  NOR2_X2 U3449 ( .A1(n5885), .A2(net224903), .ZN(n2538) );
  NAND2_X2 U3450 ( .A1(n3924), .A2(n7918), .ZN(n5921) );
  NOR2_X2 U3451 ( .A1(n5924), .A2(net224903), .ZN(n2548) );
  NOR2_X2 U3452 ( .A1(n7124), .A2(net224903), .ZN(n2528) );
  NOR2_X2 U3453 ( .A1(n5925), .A2(net224903), .ZN(n2540) );
  NOR2_X2 U3454 ( .A1(n5926), .A2(net224903), .ZN(n2545) );
  NOR2_X2 U3455 ( .A1(net224909), .A2(n3376), .ZN(n2550) );
  NOR2_X2 U3456 ( .A1(n6351), .A2(net224903), .ZN(n2541) );
  NOR2_X2 U3457 ( .A1(n5928), .A2(net224903), .ZN(n2536) );
  OAI21_X2 U3458 ( .B1(n6022), .B2(n3950), .A(n6021), .ZN(n6023) );
  NOR2_X2 U3459 ( .A1(n6027), .A2(net224903), .ZN(n2535) );
  NOR2_X2 U3460 ( .A1(n6094), .A2(net224901), .ZN(n2556) );
  INV_X4 U3461 ( .A(net224711), .ZN(net224637) );
  NOR2_X2 U3462 ( .A1(n6362), .A2(net224901), .ZN(n2559) );
  NOR2_X2 U3463 ( .A1(n7632), .A2(net224901), .ZN(\ex_mem/N47 ) );
  NOR2_X2 U3464 ( .A1(n6205), .A2(net224901), .ZN(n2557) );
  NOR2_X2 U3465 ( .A1(n6757), .A2(net224901), .ZN(n2558) );
  NOR2_X2 U3466 ( .A1(n6208), .A2(net224901), .ZN(n2534) );
  NOR2_X2 U3467 ( .A1(n6211), .A2(net224899), .ZN(n7846) );
  NOR2_X2 U3468 ( .A1(n6222), .A2(net224899), .ZN(n7845) );
  NOR2_X2 U3469 ( .A1(n7733), .A2(net224899), .ZN(\ex_mem/N131 ) );
  NOR2_X2 U3470 ( .A1(n7721), .A2(net224899), .ZN(\ex_mem/N135 ) );
  NOR2_X2 U3471 ( .A1(n7747), .A2(net224899), .ZN(\ex_mem/N136 ) );
  NOR2_X2 U3472 ( .A1(n7745), .A2(net224899), .ZN(\ex_mem/N138 ) );
  NOR2_X2 U3473 ( .A1(n7744), .A2(net224897), .ZN(\ex_mem/N139 ) );
  NOR2_X2 U3474 ( .A1(n7725), .A2(net224897), .ZN(\ex_mem/N143 ) );
  NOR2_X2 U3475 ( .A1(n7722), .A2(net224897), .ZN(\ex_mem/N144 ) );
  NOR2_X2 U3476 ( .A1(n7726), .A2(net224897), .ZN(\ex_mem/N145 ) );
  NOR2_X2 U3477 ( .A1(n7727), .A2(net224897), .ZN(\ex_mem/N146 ) );
  NOR2_X2 U3478 ( .A1(n7738), .A2(net224895), .ZN(\ex_mem/N152 ) );
  NOR2_X2 U3479 ( .A1(n7737), .A2(net224895), .ZN(\ex_mem/N153 ) );
  NOR2_X2 U3480 ( .A1(n7736), .A2(net224895), .ZN(\ex_mem/N154 ) );
  NOR2_X2 U3481 ( .A1(n7735), .A2(net224895), .ZN(\ex_mem/N155 ) );
  NOR2_X2 U3482 ( .A1(n7734), .A2(net224895), .ZN(\ex_mem/N156 ) );
  NOR2_X2 U3483 ( .A1(n7729), .A2(net224895), .ZN(\ex_mem/N157 ) );
  NOR2_X2 U3484 ( .A1(n7728), .A2(net224895), .ZN(\ex_mem/N158 ) );
  NOR2_X2 U3485 ( .A1(n7731), .A2(net224895), .ZN(\ex_mem/N159 ) );
  NOR2_X2 U3486 ( .A1(n7732), .A2(net224895), .ZN(\ex_mem/N160 ) );
  NOR2_X2 U3487 ( .A1(n7730), .A2(net224895), .ZN(\ex_mem/N161 ) );
  NOR2_X2 U3488 ( .A1(n7723), .A2(net224895), .ZN(\ex_mem/N162 ) );
  NOR2_X2 U3489 ( .A1(n6736), .A2(net224895), .ZN(n2542) );
  NOR2_X2 U3490 ( .A1(n6226), .A2(net224895), .ZN(n2551) );
  NOR2_X2 U3491 ( .A1(n6580), .A2(net224893), .ZN(n2546) );
  NOR2_X2 U3492 ( .A1(n6244), .A2(net224893), .ZN(n2539) );
  NOR2_X2 U3493 ( .A1(n6717), .A2(net224893), .ZN(n2554) );
  NOR2_X2 U3494 ( .A1(n6565), .A2(net224893), .ZN(n2553) );
  NOR2_X2 U3495 ( .A1(n6248), .A2(net224893), .ZN(n2531) );
  NOR2_X2 U3496 ( .A1(n6256), .A2(net224893), .ZN(n2533) );
  NOR2_X2 U3497 ( .A1(n6263), .A2(net224893), .ZN(n2544) );
  INV_X4 U3498 ( .A(net224711), .ZN(net224631) );
  NOR2_X2 U3499 ( .A1(n6264), .A2(net224893), .ZN(n2530) );
  NOR2_X2 U3500 ( .A1(n7470), .A2(net224893), .ZN(\ex_mem/N240 ) );
  AOI21_X2 U3501 ( .B1(n7471), .B2(n6277), .A(net224957), .ZN(n7875) );
  NOR2_X2 U3502 ( .A1(n7717), .A2(net224893), .ZN(\ex_mem/N229 ) );
  NOR2_X2 U3503 ( .A1(n7495), .A2(net224893), .ZN(\ex_mem/N230 ) );
  NOR2_X2 U3504 ( .A1(n7479), .A2(net224893), .ZN(\ex_mem/N231 ) );
  NOR2_X2 U3505 ( .A1(n7643), .A2(net224893), .ZN(\ex_mem/N233 ) );
  NOR2_X2 U3506 ( .A1(n7644), .A2(net224891), .ZN(\ex_mem/N234 ) );
  INV_X4 U3507 ( .A(net224713), .ZN(net224639) );
  NOR2_X2 U3508 ( .A1(n7716), .A2(net224891), .ZN(\ex_mem/N235 ) );
  NOR2_X2 U3509 ( .A1(n7642), .A2(net224891), .ZN(\ex_mem/N236 ) );
  NOR2_X2 U3510 ( .A1(n7477), .A2(net224891), .ZN(\ex_mem/N239 ) );
  NOR2_X2 U3511 ( .A1(net224955), .A2(n6297), .ZN(\id_ex/N42 ) );
  INV_X4 U3512 ( .A(net224727), .ZN(net224657) );
  NOR2_X2 U3513 ( .A1(net224909), .A2(n2946), .ZN(\ex_mem/N241 ) );
  NOR2_X2 U3514 ( .A1(net224909), .A2(n2854), .ZN(\ex_mem/N246 ) );
  NOR2_X2 U3515 ( .A1(net224909), .A2(n2852), .ZN(\ex_mem/N247 ) );
  NOR2_X2 U3516 ( .A1(n6299), .A2(net224891), .ZN(\ex_mem/N99 ) );
  INV_X4 U3517 ( .A(net224713), .ZN(net224633) );
  AOI21_X2 U3518 ( .B1(n6314), .B2(n2911), .A(n6313), .ZN(n6318) );
  NOR2_X2 U3519 ( .A1(n2757), .A2(n6316), .ZN(n6317) );
  NOR2_X2 U3520 ( .A1(net224909), .A2(n2853), .ZN(\ex_mem/N243 ) );
  INV_X4 U3521 ( .A(net224711), .ZN(net224659) );
  NOR2_X2 U3523 ( .A1(net224955), .A2(n2909), .ZN(n7369) );
  NOR2_X2 U3524 ( .A1(net224955), .A2(n2907), .ZN(n7370) );
  NOR2_X2 U3525 ( .A1(net224955), .A2(n2908), .ZN(n7371) );
  NOR2_X2 U3526 ( .A1(net224955), .A2(n2904), .ZN(n7372) );
  INV_X4 U3527 ( .A(n4668), .ZN(n7379) );
  NOR2_X2 U3528 ( .A1(net224909), .A2(n2850), .ZN(\ex_mem/N245 ) );
  NOR2_X2 U3529 ( .A1(net224909), .A2(n2851), .ZN(\ex_mem/N244 ) );
  INV_X4 U3530 ( .A(net224727), .ZN(net224615) );
  NOR2_X2 U3531 ( .A1(n7650), .A2(net224891), .ZN(\ex_mem/N65 ) );
  NOR2_X2 U3532 ( .A1(n7651), .A2(net224891), .ZN(\ex_mem/N64 ) );
  NOR2_X2 U3533 ( .A1(n7652), .A2(net224891), .ZN(\ex_mem/N63 ) );
  NOR2_X2 U3534 ( .A1(n7653), .A2(net224891), .ZN(\ex_mem/N62 ) );
  NOR2_X2 U3535 ( .A1(n7654), .A2(net224891), .ZN(\ex_mem/N61 ) );
  NOR2_X2 U3536 ( .A1(n7655), .A2(net224891), .ZN(\ex_mem/N60 ) );
  NOR2_X2 U3537 ( .A1(n7656), .A2(net224891), .ZN(\ex_mem/N59 ) );
  NOR2_X2 U3538 ( .A1(n7659), .A2(net224893), .ZN(\ex_mem/N56 ) );
  NOR2_X2 U3539 ( .A1(n7666), .A2(net224895), .ZN(\ex_mem/N49 ) );
  NOR2_X2 U3540 ( .A1(n7667), .A2(net224893), .ZN(\ex_mem/N48 ) );
  INV_X4 U3541 ( .A(net224713), .ZN(net224619) );
  OAI21_X1 U3542 ( .B1(n7305), .B2(n3950), .A(n6692), .ZN(n6693) );
  NOR2_X2 U3543 ( .A1(n6776), .A2(n6775), .ZN(n6787) );
  NOR2_X2 U3544 ( .A1(n6782), .A2(n6781), .ZN(n6786) );
  AOI21_X2 U3545 ( .B1(n6797), .B2(n3649), .A(n6795), .ZN(n6808) );
  NOR3_X2 U3546 ( .A1(n7119), .A2(n7120), .A3(n7121), .ZN(n7132) );
  XNOR2_X2 U3549 ( .A(n4495), .B(n3147), .ZN(n2685) );
  XNOR2_X1 U3550 ( .A(n7928), .B(n3147), .ZN(n4701) );
  INV_X8 U3552 ( .A(n8109), .ZN(n4470) );
  XNOR2_X2 U3553 ( .A(n4513), .B(iAddr[25]), .ZN(n2686) );
  NAND2_X2 U3554 ( .A1(n4516), .A2(n4518), .ZN(n4517) );
  NAND4_X2 U3557 ( .A1(n4423), .A2(n4415), .A3(n3957), .A4(n3956), .ZN(n4411)
         );
  NAND4_X2 U3559 ( .A1(n4544), .A2(n4543), .A3(iAddr[29]), .A4(iAddr[23]), 
        .ZN(n4545) );
  NAND3_X4 U3561 ( .A1(n4436), .A2(n4437), .A3(n4435), .ZN(n4340) );
  OAI221_X2 U3562 ( .B1(n7423), .B2(n4465), .C1(n4301), .C2(n4300), .A(n4299), 
        .ZN(iAddr[28]) );
  OAI221_X2 U3563 ( .B1(n7423), .B2(n4465), .C1(n2625), .C2(n4300), .A(n4299), 
        .ZN(n7907) );
  BUF_X16 U3564 ( .A(n4153), .Z(n3438) );
  INV_X1 U3565 ( .A(n4046), .ZN(n2688) );
  INV_X4 U3566 ( .A(n2688), .ZN(n2689) );
  NAND2_X1 U3567 ( .A1(n3928), .A2(n4693), .ZN(n3619) );
  MUX2_X2 U3568 ( .A(n4552), .B(n2985), .S(n3927), .Z(n1918) );
  INV_X1 U3570 ( .A(n4037), .ZN(n4164) );
  NAND2_X4 U3571 ( .A1(n7446), .A2(n7520), .ZN(n4148) );
  OAI211_X2 U3572 ( .C1(n3374), .C2(n7139), .A(n3652), .B(n7137), .ZN(n7148)
         );
  AOI21_X2 U3573 ( .B1(n7916), .B2(n4144), .A(n4001), .ZN(n4002) );
  INV_X8 U3574 ( .A(n4139), .ZN(n3987) );
  NAND4_X4 U3575 ( .A1(n5294), .A2(n5295), .A3(n5293), .A4(n5292), .ZN(n2690)
         );
  AOI21_X2 U3576 ( .B1(n4335), .B2(n2920), .A(n4334), .ZN(n4336) );
  NOR2_X4 U3577 ( .A1(n7446), .A2(n7520), .ZN(n4334) );
  OAI211_X4 U3578 ( .C1(n4067), .C2(n4334), .A(n4337), .B(n4148), .ZN(n2691)
         );
  OAI211_X2 U3579 ( .C1(n4067), .C2(n4334), .A(n4337), .B(n4148), .ZN(n4153)
         );
  BUF_X16 U3580 ( .A(n7859), .Z(iAddr[25]) );
  NAND2_X2 U3581 ( .A1(n3141), .A2(n7447), .ZN(n3980) );
  INV_X1 U3582 ( .A(n7922), .ZN(n2693) );
  INV_X4 U3583 ( .A(n2692), .ZN(n7073) );
  NAND2_X4 U3584 ( .A1(n5085), .A2(n5086), .ZN(n5091) );
  NOR2_X4 U3585 ( .A1(n3267), .A2(n2692), .ZN(n5144) );
  AOI21_X1 U3586 ( .B1(n7072), .B2(n2838), .A(n2693), .ZN(n7078) );
  AOI21_X1 U3587 ( .B1(net224843), .B2(n2693), .A(net224833), .ZN(n7076) );
  NOR2_X4 U3588 ( .A1(net228697), .A2(n4846), .ZN(n4803) );
  BUF_X32 U3589 ( .A(n3525), .Z(n2694) );
  NAND2_X4 U3590 ( .A1(n7239), .A2(n5864), .ZN(n5292) );
  NAND2_X2 U3591 ( .A1(n6730), .A2(n6729), .ZN(\ex_mem/N207 ) );
  NAND2_X2 U3593 ( .A1(n6578), .A2(n6577), .ZN(\ex_mem/N208 ) );
  NOR3_X4 U3594 ( .A1(n2606), .A2(net230622), .A3(n7564), .ZN(n4814) );
  INV_X8 U3595 ( .A(n3248), .ZN(net230622) );
  NOR3_X4 U3598 ( .A1(n6497), .A2(n6499), .A3(n6498), .ZN(n3260) );
  NOR2_X2 U3599 ( .A1(n7026), .A2(n2701), .ZN(n6746) );
  NOR3_X4 U3600 ( .A1(n6613), .A2(n6612), .A3(n6611), .ZN(n2695) );
  NOR3_X2 U3601 ( .A1(n7069), .A2(n7068), .A3(n7067), .ZN(n7070) );
  NAND2_X2 U3602 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  OAI21_X2 U3604 ( .B1(n3260), .B2(n2701), .A(n6821), .ZN(n6833) );
  INV_X4 U3605 ( .A(net224787), .ZN(net228359) );
  OAI211_X4 U3606 ( .C1(n6939), .C2(n3862), .A(n5859), .B(n5969), .ZN(n2696)
         );
  NAND3_X4 U3607 ( .A1(n4813), .A2(n4881), .A3(net225045), .ZN(n3407) );
  INV_X8 U3609 ( .A(n3856), .ZN(n3751) );
  NAND2_X2 U3610 ( .A1(n3924), .A2(n7128), .ZN(n6518) );
  NAND3_X4 U3611 ( .A1(n6515), .A2(n6517), .A3(n6516), .ZN(n7128) );
  NAND2_X2 U3612 ( .A1(n7128), .A2(n3921), .ZN(n7129) );
  NAND2_X2 U3613 ( .A1(n5994), .A2(n5993), .ZN(n6662) );
  INV_X8 U3614 ( .A(n5914), .ZN(n3440) );
  INV_X1 U3615 ( .A(n5914), .ZN(n5886) );
  OAI21_X1 U3616 ( .B1(n5915), .B2(n5914), .A(n5913), .ZN(n5916) );
  NOR2_X1 U3617 ( .A1(net225102), .A2(n3867), .ZN(n2697) );
  NAND2_X2 U3619 ( .A1(n3805), .A2(n6380), .ZN(\ex_mem/N215 ) );
  NAND2_X4 U3620 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  INV_X4 U3621 ( .A(n5150), .ZN(n4754) );
  NOR2_X1 U3622 ( .A1(n7541), .A2(n3901), .ZN(n4725) );
  AOI21_X2 U3623 ( .B1(n6004), .B2(n5967), .A(n5708), .ZN(n5719) );
  NOR2_X2 U3624 ( .A1(n6510), .A2(n6511), .ZN(n6520) );
  INV_X8 U3625 ( .A(n3865), .ZN(n2698) );
  INV_X16 U3626 ( .A(n2698), .ZN(n2699) );
  NOR3_X4 U3627 ( .A1(n2606), .A2(n3903), .A3(n7573), .ZN(n4748) );
  NOR2_X2 U3628 ( .A1(net228280), .A2(n2947), .ZN(n4953) );
  NAND2_X4 U3629 ( .A1(net230143), .A2(net224783), .ZN(n2700) );
  INV_X16 U3630 ( .A(n3937), .ZN(n3935) );
  INV_X8 U3631 ( .A(n3937), .ZN(n3936) );
  INV_X8 U3632 ( .A(n6236), .ZN(n3937) );
  NAND2_X4 U3633 ( .A1(n3128), .A2(n3511), .ZN(n6951) );
  INV_X16 U3634 ( .A(net221157), .ZN(net229330) );
  NAND3_X4 U3635 ( .A1(net221431), .A2(net230097), .A3(n6902), .ZN(net221157)
         );
  INV_X1 U3636 ( .A(n5809), .ZN(n5812) );
  OAI21_X2 U3638 ( .B1(n6980), .B2(n3954), .A(n6979), .ZN(n6998) );
  NAND2_X4 U3639 ( .A1(n4905), .A2(n4906), .ZN(n3576) );
  NAND2_X4 U3640 ( .A1(n5572), .A2(n5618), .ZN(n5573) );
  AOI22_X4 U3641 ( .A1(n7065), .A2(n7064), .B1(n7063), .B2(n7062), .ZN(n7066)
         );
  NOR2_X2 U3642 ( .A1(n4865), .A2(n2950), .ZN(n4900) );
  OAI21_X1 U3643 ( .B1(n6980), .B2(n3918), .A(n6744), .ZN(n6745) );
  OAI22_X2 U3644 ( .A1(n6100), .A2(n3954), .B1(n6980), .B2(n3923), .ZN(n6084)
         );
  INV_X2 U3646 ( .A(n7688), .ZN(n7605) );
  OAI22_X4 U3648 ( .A1(n3935), .A2(n3083), .B1(n7558), .B2(n3253), .ZN(n5396)
         );
  INV_X4 U3649 ( .A(n3590), .ZN(n3373) );
  INV_X8 U3650 ( .A(n6824), .ZN(n5462) );
  NAND2_X4 U3651 ( .A1(n3195), .A2(n7295), .ZN(n7298) );
  OAI221_X1 U3652 ( .B1(n7306), .B2(n3950), .C1(n3260), .C2(n3918), .A(n6509), 
        .ZN(n6510) );
  NOR3_X2 U3653 ( .A1(n7290), .A2(n2794), .A3(n7291), .ZN(n7294) );
  NOR3_X2 U3654 ( .A1(n4865), .A2(n7557), .A3(n4925), .ZN(n4861) );
  INV_X8 U3655 ( .A(n3899), .ZN(n3412) );
  INV_X1 U3656 ( .A(net228495), .ZN(net229037) );
  BUF_X4 U3657 ( .A(net221770), .Z(net228495) );
  NAND2_X4 U3658 ( .A1(n5399), .A2(n5500), .ZN(n5400) );
  INV_X4 U3659 ( .A(n5541), .ZN(n3658) );
  INV_X4 U3660 ( .A(net224865), .ZN(n3242) );
  INV_X2 U3661 ( .A(net224865), .ZN(net228715) );
  INV_X4 U3662 ( .A(net224703), .ZN(net224635) );
  INV_X4 U3663 ( .A(net224703), .ZN(net224641) );
  INV_X4 U3664 ( .A(net224703), .ZN(net224653) );
  INV_X4 U3665 ( .A(net224699), .ZN(net224655) );
  INV_X4 U3666 ( .A(net224699), .ZN(net224661) );
  INV_X4 U3667 ( .A(net224699), .ZN(net224663) );
  INV_X4 U3668 ( .A(\mem_wb/N41 ), .ZN(net224699) );
  OR2_X4 U3669 ( .A1(n3566), .A2(n5658), .ZN(n2701) );
  INV_X1 U3670 ( .A(net224735), .ZN(net230157) );
  INV_X4 U3671 ( .A(\mem_wb/N41 ), .ZN(net224703) );
  INV_X4 U3672 ( .A(net224713), .ZN(net224643) );
  INV_X4 U3673 ( .A(net224711), .ZN(net224645) );
  INV_X4 U3674 ( .A(net224919), .ZN(net224891) );
  INV_X1 U3675 ( .A(net224735), .ZN(net229656) );
  INV_X4 U3676 ( .A(net224919), .ZN(net224893) );
  INV_X4 U3677 ( .A(net224915), .ZN(net224903) );
  INV_X4 U3678 ( .A(net224919), .ZN(net224895) );
  INV_X8 U3679 ( .A(n2703), .ZN(n7239) );
  INV_X8 U3680 ( .A(net224967), .ZN(net224953) );
  INV_X1 U3681 ( .A(net224735), .ZN(net229061) );
  INV_X4 U3682 ( .A(net224711), .ZN(net224673) );
  INV_X4 U3683 ( .A(net224711), .ZN(net224675) );
  AND2_X4 U3684 ( .A1(n4658), .A2(net224947), .ZN(n2702) );
  INV_X8 U3685 ( .A(net224965), .ZN(net224939) );
  INV_X16 U3686 ( .A(net224965), .ZN(net224937) );
  NAND2_X4 U3687 ( .A1(n7230), .A2(n3649), .ZN(n2703) );
  INV_X16 U3688 ( .A(net224873), .ZN(net224871) );
  INV_X1 U3689 ( .A(net224735), .ZN(n3312) );
  INV_X4 U3690 ( .A(n7192), .ZN(n3917) );
  INV_X8 U3691 ( .A(net225082), .ZN(net225084) );
  INV_X4 U3692 ( .A(net224711), .ZN(net224669) );
  INV_X4 U3693 ( .A(net224711), .ZN(net224671) );
  BUF_X4 U3694 ( .A(net33204), .Z(net225622) );
  INV_X8 U3695 ( .A(n6672), .ZN(n7176) );
  NAND3_X1 U3696 ( .A1(net225622), .A2(n7254), .A3(n2786), .ZN(n2706) );
  INV_X4 U3697 ( .A(net224953), .ZN(net224947) );
  INV_X16 U3698 ( .A(net224953), .ZN(net224933) );
  INV_X4 U3699 ( .A(n2838), .ZN(net224833) );
  INV_X4 U3700 ( .A(net221340), .ZN(net224929) );
  INV_X1 U3701 ( .A(net224735), .ZN(net228909) );
  INV_X4 U3702 ( .A(net224711), .ZN(net224625) );
  INV_X4 U3703 ( .A(net224713), .ZN(net224617) );
  INV_X4 U3704 ( .A(net224713), .ZN(net224621) );
  INV_X4 U3705 ( .A(n2840), .ZN(n7358) );
  AND2_X4 U3706 ( .A1(n7713), .A2(n2868), .ZN(n2724) );
  INV_X4 U3707 ( .A(n3951), .ZN(n3950) );
  XOR2_X2 U3708 ( .A(n7461), .B(n7506), .Z(n2725) );
  INV_X4 U3709 ( .A(net224855), .ZN(net224849) );
  INV_X4 U3710 ( .A(net220517), .ZN(net224855) );
  INV_X4 U3711 ( .A(net221531), .ZN(net224967) );
  XOR2_X2 U3712 ( .A(n2856), .B(rd_2[0]), .Z(n2738) );
  NOR3_X2 U3713 ( .A1(n4549), .A2(net224891), .A3(n6271), .ZN(n4711) );
  INV_X4 U3714 ( .A(n3928), .ZN(n3931) );
  INV_X4 U3715 ( .A(n3928), .ZN(n3932) );
  XOR2_X2 U3716 ( .A(iAddr[3]), .B(iAddr[2]), .Z(n2739) );
  AND2_X4 U3717 ( .A1(net224913), .A2(net224685), .ZN(n2740) );
  INV_X4 U3718 ( .A(net224925), .ZN(net224913) );
  INV_X4 U3719 ( .A(net224915), .ZN(net224901) );
  INV_X16 U3720 ( .A(n3917), .ZN(n3918) );
  INV_X2 U3721 ( .A(n3918), .ZN(n7127) );
  INV_X1 U3722 ( .A(net224735), .ZN(net230088) );
  INV_X4 U3723 ( .A(\mem_wb/N41 ), .ZN(net224717) );
  INV_X4 U3724 ( .A(net224711), .ZN(net224627) );
  INV_X4 U3725 ( .A(net224711), .ZN(net224629) );
  INV_X4 U3726 ( .A(net224713), .ZN(net224623) );
  INV_X4 U3727 ( .A(n2653), .ZN(n5646) );
  AND2_X4 U3728 ( .A1(n7719), .A2(net225605), .ZN(n2756) );
  AND3_X4 U3729 ( .A1(net224933), .A2(n7708), .A3(n2724), .ZN(n2757) );
  AND2_X4 U3730 ( .A1(n6358), .A2(n3133), .ZN(n2759) );
  AND2_X4 U3731 ( .A1(n6309), .A2(n4683), .ZN(n2772) );
  AND2_X4 U3732 ( .A1(n4591), .A2(n7555), .ZN(n2788) );
  AND2_X4 U3733 ( .A1(n3925), .A2(net224903), .ZN(n2789) );
  INV_X4 U3734 ( .A(net224849), .ZN(net224843) );
  AND2_X4 U3735 ( .A1(n7230), .A2(n3725), .ZN(n2790) );
  XOR2_X2 U3736 ( .A(n6799), .B(n3754), .Z(n2794) );
  AND2_X4 U3737 ( .A1(net224933), .A2(n2849), .ZN(n2795) );
  INV_X4 U3738 ( .A(net224967), .ZN(net224965) );
  AND2_X4 U3739 ( .A1(n7475), .A2(n2758), .ZN(n2796) );
  AND2_X4 U3740 ( .A1(n2723), .A2(n2758), .ZN(n2797) );
  INV_X4 U3741 ( .A(n4326), .ZN(n3894) );
  NAND2_X2 U3742 ( .A1(n7474), .A2(net224925), .ZN(n4326) );
  INV_X8 U3743 ( .A(n3894), .ZN(n3895) );
  OR2_X4 U3744 ( .A1(n3933), .A2(n3010), .ZN(n2798) );
  XOR2_X2 U3745 ( .A(n6599), .B(n3535), .Z(n2823) );
  AND2_X4 U3746 ( .A1(net224937), .A2(n2963), .ZN(n2835) );
  AND3_X4 U3747 ( .A1(n7497), .A2(n7492), .A3(n7498), .ZN(n2836) );
  NAND3_X4 U3748 ( .A1(n2756), .A2(n7254), .A3(n4968), .ZN(n2838) );
  INV_X1 U3749 ( .A(n3321), .ZN(net225605) );
  INV_X4 U3750 ( .A(net224929), .ZN(net224925) );
  INV_X4 U3751 ( .A(net224925), .ZN(net224915) );
  INV_X4 U3752 ( .A(net224925), .ZN(net224919) );
  NAND2_X2 U3753 ( .A1(net224913), .A2(n2767), .ZN(n2840) );
  INV_X8 U3754 ( .A(net225015), .ZN(net225011) );
  INV_X4 U3755 ( .A(n4711), .ZN(n3928) );
  INV_X16 U3756 ( .A(net224751), .ZN(net224741) );
  INV_X4 U3757 ( .A(\mem_wb/N41 ), .ZN(net224727) );
  INV_X4 U3758 ( .A(\mem_wb/N41 ), .ZN(net224713) );
  INV_X4 U3759 ( .A(\mem_wb/N41 ), .ZN(net224711) );
  INV_X1 U3760 ( .A(n6568), .ZN(n3261) );
  INV_X4 U3761 ( .A(n7081), .ZN(n3653) );
  XOR2_X2 U3762 ( .A(n5643), .B(n5642), .Z(n2842) );
  INV_X4 U3763 ( .A(n3867), .ZN(n4722) );
  INV_X4 U3764 ( .A(n5468), .ZN(n5467) );
  INV_X4 U3765 ( .A(n3296), .ZN(net220663) );
  INV_X8 U3766 ( .A(n4248), .ZN(n4346) );
  AND2_X4 U3767 ( .A1(n3162), .A2(n3163), .ZN(n2863) );
  INV_X4 U3768 ( .A(net222155), .ZN(net230199) );
  INV_X4 U3769 ( .A(n3868), .ZN(n3622) );
  AND2_X4 U3770 ( .A1(n7710), .A2(n7708), .ZN(n2911) );
  AND2_X4 U3771 ( .A1(n6552), .A2(n6699), .ZN(n2912) );
  AND3_X4 U3772 ( .A1(n7254), .A2(n2786), .A3(n2704), .ZN(n2914) );
  AND3_X4 U3773 ( .A1(n4615), .A2(n4550), .A3(n4572), .ZN(n2919) );
  XOR2_X1 U3774 ( .A(n7446), .B(n7520), .Z(n2920) );
  OAI22_X2 U3775 ( .A1(n7536), .A2(n3752), .B1(n7679), .B2(net225243), .ZN(
        n5063) );
  INV_X2 U3776 ( .A(n7675), .ZN(n7607) );
  AND2_X4 U3777 ( .A1(rs1[3]), .A2(net224947), .ZN(n2926) );
  AND2_X4 U3778 ( .A1(net220601), .A2(n6121), .ZN(n2929) );
  AND2_X2 U3779 ( .A1(n5996), .A2(n5997), .ZN(n2940) );
  AND2_X2 U3780 ( .A1(n4524), .A2(n4188), .ZN(n2942) );
  OR2_X4 U3781 ( .A1(net224733), .A2(n7720), .ZN(n2943) );
  INV_X4 U3782 ( .A(n2796), .ZN(net224767) );
  INV_X4 U3783 ( .A(n2796), .ZN(net224765) );
  AND3_X4 U3784 ( .A1(n4582), .A2(n7712), .A3(n2765), .ZN(n2944) );
  INV_X1 U3785 ( .A(n6861), .ZN(n6264) );
  INV_X4 U3786 ( .A(n2797), .ZN(net224759) );
  INV_X4 U3787 ( .A(n2797), .ZN(net224755) );
  INV_X4 U3788 ( .A(n7123), .ZN(n3923) );
  INV_X4 U3789 ( .A(n3923), .ZN(n3924) );
  NOR2_X2 U3790 ( .A1(n3566), .A2(n5730), .ZN(n7123) );
  OR2_X4 U3791 ( .A1(n7416), .A2(n4465), .ZN(n2961) );
  OR2_X4 U3792 ( .A1(n7467), .A2(n4465), .ZN(n2962) );
  INV_X4 U3793 ( .A(net224913), .ZN(net224909) );
  INV_X4 U3794 ( .A(net224915), .ZN(net224897) );
  INV_X4 U3795 ( .A(net224919), .ZN(net224899) );
  OR2_X4 U3796 ( .A1(net224733), .A2(n7733), .ZN(n2970) );
  OR2_X4 U3798 ( .A1(n3167), .A2(n3839), .ZN(n2975) );
  AND3_X4 U3799 ( .A1(n5438), .A2(n2596), .A3(n5436), .ZN(n2978) );
  INV_X4 U3800 ( .A(n3269), .ZN(net221881) );
  AND2_X4 U3801 ( .A1(n4416), .A2(n2741), .ZN(n2980) );
  NAND2_X1 U3802 ( .A1(n4394), .A2(n4013), .ZN(n2986) );
  AND3_X4 U3803 ( .A1(n5498), .A2(n3133), .A3(n3945), .ZN(n2989) );
  INV_X1 U3804 ( .A(n7445), .ZN(n3583) );
  OR2_X4 U3805 ( .A1(n7465), .A2(n7502), .ZN(n2994) );
  INV_X4 U3806 ( .A(n3709), .ZN(n3716) );
  AND2_X2 U3807 ( .A1(\wb/dsize_reg/z2 [26]), .A2(net224735), .ZN(n2995) );
  INV_X4 U3808 ( .A(n2591), .ZN(n3765) );
  OR2_X4 U3809 ( .A1(n6271), .A2(n2922), .ZN(n3008) );
  AND2_X4 U3810 ( .A1(net220310), .A2(n2841), .ZN(n3011) );
  INV_X4 U3811 ( .A(n3953), .ZN(n3952) );
  INV_X4 U3812 ( .A(n3953), .ZN(n3954) );
  AND3_X2 U3813 ( .A1(n5741), .A2(n5742), .A3(n5743), .ZN(n3041) );
  NAND4_X1 U3814 ( .A1(n3814), .A2(n3846), .A3(n6895), .A4(n6884), .ZN(n3042)
         );
  INV_X4 U3815 ( .A(n7674), .ZN(n7606) );
  AND3_X4 U3817 ( .A1(n7719), .A2(n7254), .A3(n2839), .ZN(n3069) );
  INV_X4 U3818 ( .A(n3530), .ZN(n3531) );
  AND2_X4 U3819 ( .A1(net224937), .A2(n2952), .ZN(n3071) );
  AND2_X4 U3820 ( .A1(net224937), .A2(n2953), .ZN(n3072) );
  AND2_X4 U3821 ( .A1(net224937), .A2(n2954), .ZN(n3073) );
  AND2_X4 U3822 ( .A1(net224937), .A2(n2968), .ZN(n3074) );
  INV_X4 U3823 ( .A(net36084), .ZN(net224777) );
  INV_X4 U3824 ( .A(net224777), .ZN(net224773) );
  OR2_X4 U3825 ( .A1(n3952), .A2(n3914), .ZN(n3088) );
  OR2_X4 U3826 ( .A1(reg31Val_3[0]), .A2(n4462), .ZN(n3091) );
  OR3_X2 U3827 ( .A1(net230741), .A2(n3864), .A3(n4982), .ZN(n3092) );
  AND2_X2 U3828 ( .A1(n4008), .A2(n4007), .ZN(n3094) );
  AND2_X4 U3829 ( .A1(n6319), .A2(n4683), .ZN(n3095) );
  OR2_X4 U3830 ( .A1(instr_2[5]), .A2(n7495), .ZN(n3117) );
  AND2_X4 U3831 ( .A1(n7378), .A2(n7554), .ZN(n3119) );
  INV_X1 U3832 ( .A(n5441), .ZN(n4805) );
  AND2_X4 U3833 ( .A1(n6629), .A2(n6628), .ZN(n3123) );
  AND2_X2 U3834 ( .A1(n6658), .A2(n6657), .ZN(n3124) );
  AND4_X4 U3835 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n3125)
         );
  AND2_X2 U3836 ( .A1(n3402), .A2(n3197), .ZN(n3128) );
  NAND2_X2 U3837 ( .A1(n3506), .A2(n3507), .ZN(net222371) );
  INV_X4 U3838 ( .A(net222371), .ZN(n3355) );
  NAND2_X2 U3839 ( .A1(n4475), .A2(n3181), .ZN(n4479) );
  NAND2_X2 U3840 ( .A1(n5356), .A2(\wb/dsize_reg/z2 [31]), .ZN(n4941) );
  INV_X4 U3841 ( .A(n4941), .ZN(n4942) );
  AND2_X2 U3842 ( .A1(n8096), .A2(n2869), .ZN(n3130) );
  NOR2_X2 U3843 ( .A1(n4791), .A2(n4790), .ZN(n4792) );
  NOR2_X2 U3844 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  INV_X8 U3846 ( .A(n2790), .ZN(n3914) );
  INV_X4 U3847 ( .A(n3928), .ZN(n3929) );
  INV_X16 U3848 ( .A(net224865), .ZN(net224859) );
  INV_X4 U3849 ( .A(n2706), .ZN(n3951) );
  INV_X4 U3850 ( .A(net224943), .ZN(net224957) );
  INV_X4 U3851 ( .A(\mem_wb/N41 ), .ZN(net224691) );
  INV_X4 U3852 ( .A(net224717), .ZN(net224611) );
  INV_X4 U3853 ( .A(net224711), .ZN(net224613) );
  INV_X4 U3854 ( .A(net224693), .ZN(net224679) );
  NAND2_X1 U3855 ( .A1(n4442), .A2(iAddr[5]), .ZN(n4448) );
  NAND4_X1 U3856 ( .A1(n6290), .A2(n6289), .A3(n6321), .A4(n6288), .ZN(n6296)
         );
  MUX2_X2 U3857 ( .A(n4703), .B(n3044), .S(n3927), .Z(n2004) );
  BUF_X4 U3858 ( .A(n4156), .Z(n3159) );
  MUX2_X2 U3859 ( .A(n4694), .B(n3049), .S(n3927), .Z(n2013) );
  NAND2_X1 U3860 ( .A1(n4440), .A2(n4473), .ZN(n4441) );
  MUX2_X2 U3861 ( .A(n4700), .B(n3051), .S(n3927), .Z(n2007) );
  INV_X8 U3862 ( .A(n4546), .ZN(n3927) );
  MUX2_X2 U3863 ( .A(n2984), .B(n4707), .S(n3925), .Z(n2000) );
  INV_X4 U3864 ( .A(n4692), .ZN(n3135) );
  INV_X4 U3865 ( .A(n7709), .ZN(n4692) );
  INV_X1 U3866 ( .A(n3965), .ZN(n4394) );
  NAND2_X1 U3867 ( .A1(n2724), .A2(n7707), .ZN(n4615) );
  MUX2_X2 U3868 ( .A(n4708), .B(n3043), .S(n3927), .Z(n1999) );
  AND3_X2 U3869 ( .A1(n4682), .A2(n4587), .A3(n4586), .ZN(n4588) );
  NOR2_X1 U3870 ( .A1(n7427), .A2(n4421), .ZN(n4418) );
  NOR2_X1 U3871 ( .A1(n7427), .A2(n7426), .ZN(n3957) );
  MUX2_X2 U3872 ( .A(n4702), .B(n3009), .S(n3927), .Z(n2005) );
  INV_X1 U3873 ( .A(n4343), .ZN(n3136) );
  INV_X8 U3874 ( .A(n4343), .ZN(n4486) );
  NAND2_X2 U3875 ( .A1(n4505), .A2(n3591), .ZN(n4506) );
  INV_X1 U3876 ( .A(n4544), .ZN(n3591) );
  INV_X2 U3877 ( .A(n4089), .ZN(n4048) );
  MUX2_X2 U3878 ( .A(n4699), .B(n3046), .S(n3927), .Z(n2008) );
  INV_X4 U3879 ( .A(n3927), .ZN(n3925) );
  OAI21_X2 U3880 ( .B1(n4449), .B2(iAddr[6]), .A(n4448), .ZN(n4450) );
  NAND2_X1 U3881 ( .A1(n4094), .A2(n4105), .ZN(n4076) );
  INV_X16 U3882 ( .A(net224999), .ZN(net225216) );
  INV_X16 U3883 ( .A(net224999), .ZN(net225214) );
  NOR2_X2 U3884 ( .A1(n5173), .A2(n4801), .ZN(n5101) );
  INV_X2 U3885 ( .A(n5371), .ZN(n5176) );
  INV_X8 U3886 ( .A(n4178), .ZN(n4323) );
  OAI21_X4 U3887 ( .B1(n4329), .B2(n4328), .A(n4327), .ZN(n4498) );
  NAND2_X4 U3888 ( .A1(n3589), .A2(n4324), .ZN(n4328) );
  AOI21_X4 U3889 ( .B1(n4328), .B2(n4329), .A(n3895), .ZN(n4327) );
  INV_X2 U3890 ( .A(iAddr[21]), .ZN(n4496) );
  NOR2_X2 U3891 ( .A1(n4533), .A2(n4532), .ZN(n4534) );
  INV_X4 U3892 ( .A(net225082), .ZN(net225083) );
  NAND2_X2 U3894 ( .A1(n7906), .A2(iAddr[28]), .ZN(n4316) );
  INV_X4 U3895 ( .A(n3690), .ZN(n3137) );
  INV_X32 U3896 ( .A(n3909), .ZN(n5710) );
  NAND2_X1 U3898 ( .A1(n4500), .A2(iAddr[21]), .ZN(n4502) );
  NOR2_X2 U3899 ( .A1(n7710), .A2(net224955), .ZN(\id_ex/N33 ) );
  NAND2_X4 U3900 ( .A1(n4574), .A2(n7710), .ZN(n6315) );
  INV_X8 U3901 ( .A(n4221), .ZN(n4223) );
  INV_X1 U3903 ( .A(n7519), .ZN(n3140) );
  INV_X2 U3904 ( .A(n3140), .ZN(n3141) );
  NOR2_X2 U3905 ( .A1(n7438), .A2(n3247), .ZN(n4116) );
  INV_X8 U3906 ( .A(n3246), .ZN(n3247) );
  OAI21_X2 U3907 ( .B1(n3156), .B2(n7917), .A(n4140), .ZN(n4143) );
  NOR2_X2 U3908 ( .A1(n7715), .A2(net224899), .ZN(\ex_mem/N35 ) );
  INV_X1 U3909 ( .A(n3726), .ZN(n3144) );
  INV_X4 U3910 ( .A(n3144), .ZN(iAddr[20]) );
  NAND2_X4 U3911 ( .A1(n2741), .A2(n2988), .ZN(n4070) );
  INV_X8 U3912 ( .A(n4044), .ZN(n4077) );
  OR2_X1 U3913 ( .A1(n3553), .A2(n7514), .ZN(n3146) );
  NOR2_X2 U3914 ( .A1(n4002), .A2(n4046), .ZN(n4006) );
  NOR2_X2 U3915 ( .A1(n7657), .A2(net224891), .ZN(\ex_mem/N58 ) );
  NOR2_X1 U3916 ( .A1(net224999), .A2(n5271), .ZN(n5272) );
  NAND2_X4 U3917 ( .A1(n3582), .A2(n3979), .ZN(n3981) );
  INV_X16 U3918 ( .A(n5947), .ZN(n5967) );
  NAND2_X4 U3919 ( .A1(n3862), .A2(n3916), .ZN(n5947) );
  NOR2_X2 U3921 ( .A1(n6725), .A2(n3923), .ZN(n5850) );
  MUX2_X2 U3922 ( .A(n7911), .B(n3048), .S(n3927), .Z(n2014) );
  OAI21_X2 U3923 ( .B1(n4156), .B2(n4155), .A(n4154), .ZN(n4157) );
  AOI21_X2 U3924 ( .B1(n3987), .B2(n4000), .A(n4047), .ZN(n3988) );
  BUF_X8 U3925 ( .A(n4185), .Z(n3150) );
  NAND2_X1 U3927 ( .A1(n3136), .A2(iAddr[16]), .ZN(n4482) );
  MUX2_X2 U3928 ( .A(n6606), .B(n7193), .S(n7205), .Z(n6800) );
  NOR2_X4 U3929 ( .A1(n3232), .A2(n7149), .ZN(n7154) );
  INV_X4 U3931 ( .A(n3152), .ZN(n6543) );
  INV_X2 U3932 ( .A(n4067), .ZN(n4085) );
  OAI211_X4 U3933 ( .C1(n3154), .C2(n6532), .A(n3155), .B(n3153), .ZN(n3152)
         );
  AND2_X4 U3934 ( .A1(n6523), .A2(n2838), .ZN(n3154) );
  NAND2_X1 U3935 ( .A1(n4098), .A2(n4099), .ZN(n3156) );
  AND2_X2 U3936 ( .A1(n4157), .A2(n3894), .ZN(n4158) );
  INV_X4 U3937 ( .A(n3894), .ZN(n3896) );
  AOI211_X2 U3938 ( .C1(n5919), .C2(n5918), .A(n5916), .B(n5917), .ZN(n5922)
         );
  NOR2_X2 U3939 ( .A1(n6672), .A2(n6606), .ZN(n6009) );
  NAND2_X4 U3940 ( .A1(n4165), .A2(n4036), .ZN(n4208) );
  NOR2_X2 U3941 ( .A1(n7665), .A2(net224895), .ZN(\ex_mem/N50 ) );
  NAND3_X2 U3942 ( .A1(n3981), .A2(n2691), .A3(n4152), .ZN(n3984) );
  OAI21_X2 U3943 ( .B1(n5819), .B2(n3950), .A(n5818), .ZN(n5824) );
  NOR2_X2 U3944 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  NAND4_X2 U3945 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n7122)
         );
  NAND3_X4 U3946 ( .A1(n4059), .A2(n4058), .A3(n2961), .ZN(iAddr[14]) );
  INV_X8 U3947 ( .A(iAddr[14]), .ZN(n4477) );
  NAND2_X4 U3948 ( .A1(n5762), .A2(n3955), .ZN(n5747) );
  XOR2_X2 U3949 ( .A(n3385), .B(n7437), .Z(n4458) );
  INV_X2 U3950 ( .A(n4072), .ZN(n4073) );
  NAND3_X4 U3951 ( .A1(iAddr[3]), .A2(iAddr[4]), .A3(iAddr[2]), .ZN(n4453) );
  NAND2_X1 U3952 ( .A1(n7176), .A2(n3878), .ZN(n6665) );
  OAI21_X2 U3953 ( .B1(n3171), .B2(n4150), .A(n4152), .ZN(n4160) );
  INV_X2 U3954 ( .A(n7453), .ZN(n4012) );
  INV_X2 U3955 ( .A(n4050), .ZN(n4055) );
  NAND2_X4 U3956 ( .A1(n5875), .A2(n5874), .ZN(n3878) );
  NOR2_X2 U3957 ( .A1(n3260), .A2(n3954), .ZN(n7119) );
  INV_X8 U3958 ( .A(n5986), .ZN(n6956) );
  NAND2_X4 U3959 ( .A1(n7242), .A2(n3862), .ZN(n5986) );
  MUX2_X2 U3960 ( .A(n4697), .B(n3045), .S(n3927), .Z(n2010) );
  AND3_X4 U3961 ( .A1(n7907), .A2(n7859), .A3(iAddr[24]), .ZN(n4529) );
  NOR2_X2 U3962 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  INV_X4 U3964 ( .A(n7515), .ZN(n4391) );
  INV_X4 U3965 ( .A(n4183), .ZN(n4185) );
  BUF_X32 U3966 ( .A(n6579), .Z(n3160) );
  OAI21_X2 U3967 ( .B1(n2668), .B2(n4103), .A(n4077), .ZN(n4089) );
  NOR4_X1 U3968 ( .A1(n4048), .A2(n4075), .A3(n4047), .A4(n2689), .ZN(n4057)
         );
  AOI21_X2 U3969 ( .B1(n4127), .B2(n4128), .A(n3993), .ZN(n3161) );
  INV_X4 U3970 ( .A(n4128), .ZN(n3994) );
  NAND2_X2 U3971 ( .A1(n4843), .A2(n5413), .ZN(n5416) );
  OAI21_X2 U3972 ( .B1(n3936), .B2(n5417), .A(n5413), .ZN(n5410) );
  AND2_X2 U3973 ( .A1(n3162), .A2(n2965), .ZN(n3164) );
  NOR2_X4 U3974 ( .A1(net225238), .A2(n2967), .ZN(n4882) );
  XNOR2_X2 U3975 ( .A(n4122), .B(n4121), .ZN(n4125) );
  NAND2_X2 U3976 ( .A1(n4126), .A2(n4120), .ZN(n4122) );
  INV_X8 U3977 ( .A(n5838), .ZN(n6725) );
  NAND2_X4 U3978 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  NAND3_X2 U3979 ( .A1(n3460), .A2(n2649), .A3(n5952), .ZN(n3891) );
  NAND2_X1 U3980 ( .A1(n5949), .A2(n6583), .ZN(n3460) );
  NAND3_X2 U3981 ( .A1(n4137), .A2(n4136), .A3(n4135), .ZN(iAddr[9]) );
  OAI211_X4 U3982 ( .C1(n4147), .C2(n3896), .A(n4146), .B(n4145), .ZN(
        iAddr[13]) );
  NOR2_X2 U3983 ( .A1(n6980), .A2(n2701), .ZN(n6024) );
  MUX2_X2 U3984 ( .A(n4747), .B(n7736), .S(net230157), .Z(n3165) );
  INV_X1 U3986 ( .A(n5030), .ZN(n3167) );
  OAI21_X4 U3987 ( .B1(n7205), .B2(n6610), .A(n6006), .ZN(n6007) );
  NOR3_X2 U3988 ( .A1(n7101), .A2(n7099), .A3(n7100), .ZN(n7102) );
  NOR2_X2 U3989 ( .A1(n7098), .A2(n3954), .ZN(n7099) );
  OAI21_X2 U3990 ( .B1(n3260), .B2(n3923), .A(n7079), .ZN(n7101) );
  MUX2_X2 U3991 ( .A(n4695), .B(n3050), .S(n3927), .Z(n2012) );
  XNOR2_X1 U3992 ( .A(n4473), .B(iAddr[13]), .ZN(n4709) );
  BUF_X16 U3993 ( .A(n4356), .Z(n3169) );
  NAND2_X2 U3994 ( .A1(n3583), .A2(n7426), .ZN(n3585) );
  INV_X1 U3995 ( .A(n7426), .ZN(n3584) );
  NAND2_X2 U3996 ( .A1(n3951), .A2(n3539), .ZN(n6970) );
  NAND2_X4 U3998 ( .A1(n6663), .A2(n3878), .ZN(n5879) );
  XNOR2_X1 U3999 ( .A(n7428), .B(n2980), .ZN(n4420) );
  INV_X8 U4000 ( .A(n5858), .ZN(n6939) );
  AND2_X4 U4001 ( .A1(n2696), .A2(n7239), .ZN(n3275) );
  NAND2_X2 U4002 ( .A1(n4934), .A2(n4935), .ZN(n5040) );
  INV_X4 U4003 ( .A(n6165), .ZN(n4934) );
  NOR2_X4 U4004 ( .A1(n5161), .A2(n3267), .ZN(n3266) );
  XNOR2_X1 U4005 ( .A(n7516), .B(n4389), .ZN(n4390) );
  INV_X1 U4006 ( .A(n4208), .ZN(n4210) );
  NOR2_X4 U4007 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NOR2_X2 U4008 ( .A1(n3914), .A2(n6607), .ZN(n6008) );
  AOI21_X2 U4009 ( .B1(n6835), .B2(n3921), .A(n6764), .ZN(n6765) );
  INV_X8 U4010 ( .A(n6660), .ZN(n6619) );
  BUF_X8 U4011 ( .A(n5663), .Z(n3511) );
  INV_X4 U4012 ( .A(n3879), .ZN(n3880) );
  NOR2_X2 U4013 ( .A1(n6123), .A2(n6122), .ZN(n6135) );
  NAND3_X4 U4014 ( .A1(n7198), .A2(n3888), .A3(n5965), .ZN(n5966) );
  NAND2_X4 U4015 ( .A1(n7242), .A2(n5960), .ZN(n7198) );
  NAND2_X2 U4016 ( .A1(n7127), .A2(n6545), .ZN(n6379) );
  MUX2_X2 U4017 ( .A(n6669), .B(n7255), .S(n7205), .Z(n6859) );
  NAND2_X2 U4019 ( .A1(n2681), .A2(n7176), .ZN(n6437) );
  INV_X8 U4020 ( .A(n3270), .ZN(n6608) );
  NAND2_X4 U4021 ( .A1(n3311), .A2(n5992), .ZN(n3170) );
  NAND2_X2 U4022 ( .A1(n3311), .A2(n5992), .ZN(n3310) );
  NAND2_X4 U4024 ( .A1(n6477), .A2(n3395), .ZN(n6964) );
  NAND2_X4 U4026 ( .A1(n4062), .A2(n4347), .ZN(n3519) );
  NAND2_X2 U4027 ( .A1(n4134), .A2(n4156), .ZN(n3171) );
  INV_X4 U4028 ( .A(n5722), .ZN(n3172) );
  NAND2_X4 U4029 ( .A1(n3887), .A2(n7169), .ZN(n3311) );
  NOR2_X2 U4030 ( .A1(n6800), .A2(n3923), .ZN(n6387) );
  NOR2_X2 U4031 ( .A1(n6800), .A2(n3954), .ZN(n6653) );
  NOR2_X2 U4032 ( .A1(n6800), .A2(n2701), .ZN(n6782) );
  INV_X2 U4033 ( .A(n6800), .ZN(n6802) );
  AOI211_X2 U4034 ( .C1(n6389), .C2(n6388), .A(n6387), .B(n6386), .ZN(n6484)
         );
  NOR2_X4 U4035 ( .A1(n5918), .A2(n5154), .ZN(n5158) );
  NAND2_X2 U4036 ( .A1(n6621), .A2(n6663), .ZN(n6516) );
  INV_X4 U4037 ( .A(n3173), .ZN(n3174) );
  NOR2_X2 U4038 ( .A1(n7633), .A2(net224901), .ZN(\ex_mem/N44 ) );
  OAI21_X4 U4039 ( .B1(n4820), .B2(net223242), .A(n4819), .ZN(n4821) );
  INV_X1 U4040 ( .A(n3160), .ZN(n4833) );
  INV_X8 U4041 ( .A(n6602), .ZN(n6667) );
  NAND2_X2 U4042 ( .A1(n5873), .A2(n3922), .ZN(n5863) );
  NAND3_X1 U4043 ( .A1(n4499), .A2(n4497), .A3(n4498), .ZN(iAddr[22]) );
  AOI21_X1 U4044 ( .B1(n4154), .B2(n7916), .A(n4138), .ZN(n4140) );
  NAND2_X2 U4045 ( .A1(net222161), .A2(net229596), .ZN(n3202) );
  NAND2_X4 U4046 ( .A1(n4338), .A2(n4524), .ZN(n4436) );
  BUF_X4 U4047 ( .A(n3283), .Z(n3175) );
  NAND2_X2 U4048 ( .A1(n6930), .A2(n7001), .ZN(n3176) );
  NAND2_X2 U4049 ( .A1(n7001), .A2(n6930), .ZN(n7338) );
  NAND2_X2 U4050 ( .A1(n3643), .A2(memAddr[17]), .ZN(n3678) );
  OAI21_X4 U4051 ( .B1(n4742), .B2(net230741), .A(n4741), .ZN(n6060) );
  INV_X4 U4052 ( .A(n6107), .ZN(n3508) );
  NAND2_X4 U4053 ( .A1(n6868), .A2(n6869), .ZN(n6871) );
  MUX2_X2 U4055 ( .A(memRdData[26]), .B(\wb/dsize_reg/z2 [26]), .S(net224723), 
        .Z(n2241) );
  NAND3_X1 U4056 ( .A1(n4483), .A2(n4484), .A3(n4485), .ZN(iAddr[18]) );
  INV_X4 U4057 ( .A(n3177), .ZN(n3178) );
  NOR2_X2 U4058 ( .A1(n7663), .A2(net224895), .ZN(\ex_mem/N52 ) );
  INV_X1 U4059 ( .A(n2621), .ZN(n6708) );
  INV_X2 U4060 ( .A(net228940), .ZN(net228942) );
  INV_X8 U4061 ( .A(n4844), .ZN(n5111) );
  INV_X1 U4062 ( .A(n2582), .ZN(n6532) );
  NAND2_X1 U4063 ( .A1(net225237), .A2(reg31Val_0[25]), .ZN(n4757) );
  INV_X1 U4064 ( .A(n6390), .ZN(n3179) );
  NAND2_X2 U4066 ( .A1(n3212), .A2(n3843), .ZN(n3370) );
  NAND2_X4 U4067 ( .A1(n3370), .A2(n3371), .ZN(n6139) );
  NAND2_X2 U4068 ( .A1(n6944), .A2(n3293), .ZN(n5718) );
  INV_X4 U4069 ( .A(n6853), .ZN(n6086) );
  NOR3_X4 U4070 ( .A1(n6024), .A2(n6025), .A3(n6023), .ZN(n6026) );
  NAND2_X2 U4071 ( .A1(n5146), .A2(n5145), .ZN(n5052) );
  XNOR2_X1 U4072 ( .A(n7913), .B(n3070), .ZN(n3180) );
  INV_X1 U4073 ( .A(n4477), .ZN(n3181) );
  INV_X2 U4075 ( .A(n7282), .ZN(n6573) );
  NAND2_X4 U4077 ( .A1(n3183), .A2(n5952), .ZN(n6941) );
  INV_X4 U4078 ( .A(n3182), .ZN(n3183) );
  NAND2_X2 U4079 ( .A1(n3426), .A2(n5869), .ZN(n5953) );
  NAND2_X2 U4080 ( .A1(n2588), .A2(n5366), .ZN(n5078) );
  NAND2_X2 U4081 ( .A1(n6062), .A2(n3184), .ZN(n3185) );
  NAND2_X1 U4082 ( .A1(n7736), .A2(net225434), .ZN(n3186) );
  NAND2_X4 U4083 ( .A1(n3185), .A2(n3186), .ZN(n6063) );
  INV_X1 U4084 ( .A(net225434), .ZN(n3184) );
  NAND2_X1 U4085 ( .A1(n6059), .A2(net224861), .ZN(n3189) );
  NAND2_X2 U4086 ( .A1(n3189), .A2(n3190), .ZN(net221757) );
  INV_X4 U4087 ( .A(n6059), .ZN(n3187) );
  INV_X1 U4088 ( .A(net224861), .ZN(n3188) );
  NAND2_X2 U4089 ( .A1(n3191), .A2(n3192), .ZN(n3194) );
  NAND2_X4 U4090 ( .A1(n3193), .A2(n3194), .ZN(net220619) );
  INV_X2 U4091 ( .A(net220651), .ZN(n3192) );
  NOR2_X4 U4092 ( .A1(n6162), .A2(n6163), .ZN(n6168) );
  NAND2_X2 U4093 ( .A1(n7327), .A2(n7326), .ZN(n7328) );
  NAND3_X1 U4095 ( .A1(net221442), .A2(n6401), .A3(n3549), .ZN(n6402) );
  NAND3_X1 U4096 ( .A1(net223339), .A2(net223338), .A3(n3279), .ZN(net222161)
         );
  NAND2_X4 U4097 ( .A1(n5843), .A2(net220849), .ZN(n7004) );
  INV_X4 U4098 ( .A(n3555), .ZN(n3556) );
  NAND3_X4 U4099 ( .A1(n3871), .A2(n3872), .A3(n3873), .ZN(n3870) );
  INV_X8 U4100 ( .A(n3870), .ZN(n5228) );
  AOI22_X2 U4101 ( .A1(n4894), .A2(net225047), .B1(n4893), .B2(net225047), 
        .ZN(n5047) );
  NAND2_X1 U4103 ( .A1(n6634), .A2(n3272), .ZN(n3210) );
  NAND2_X2 U4104 ( .A1(n6631), .A2(n6411), .ZN(n3430) );
  INV_X4 U4106 ( .A(n3502), .ZN(n3383) );
  XNOR2_X1 U4108 ( .A(n7997), .B(net228715), .ZN(net230245) );
  INV_X2 U4109 ( .A(n3647), .ZN(n3648) );
  INV_X8 U4110 ( .A(n4859), .ZN(n5189) );
  OR2_X2 U4111 ( .A1(n7297), .A2(n7296), .ZN(n3195) );
  INV_X1 U4112 ( .A(n7181), .ZN(n3196) );
  INV_X4 U4113 ( .A(n6839), .ZN(n7295) );
  INV_X4 U4114 ( .A(n7179), .ZN(n7181) );
  NAND2_X2 U4115 ( .A1(n5487), .A2(n5821), .ZN(n3198) );
  NAND2_X4 U4116 ( .A1(n3198), .A2(n3199), .ZN(n3634) );
  INV_X8 U4117 ( .A(n5821), .ZN(n3197) );
  NAND4_X4 U4118 ( .A1(n5143), .A2(n3201), .A3(n5142), .A4(n5144), .ZN(n5166)
         );
  NAND2_X2 U4119 ( .A1(n2844), .A2(net223245), .ZN(n3677) );
  OAI221_X4 U4120 ( .B1(n7521), .B2(n4465), .C1(n4087), .C2(n3895), .A(n4086), 
        .ZN(n8109) );
  NAND2_X2 U4121 ( .A1(n2900), .A2(net228981), .ZN(n3203) );
  NAND2_X4 U4122 ( .A1(n3202), .A2(n3203), .ZN(net222155) );
  INV_X4 U4123 ( .A(n3802), .ZN(n3803) );
  BUF_X8 U4124 ( .A(n5813), .Z(n3204) );
  INV_X4 U4125 ( .A(n4924), .ZN(n3206) );
  NAND2_X1 U4126 ( .A1(n4950), .A2(net224995), .ZN(n4951) );
  AOI21_X2 U4127 ( .B1(n3955), .B2(n6602), .A(n5999), .ZN(n6000) );
  AOI21_X4 U4128 ( .B1(net225216), .B2(n3550), .A(n2676), .ZN(n3549) );
  OAI211_X1 U4131 ( .C1(n7142), .C2(n7141), .A(n7143), .B(n3672), .ZN(n7147)
         );
  NAND2_X1 U4132 ( .A1(n3955), .A2(n6514), .ZN(n5789) );
  INV_X2 U4134 ( .A(n4886), .ZN(n5156) );
  NAND2_X4 U4135 ( .A1(n4851), .A2(n4850), .ZN(n5382) );
  INV_X1 U4136 ( .A(n7476), .ZN(n4867) );
  NOR3_X2 U4137 ( .A1(n6833), .A2(n6832), .A3(n6831), .ZN(n6834) );
  INV_X8 U4138 ( .A(n5359), .ZN(n3785) );
  AOI21_X1 U4139 ( .B1(net224843), .B2(n3323), .A(net224835), .ZN(net221858)
         );
  AOI21_X1 U4140 ( .B1(net221862), .B2(n2838), .A(n3323), .ZN(net221856) );
  NAND2_X2 U4141 ( .A1(n3323), .A2(net221864), .ZN(n3329) );
  INV_X2 U4142 ( .A(n3323), .ZN(n3327) );
  NAND2_X4 U4143 ( .A1(n6098), .A2(n6663), .ZN(n6099) );
  NAND2_X4 U4144 ( .A1(n3209), .A2(net228715), .ZN(n3211) );
  NAND2_X4 U4145 ( .A1(n3210), .A2(n3211), .ZN(n6411) );
  NAND2_X2 U4146 ( .A1(n3825), .A2(n3212), .ZN(n3213) );
  NAND2_X2 U4147 ( .A1(n7731), .A2(n3299), .ZN(n3214) );
  INV_X4 U4148 ( .A(n3299), .ZN(n3212) );
  INV_X2 U4149 ( .A(net224735), .ZN(n3299) );
  NAND3_X2 U4150 ( .A1(n5184), .A2(n5185), .A3(n5142), .ZN(n5186) );
  INV_X32 U4151 ( .A(n3934), .ZN(n3933) );
  NOR2_X2 U4152 ( .A1(net225015), .A2(n5389), .ZN(n5390) );
  NOR2_X4 U4153 ( .A1(n7942), .A2(n3217), .ZN(n3215) );
  INV_X4 U4154 ( .A(n3215), .ZN(n5154) );
  AND2_X4 U4155 ( .A1(n2932), .A2(net229784), .ZN(n3217) );
  NOR2_X4 U4156 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  INV_X8 U4157 ( .A(n6392), .ZN(n3829) );
  NAND2_X4 U4158 ( .A1(n2646), .A2(net229005), .ZN(n6885) );
  NAND4_X4 U4159 ( .A1(n5068), .A2(net224737), .A3(n5067), .A4(n5066), .ZN(
        n5069) );
  NAND2_X4 U4160 ( .A1(n2635), .A2(n3218), .ZN(n3219) );
  NAND2_X4 U4161 ( .A1(n3219), .A2(n4744), .ZN(n6061) );
  INV_X1 U4162 ( .A(net230741), .ZN(n3218) );
  NAND2_X2 U4164 ( .A1(n4743), .A2(net225047), .ZN(n4744) );
  NAND2_X2 U4166 ( .A1(n3221), .A2(n6124), .ZN(n6936) );
  INV_X4 U4167 ( .A(n3220), .ZN(n3221) );
  INV_X8 U4168 ( .A(n6845), .ZN(n6840) );
  NAND2_X1 U4169 ( .A1(n7358), .A2(n6175), .ZN(n6176) );
  INV_X4 U4170 ( .A(n6878), .ZN(n6897) );
  OAI21_X4 U4172 ( .B1(n3683), .B2(n5795), .A(n3615), .ZN(n5797) );
  NAND3_X2 U4173 ( .A1(n2691), .A2(n3981), .A3(n4152), .ZN(n3223) );
  NAND2_X4 U4174 ( .A1(n3723), .A2(n3149), .ZN(n4152) );
  INV_X4 U4175 ( .A(n7213), .ZN(n3953) );
  OAI211_X2 U4176 ( .C1(n6552), .C2(n3615), .A(n3765), .B(n6699), .ZN(n5898)
         );
  NAND2_X2 U4177 ( .A1(n6421), .A2(n3631), .ZN(n3227) );
  NAND2_X4 U4178 ( .A1(n3225), .A2(n3226), .ZN(n3228) );
  NAND2_X4 U4179 ( .A1(n3227), .A2(n3228), .ZN(n7335) );
  INV_X4 U4180 ( .A(n6421), .ZN(n3225) );
  INV_X4 U4181 ( .A(n3631), .ZN(n3226) );
  NAND2_X2 U4182 ( .A1(n3229), .A2(n5203), .ZN(n3230) );
  NAND2_X2 U4183 ( .A1(n2763), .A2(net229173), .ZN(n3231) );
  INV_X4 U4185 ( .A(net229173), .ZN(n3229) );
  INV_X1 U4186 ( .A(net224735), .ZN(net229173) );
  INV_X4 U4187 ( .A(n3774), .ZN(n3775) );
  NAND2_X4 U4188 ( .A1(net224737), .A2(n3449), .ZN(n6395) );
  CLKBUF_X3 U4189 ( .A(n7301), .Z(n3232) );
  INV_X4 U4190 ( .A(n6919), .ZN(n3233) );
  NAND2_X4 U4192 ( .A1(n3235), .A2(n3234), .ZN(n3237) );
  NAND2_X4 U4193 ( .A1(n3236), .A2(n3237), .ZN(n6391) );
  INV_X1 U4194 ( .A(net227884), .ZN(n3234) );
  INV_X4 U4195 ( .A(n6423), .ZN(n3235) );
  INV_X1 U4196 ( .A(n4537), .ZN(n3238) );
  INV_X4 U4197 ( .A(n4512), .ZN(n3239) );
  MUX2_X1 U4198 ( .A(n3054), .B(n4698), .S(n3926), .Z(n2009) );
  NAND2_X4 U4199 ( .A1(n3343), .A2(n3342), .ZN(n3345) );
  INV_X4 U4200 ( .A(n3548), .ZN(n5895) );
  MUX2_X2 U4201 ( .A(n4701), .B(n3084), .S(n3927), .Z(n2006) );
  INV_X4 U4202 ( .A(n3927), .ZN(n3926) );
  NAND2_X4 U4203 ( .A1(n3364), .A2(n3365), .ZN(n5485) );
  INV_X16 U4204 ( .A(n7053), .ZN(n6985) );
  NAND2_X2 U4205 ( .A1(n7053), .A2(n3652), .ZN(n6041) );
  NOR2_X2 U4206 ( .A1(n7724), .A2(net224897), .ZN(\ex_mem/N142 ) );
  NAND2_X1 U4207 ( .A1(net224865), .A2(n6112), .ZN(n3244) );
  NAND2_X4 U4208 ( .A1(n3242), .A2(n3243), .ZN(n3245) );
  NAND2_X4 U4209 ( .A1(n3244), .A2(n3245), .ZN(n6113) );
  INV_X2 U4210 ( .A(n6112), .ZN(n3243) );
  NAND2_X4 U4211 ( .A1(n3530), .A2(n7932), .ZN(n4127) );
  INV_X4 U4212 ( .A(n7433), .ZN(n3246) );
  NAND4_X4 U4213 ( .A1(n5748), .A2(n5749), .A3(n5750), .A4(n5747), .ZN(n6521)
         );
  XNOR2_X2 U4215 ( .A(n6059), .B(net224861), .ZN(n3269) );
  INV_X4 U4216 ( .A(n6189), .ZN(n5974) );
  NAND2_X4 U4217 ( .A1(n6487), .A2(n2615), .ZN(n3284) );
  NAND2_X4 U4218 ( .A1(net220312), .A2(net220313), .ZN(n3249) );
  INV_X4 U4219 ( .A(n6167), .ZN(n3408) );
  NAND2_X2 U4220 ( .A1(n3537), .A2(n3538), .ZN(n3250) );
  NAND2_X2 U4221 ( .A1(n3538), .A2(n3537), .ZN(n7323) );
  NOR2_X1 U4222 ( .A1(n3950), .A2(n7326), .ZN(n7067) );
  NAND2_X4 U4223 ( .A1(n3598), .A2(n3599), .ZN(n5205) );
  AOI21_X1 U4224 ( .B1(n4478), .B2(n4477), .A(n4476), .ZN(n4708) );
  INV_X1 U4225 ( .A(n3552), .ZN(n4401) );
  NAND3_X2 U4226 ( .A1(n7055), .A2(n3204), .A3(n3424), .ZN(n7138) );
  INV_X16 U4227 ( .A(net221652), .ZN(net230144) );
  NAND2_X4 U4228 ( .A1(n3732), .A2(net229719), .ZN(n3574) );
  OAI21_X2 U4229 ( .B1(n3850), .B2(n3170), .A(n7239), .ZN(n7251) );
  NAND2_X2 U4230 ( .A1(n4862), .A2(n4863), .ZN(n4864) );
  INV_X8 U4231 ( .A(n5065), .ZN(n5066) );
  NOR2_X4 U4233 ( .A1(net225238), .A2(n2937), .ZN(n4866) );
  OAI21_X4 U4234 ( .B1(n4129), .B2(n3377), .A(n4127), .ZN(n4130) );
  INV_X16 U4235 ( .A(n3939), .ZN(n3938) );
  INV_X8 U4239 ( .A(n4349), .ZN(n4238) );
  INV_X4 U4240 ( .A(n6531), .ZN(n3635) );
  NAND2_X2 U4241 ( .A1(n3406), .A2(n6531), .ZN(n3636) );
  NOR2_X4 U4242 ( .A1(n3263), .A2(net224871), .ZN(n5345) );
  NAND2_X1 U4243 ( .A1(n5080), .A2(n3257), .ZN(n3258) );
  NAND2_X2 U4244 ( .A1(n7732), .A2(net227817), .ZN(n3259) );
  NAND2_X2 U4245 ( .A1(n3258), .A2(n3259), .ZN(n5206) );
  INV_X4 U4246 ( .A(net227817), .ZN(n3257) );
  INV_X8 U4247 ( .A(n3851), .ZN(n5080) );
  INV_X1 U4248 ( .A(net224735), .ZN(net227817) );
  NOR2_X2 U4249 ( .A1(n5333), .A2(n7943), .ZN(n5335) );
  INV_X4 U4250 ( .A(n4858), .ZN(n3307) );
  INV_X2 U4251 ( .A(n6620), .ZN(n5721) );
  NOR2_X1 U4252 ( .A1(n7302), .A2(n3950), .ZN(n6831) );
  NAND4_X2 U4253 ( .A1(net224737), .A2(n5004), .A3(n3907), .A4(n5003), .ZN(
        n5545) );
  OAI21_X1 U4254 ( .B1(net224833), .B2(n7152), .A(n5154), .ZN(n7153) );
  INV_X2 U4255 ( .A(n7959), .ZN(n3482) );
  INV_X4 U4256 ( .A(n6185), .ZN(n6568) );
  NAND2_X2 U4257 ( .A1(n5234), .A2(n5440), .ZN(n5237) );
  NAND2_X2 U4258 ( .A1(n5368), .A2(n5440), .ZN(n5370) );
  NAND2_X2 U4259 ( .A1(n6462), .A2(n6504), .ZN(n5288) );
  NAND2_X2 U4260 ( .A1(n3773), .A2(n6462), .ZN(n5854) );
  NOR2_X2 U4261 ( .A1(net221878), .A2(net221425), .ZN(n3326) );
  NOR2_X2 U4262 ( .A1(net221762), .A2(net221425), .ZN(net221761) );
  NAND2_X4 U4264 ( .A1(n3264), .A2(n5325), .ZN(n5304) );
  NAND2_X4 U4265 ( .A1(n5084), .A2(n3265), .ZN(n3264) );
  NOR2_X4 U4266 ( .A1(n3412), .A2(net224747), .ZN(n3265) );
  NAND2_X4 U4267 ( .A1(n5042), .A2(n3266), .ZN(n5046) );
  INV_X1 U4268 ( .A(n8013), .ZN(n5756) );
  OAI222_X1 U4269 ( .A1(n7382), .A2(net224767), .B1(net224755), .B2(n2736), 
        .C1(net224773), .C2(n7540), .ZN(memWrData[21]) );
  NAND2_X4 U4270 ( .A1(n5257), .A2(n6232), .ZN(n5351) );
  NAND3_X2 U4271 ( .A1(n6232), .A2(n6231), .A3(n6230), .ZN(regWrData[8]) );
  NAND2_X4 U4272 ( .A1(n3738), .A2(n3739), .ZN(n3268) );
  NAND2_X2 U4273 ( .A1(n5303), .A2(n3746), .ZN(n5086) );
  NAND3_X2 U4274 ( .A1(n5532), .A2(n5531), .A3(n5530), .ZN(n5536) );
  NAND2_X4 U4275 ( .A1(n3397), .A2(n5531), .ZN(n5061) );
  INV_X8 U4276 ( .A(n5534), .ZN(n5531) );
  INV_X8 U4277 ( .A(n4854), .ZN(n5132) );
  NAND2_X2 U4278 ( .A1(n6788), .A2(n6944), .ZN(n6465) );
  NOR3_X2 U4280 ( .A1(n3935), .A2(n5386), .A3(n3920), .ZN(n5391) );
  NOR2_X4 U4283 ( .A1(net229481), .A2(n6120), .ZN(n3271) );
  OAI21_X2 U4284 ( .B1(n5122), .B2(n5121), .A(n5330), .ZN(n5196) );
  OAI21_X2 U4285 ( .B1(n5978), .B2(n3560), .A(n6956), .ZN(n5979) );
  NAND2_X4 U4286 ( .A1(n3430), .A2(n3431), .ZN(n6873) );
  NAND2_X4 U4287 ( .A1(n3428), .A2(n3429), .ZN(n3431) );
  INV_X2 U4288 ( .A(n3755), .ZN(n3523) );
  AOI21_X4 U4289 ( .B1(net225216), .B2(n3550), .A(n3551), .ZN(n3273) );
  NAND4_X2 U4290 ( .A1(n5221), .A2(n5220), .A3(n3811), .A4(n3208), .ZN(n5222)
         );
  OAI22_X2 U4291 ( .A1(n7411), .A2(n3912), .B1(n7699), .B2(n3909), .ZN(n5653)
         );
  XNOR2_X2 U4294 ( .A(n3278), .B(n3137), .ZN(n3277) );
  INV_X4 U4295 ( .A(n3277), .ZN(n7300) );
  NAND2_X2 U4296 ( .A1(n6732), .A2(n6731), .ZN(n3278) );
  AOI21_X4 U4297 ( .B1(net223341), .B2(net225251), .A(net223342), .ZN(n3279)
         );
  OAI21_X4 U4298 ( .B1(net225243), .B2(net33280), .A(net223343), .ZN(net223342) );
  NAND2_X4 U4300 ( .A1(n5036), .A2(n3407), .ZN(n3280) );
  INV_X2 U4301 ( .A(n5342), .ZN(n5349) );
  INV_X2 U4302 ( .A(n7084), .ZN(n5843) );
  XNOR2_X2 U4303 ( .A(n3281), .B(n7499), .ZN(n3974) );
  OAI22_X4 U4304 ( .A1(n2699), .A2(n4759), .B1(n3252), .B2(n4758), .ZN(n5065)
         );
  NAND2_X2 U4305 ( .A1(net225237), .A2(\wb/dsize_reg/z2 [25]), .ZN(n4759) );
  INV_X16 U4306 ( .A(net225055), .ZN(net225251) );
  INV_X1 U4307 ( .A(n6706), .ZN(n3522) );
  NAND2_X4 U4308 ( .A1(n5566), .A2(n5485), .ZN(n5488) );
  NOR2_X2 U4309 ( .A1(net224745), .A2(n5311), .ZN(n5305) );
  AOI21_X4 U4310 ( .B1(n5311), .B2(n3746), .A(net224745), .ZN(n5089) );
  INV_X8 U4311 ( .A(net224789), .ZN(n3283) );
  INV_X16 U4312 ( .A(net224789), .ZN(net224787) );
  NAND2_X2 U4313 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  NAND2_X4 U4314 ( .A1(n4093), .A2(n4094), .ZN(n4103) );
  OAI211_X4 U4315 ( .C1(net225015), .C2(n7973), .A(n4843), .B(n5413), .ZN(
        n4844) );
  NAND2_X2 U4316 ( .A1(n5551), .A2(n5550), .ZN(n3617) );
  NAND2_X2 U4317 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  NAND2_X4 U4318 ( .A1(net228707), .A2(net228708), .ZN(net228710) );
  NOR2_X4 U4319 ( .A1(n3625), .A2(n6647), .ZN(n6648) );
  NAND2_X1 U4320 ( .A1(n6470), .A2(n3948), .ZN(n5942) );
  NOR2_X1 U4321 ( .A1(n7569), .A2(net225015), .ZN(n6237) );
  INV_X1 U4322 ( .A(n6598), .ZN(n3285) );
  OAI21_X4 U4324 ( .B1(n3288), .B2(n3289), .A(n3287), .ZN(n3286) );
  INV_X4 U4325 ( .A(n3286), .ZN(n5565) );
  OR2_X1 U4326 ( .A1(n5559), .A2(n5563), .ZN(n3288) );
  OR2_X2 U4327 ( .A1(n5562), .A2(n5561), .ZN(n3289) );
  NOR2_X1 U4328 ( .A1(n3710), .A2(n2734), .ZN(n4785) );
  INV_X8 U4329 ( .A(net225229), .ZN(n3290) );
  INV_X4 U4330 ( .A(net225229), .ZN(net225230) );
  OAI22_X1 U4331 ( .A1(n7747), .A2(net224943), .B1(n4658), .B2(n4656), .ZN(
        n7883) );
  NAND2_X1 U4332 ( .A1(n7030), .A2(n7358), .ZN(n7031) );
  NOR2_X1 U4333 ( .A1(n7030), .A2(n6686), .ZN(n6338) );
  NAND3_X2 U4334 ( .A1(n4778), .A2(net228287), .A3(net225045), .ZN(n5073) );
  INV_X8 U4335 ( .A(net224991), .ZN(n3291) );
  INV_X4 U4336 ( .A(n5014), .ZN(n3855) );
  INV_X16 U4337 ( .A(net224997), .ZN(net224991) );
  INV_X8 U4339 ( .A(n7083), .ZN(n7086) );
  NOR2_X4 U4340 ( .A1(n3485), .A2(n5187), .ZN(n5139) );
  NAND2_X4 U4342 ( .A1(n5759), .A2(n7172), .ZN(n5971) );
  AOI21_X2 U4343 ( .B1(n7172), .B2(n2649), .A(n7201), .ZN(n7173) );
  NAND2_X2 U4344 ( .A1(n5491), .A2(n5492), .ZN(n5495) );
  NAND2_X1 U4345 ( .A1(n5429), .A2(n5428), .ZN(n3294) );
  NOR2_X4 U4346 ( .A1(n6401), .A2(n3920), .ZN(n6398) );
  INV_X2 U4347 ( .A(n6404), .ZN(n6405) );
  NAND2_X1 U4348 ( .A1(n3746), .A2(n5325), .ZN(n5327) );
  AOI21_X1 U4349 ( .B1(n5177), .B2(n5176), .A(n5445), .ZN(n5181) );
  OAI21_X2 U4351 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n6830) );
  BUF_X32 U4352 ( .A(n4337), .Z(n3546) );
  NAND2_X4 U4353 ( .A1(n3656), .A2(n3657), .ZN(n3295) );
  INV_X1 U4354 ( .A(net221153), .ZN(n3296) );
  OAI21_X4 U4356 ( .B1(n5375), .B2(n5376), .A(n3615), .ZN(n5435) );
  INV_X1 U4357 ( .A(net229071), .ZN(n3297) );
  INV_X1 U4358 ( .A(net228597), .ZN(n3298) );
  NAND2_X4 U4359 ( .A1(n5958), .A2(n5959), .ZN(n3753) );
  NAND2_X2 U4361 ( .A1(n5948), .A2(n6944), .ZN(n5664) );
  INV_X1 U4362 ( .A(n6500), .ZN(n4855) );
  NOR2_X2 U4363 ( .A1(n7545), .A2(net225015), .ZN(n4940) );
  NAND3_X2 U4364 ( .A1(n2603), .A2(n4989), .A3(net224731), .ZN(n5567) );
  INV_X16 U4365 ( .A(net224743), .ZN(net224731) );
  NAND3_X1 U4366 ( .A1(n4053), .A2(n4049), .A3(n4052), .ZN(n4056) );
  XNOR2_X2 U4367 ( .A(n6715), .B(n6553), .ZN(n3300) );
  NAND2_X4 U4368 ( .A1(n2614), .A2(n3799), .ZN(n3301) );
  NAND2_X4 U4369 ( .A1(n2604), .A2(net220637), .ZN(n7083) );
  NOR2_X2 U4371 ( .A1(n7018), .A2(n7024), .ZN(n3303) );
  NAND2_X4 U4372 ( .A1(net230730), .A2(net221416), .ZN(n3340) );
  INV_X8 U4373 ( .A(n6985), .ZN(n3776) );
  NAND2_X4 U4374 ( .A1(n7054), .A2(n6985), .ZN(n5511) );
  NAND2_X4 U4375 ( .A1(n6890), .A2(n6141), .ZN(n6639) );
  CLKBUF_X3 U4376 ( .A(n6890), .Z(n3661) );
  NAND2_X4 U4377 ( .A1(net220780), .A2(net230245), .ZN(n6890) );
  NAND2_X4 U4379 ( .A1(n6931), .A2(n3176), .ZN(n3305) );
  NAND2_X2 U4380 ( .A1(n6931), .A2(n3176), .ZN(net220313) );
  INV_X4 U4381 ( .A(n5199), .ZN(n3645) );
  NAND2_X4 U4382 ( .A1(n4857), .A2(n3306), .ZN(n4859) );
  NAND3_X2 U4383 ( .A1(n4856), .A2(\wb/dsize_reg/z2 [30]), .A3(n3898), .ZN(
        n4858) );
  INV_X32 U4384 ( .A(n3862), .ZN(n7201) );
  OAI21_X1 U4385 ( .B1(net221488), .B2(net221489), .A(net221490), .ZN(
        net221487) );
  INV_X8 U4386 ( .A(n6637), .ZN(n6631) );
  OAI21_X4 U4387 ( .B1(n5673), .B2(n6257), .A(n5672), .ZN(n3309) );
  NAND3_X2 U4388 ( .A1(n3888), .A2(n5988), .A3(n5987), .ZN(n3887) );
  AOI22_X4 U4390 ( .A1(net223245), .A2(n2708), .B1(n7995), .B2(memAddr[29]), 
        .ZN(n4819) );
  OAI22_X2 U4392 ( .A1(n7420), .A2(n3911), .B1(n7689), .B2(n3909), .ZN(n5514)
         );
  NAND2_X1 U4393 ( .A1(n4148), .A2(n3546), .ZN(n4150) );
  INV_X1 U4394 ( .A(n7001), .ZN(n7017) );
  NOR2_X1 U4396 ( .A1(n3952), .A2(n2703), .ZN(n7194) );
  INV_X8 U4397 ( .A(n6521), .ZN(n6546) );
  AOI22_X1 U4398 ( .A1(memAddr[21]), .A2(n3910), .B1(n7603), .B2(n3908), .ZN(
        n3314) );
  INV_X2 U4399 ( .A(n3314), .ZN(n6054) );
  AOI22_X4 U4400 ( .A1(n3910), .A2(memAddr[7]), .B1(n5710), .B2(n7605), .ZN(
        net228921) );
  NAND3_X2 U4401 ( .A1(n5189), .A2(n5190), .A3(net33207), .ZN(n5191) );
  AND3_X4 U4402 ( .A1(n4276), .A2(n4290), .A3(n3466), .ZN(n4028) );
  NAND3_X2 U4403 ( .A1(net221875), .A2(net221876), .A3(net220875), .ZN(
        net229737) );
  NOR2_X4 U4404 ( .A1(net220285), .A2(net220286), .ZN(net133771) );
  OAI21_X4 U4405 ( .B1(net220287), .B2(net220288), .A(net220289), .ZN(
        net220286) );
  NAND2_X4 U4406 ( .A1(n3315), .A2(n3316), .ZN(net220289) );
  INV_X2 U4407 ( .A(net220292), .ZN(n3316) );
  INV_X2 U4408 ( .A(net220293), .ZN(n3315) );
  NAND2_X4 U4409 ( .A1(net220409), .A2(net228541), .ZN(net220288) );
  NOR3_X4 U4410 ( .A1(net220294), .A2(net220295), .A3(net220296), .ZN(
        net220287) );
  OAI221_X2 U4411 ( .B1(net220297), .B2(net220298), .C1(net220299), .C2(
        net220300), .A(net220301), .ZN(net220296) );
  AOI221_X1 U4412 ( .B1(n3317), .B2(n2848), .C1(n3318), .C2(n3255), .A(n2839), 
        .ZN(net220301) );
  INV_X4 U4413 ( .A(net33219), .ZN(n3321) );
  INV_X4 U4414 ( .A(n3320), .ZN(n3318) );
  OAI211_X2 U4415 ( .C1(net220310), .C2(net220307), .A(setInv_2), .B(n2841), 
        .ZN(n3320) );
  NAND2_X2 U4416 ( .A1(net224957), .A2(n2841), .ZN(net223781) );
  INV_X1 U4417 ( .A(net220305), .ZN(net220307) );
  NAND2_X2 U4419 ( .A1(net220307), .A2(n2848), .ZN(net220354) );
  NAND3_X2 U4420 ( .A1(net228677), .A2(n3305), .A3(net220314), .ZN(net220300)
         );
  INV_X4 U4421 ( .A(net220354), .ZN(net220314) );
  NAND2_X2 U4422 ( .A1(net220314), .A2(n3305), .ZN(net228093) );
  NAND2_X4 U4423 ( .A1(net229736), .A2(net229737), .ZN(net220323) );
  NAND2_X4 U4424 ( .A1(n3329), .A2(n3330), .ZN(net221769) );
  INV_X8 U4425 ( .A(net221769), .ZN(net220875) );
  NAND2_X2 U4426 ( .A1(net220876), .A2(net221769), .ZN(net221766) );
  NAND2_X4 U4427 ( .A1(n3327), .A2(n3328), .ZN(n3330) );
  INV_X4 U4428 ( .A(net221864), .ZN(n3328) );
  NAND2_X4 U4429 ( .A1(net221875), .A2(net221876), .ZN(net221863) );
  OAI21_X2 U4430 ( .B1(n3324), .B2(net221878), .A(n3325), .ZN(net221876) );
  NAND2_X2 U4431 ( .A1(n3326), .A2(n3322), .ZN(n3325) );
  INV_X4 U4432 ( .A(net221426), .ZN(n3322) );
  NAND2_X2 U4433 ( .A1(n3322), .A2(net221802), .ZN(net221800) );
  NAND2_X4 U4435 ( .A1(net221425), .A2(net221152), .ZN(net221163) );
  NOR2_X1 U4436 ( .A1(net228708), .A2(n8003), .ZN(n3324) );
  INV_X1 U4437 ( .A(net228056), .ZN(net228708) );
  INV_X4 U4438 ( .A(net228940), .ZN(net228056) );
  NAND2_X2 U4439 ( .A1(net221431), .A2(net228056), .ZN(net221812) );
  INV_X16 U4440 ( .A(net228615), .ZN(net228029) );
  NAND2_X4 U4441 ( .A1(net225091), .A2(net228615), .ZN(net223262) );
  INV_X16 U4442 ( .A(net225095), .ZN(net225096) );
  INV_X4 U4443 ( .A(net34717), .ZN(net225095) );
  NOR2_X1 U4444 ( .A1(net34763), .A2(net225091), .ZN(n3331) );
  INV_X16 U4445 ( .A(n3332), .ZN(net225091) );
  INV_X4 U4446 ( .A(net34726), .ZN(n3332) );
  OAI222_X2 U4447 ( .A1(net34613), .A2(net224767), .B1(net224755), .B2(n2735), 
        .C1(net36084), .C2(net34763), .ZN(memWrData[19]) );
  MUX2_X1 U4448 ( .A(net34763), .B(net35052), .S(net224719), .Z(net35483) );
  NAND3_X2 U4449 ( .A1(net227945), .A2(net220714), .A3(net228056), .ZN(
        net228479) );
  NAND2_X2 U4450 ( .A1(net228056), .A2(net229330), .ZN(net228058) );
  INV_X8 U4451 ( .A(net220747), .ZN(net228940) );
  XNOR2_X2 U4452 ( .A(n3333), .B(net220775), .ZN(net220747) );
  XNOR2_X2 U4453 ( .A(net220778), .B(net228715), .ZN(n3333) );
  INV_X32 U4454 ( .A(net224871), .ZN(net224865) );
  INV_X8 U4456 ( .A(net220323), .ZN(net220316) );
  XNOR2_X2 U4458 ( .A(net222158), .B(net224865), .ZN(net222156) );
  NAND2_X2 U4459 ( .A1(n2900), .A2(net228981), .ZN(net228982) );
  AOI22_X2 U4460 ( .A1(net224957), .A2(n2900), .B1(n2702), .B2(n2761), .ZN(
        net223721) );
  NAND3_X2 U4461 ( .A1(n3279), .A2(net223338), .A3(net223339), .ZN(net227823)
         );
  NAND3_X2 U4463 ( .A1(net223339), .A2(net223340), .A3(net223338), .ZN(
        net229624) );
  INV_X8 U4464 ( .A(net222353), .ZN(net225055) );
  INV_X16 U4465 ( .A(net225055), .ZN(net225053) );
  NAND2_X4 U4466 ( .A1(net225581), .A2(n3334), .ZN(net222353) );
  INV_X4 U4467 ( .A(net35047), .ZN(n3334) );
  NAND2_X4 U4468 ( .A1(net225581), .A2(n3334), .ZN(net221648) );
  NAND2_X4 U4469 ( .A1(net225581), .A2(n3334), .ZN(net223437) );
  INV_X4 U4470 ( .A(net225580), .ZN(net225581) );
  NOR3_X4 U4471 ( .A1(n2606), .A2(net228029), .A3(n3336), .ZN(net223347) );
  INV_X2 U4472 ( .A(n3335), .ZN(n3336) );
  INV_X16 U4473 ( .A(net225091), .ZN(net223348) );
  NOR3_X4 U4474 ( .A1(net220315), .A2(net220316), .A3(n3337), .ZN(net220299)
         );
  OAI211_X4 U4475 ( .C1(net220318), .C2(net220319), .A(net220320), .B(n3338), 
        .ZN(n3337) );
  NAND2_X4 U4476 ( .A1(n3344), .A2(n3345), .ZN(net221432) );
  INV_X4 U4477 ( .A(net221820), .ZN(n3343) );
  INV_X4 U4479 ( .A(net221798), .ZN(net221799) );
  INV_X8 U4480 ( .A(net220322), .ZN(net220318) );
  NAND3_X4 U4481 ( .A1(n3341), .A2(n3339), .A3(n2929), .ZN(net220322) );
  INV_X8 U4482 ( .A(n3340), .ZN(n3339) );
  NAND3_X1 U4483 ( .A1(n3341), .A2(n2929), .A3(n3339), .ZN(net230733) );
  NAND2_X4 U4484 ( .A1(net228081), .A2(n3339), .ZN(net220320) );
  INV_X4 U4485 ( .A(net221807), .ZN(net221805) );
  BUF_X4 U4486 ( .A(net221793), .Z(n3341) );
  INV_X8 U4487 ( .A(net220316), .ZN(net229367) );
  NAND2_X4 U4488 ( .A1(net221473), .A2(n3348), .ZN(n3347) );
  NAND4_X2 U4489 ( .A1(n8002), .A2(n3347), .A3(net228768), .A4(net220767), 
        .ZN(net221817) );
  INV_X4 U4490 ( .A(n3347), .ZN(net229270) );
  NAND3_X2 U4491 ( .A1(net220766), .A2(n3347), .A3(net220767), .ZN(net228148)
         );
  INV_X4 U4492 ( .A(n3346), .ZN(n3348) );
  NAND2_X1 U4493 ( .A1(n2604), .A2(n3348), .ZN(net220729) );
  INV_X8 U4495 ( .A(net220889), .ZN(n3346) );
  NOR3_X4 U4496 ( .A1(net221758), .A2(net220644), .A3(n3346), .ZN(net220637)
         );
  INV_X8 U4497 ( .A(net229486), .ZN(net221473) );
  INV_X8 U4498 ( .A(net221473), .ZN(net220851) );
  XNOR2_X2 U4499 ( .A(net222156), .B(net221488), .ZN(net229486) );
  AOI21_X4 U4500 ( .B1(n7988), .B2(n3133), .A(net224873), .ZN(net222745) );
  XNOR2_X2 U4501 ( .A(net224873), .B(n2902), .ZN(net222672) );
  NAND2_X4 U4502 ( .A1(net224873), .A2(net224731), .ZN(net222515) );
  OAI21_X4 U4503 ( .B1(net33205), .B2(n3321), .A(net225622), .ZN(net220524) );
  NAND2_X4 U4504 ( .A1(net225229), .A2(net230143), .ZN(net221652) );
  NAND2_X4 U4505 ( .A1(net224785), .A2(net225102), .ZN(net222698) );
  INV_X16 U4506 ( .A(net225101), .ZN(net225102) );
  INV_X4 U4507 ( .A(net220540), .ZN(net228677) );
  AOI21_X4 U4508 ( .B1(net229575), .B2(net221817), .A(net221890), .ZN(
        net221889) );
  OAI211_X4 U4509 ( .C1(net221888), .C2(net221807), .A(net221889), .B(
        net221416), .ZN(net221875) );
  AND3_X4 U4510 ( .A1(net225601), .A2(net221152), .A3(net225587), .ZN(n3349)
         );
  INV_X8 U4511 ( .A(net220619), .ZN(net225587) );
  XNOR2_X2 U4513 ( .A(net229691), .B(net221905), .ZN(net229291) );
  INV_X4 U4514 ( .A(net221813), .ZN(net221152) );
  INV_X16 U4515 ( .A(net225242), .ZN(net225243) );
  INV_X8 U4516 ( .A(net222771), .ZN(net225242) );
  NAND2_X2 U4517 ( .A1(net225091), .A2(net225096), .ZN(net222771) );
  NAND2_X4 U4518 ( .A1(net221491), .A2(net225029), .ZN(net221488) );
  INV_X8 U4519 ( .A(net221488), .ZN(net221494) );
  INV_X32 U4520 ( .A(net225084), .ZN(net225029) );
  NAND2_X4 U4521 ( .A1(net221817), .A2(net229575), .ZN(net220601) );
  NAND2_X4 U4522 ( .A1(n3353), .A2(n3352), .ZN(net228768) );
  NAND2_X4 U4523 ( .A1(net228149), .A2(n7992), .ZN(net220753) );
  INV_X4 U4524 ( .A(net221924), .ZN(n3352) );
  NOR2_X4 U4525 ( .A1(net221479), .A2(net220640), .ZN(n3353) );
  INV_X8 U4526 ( .A(net220632), .ZN(net220640) );
  INV_X8 U4527 ( .A(n3351), .ZN(net221479) );
  NAND2_X4 U4528 ( .A1(n3356), .A2(n3357), .ZN(n3351) );
  NAND2_X4 U4529 ( .A1(n3354), .A2(n3355), .ZN(n3357) );
  INV_X4 U4530 ( .A(net222370), .ZN(n3354) );
  NAND2_X2 U4531 ( .A1(net222370), .A2(net222371), .ZN(n3356) );
  NAND2_X2 U4532 ( .A1(net229624), .A2(net224737), .ZN(n3702) );
  NOR2_X1 U4534 ( .A1(n7921), .A2(n3126), .ZN(n4883) );
  NAND2_X2 U4535 ( .A1(net221758), .A2(net225587), .ZN(n6150) );
  INV_X1 U4536 ( .A(net225588), .ZN(net228720) );
  NAND2_X2 U4537 ( .A1(n5842), .A2(net221494), .ZN(n3411) );
  NAND2_X4 U4538 ( .A1(n5937), .A2(n7108), .ZN(n5289) );
  OAI211_X4 U4540 ( .C1(n5852), .C2(n3261), .A(n5851), .B(n3947), .ZN(n5853)
         );
  NOR2_X2 U4541 ( .A1(n3386), .A2(n6906), .ZN(n3358) );
  NOR2_X4 U4543 ( .A1(n5420), .A2(n5419), .ZN(n5425) );
  INV_X4 U4544 ( .A(n4718), .ZN(regWrData[7]) );
  NAND2_X4 U4545 ( .A1(n5034), .A2(net224737), .ZN(n3735) );
  NOR2_X2 U4546 ( .A1(n5914), .A2(n2680), .ZN(n5566) );
  NOR2_X1 U4547 ( .A1(n5468), .A2(n3920), .ZN(n5472) );
  INV_X4 U4548 ( .A(n5025), .ZN(n5030) );
  INV_X1 U4549 ( .A(n6588), .ZN(n3361) );
  AOI22_X4 U4550 ( .A1(n3643), .A2(memAddr[10]), .B1(net223245), .B2(n2711), 
        .ZN(n4851) );
  NAND2_X2 U4551 ( .A1(net220663), .A2(n7066), .ZN(n3562) );
  NAND2_X4 U4552 ( .A1(n3362), .A2(n3363), .ZN(n3365) );
  INV_X4 U4553 ( .A(n5820), .ZN(n3362) );
  INV_X4 U4554 ( .A(n5484), .ZN(n3363) );
  NAND2_X1 U4555 ( .A1(n4942), .A2(net224993), .ZN(n3366) );
  NAND2_X1 U4556 ( .A1(\wb/dsize_reg/z2 [15]), .A2(n3934), .ZN(n3367) );
  AND2_X4 U4557 ( .A1(n3366), .A2(n3367), .ZN(n4943) );
  INV_X4 U4558 ( .A(n5816), .ZN(n5820) );
  INV_X4 U4559 ( .A(n6809), .ZN(n7103) );
  NAND2_X1 U4560 ( .A1(n5183), .A2(net230760), .ZN(n3368) );
  NAND2_X1 U4561 ( .A1(n2915), .A2(net224743), .ZN(n3369) );
  INV_X1 U4562 ( .A(net224743), .ZN(net230760) );
  INV_X2 U4563 ( .A(n6141), .ZN(n3483) );
  NAND2_X2 U4565 ( .A1(n2928), .A2(net230157), .ZN(n3371) );
  NAND2_X2 U4566 ( .A1(n4917), .A2(net225214), .ZN(n4921) );
  NOR2_X1 U4568 ( .A1(n3135), .A2(net224955), .ZN(\id_ex/N31 ) );
  OAI22_X1 U4569 ( .A1(n7716), .A2(net224943), .B1(n4683), .B2(n4668), .ZN(
        n7881) );
  OAI221_X1 U4570 ( .B1(n4675), .B2(n6332), .C1(n3135), .C2(n4671), .A(n4661), 
        .ZN(n2123) );
  OAI21_X1 U4571 ( .B1(n4596), .B2(n2757), .A(n4595), .ZN(n4601) );
  AOI21_X1 U4572 ( .B1(n4660), .B2(n3135), .A(n7925), .ZN(n4571) );
  NAND2_X1 U4573 ( .A1(n7709), .A2(n2855), .ZN(n4663) );
  NAND2_X1 U4574 ( .A1(n4551), .A2(n4683), .ZN(n4667) );
  NAND3_X1 U4575 ( .A1(n7710), .A2(n7713), .A3(n7709), .ZN(n4572) );
  INV_X32 U4576 ( .A(net224997), .ZN(net224995) );
  INV_X8 U4577 ( .A(regWrData[22]), .ZN(n5681) );
  OAI211_X4 U4578 ( .C1(n5814), .C2(n6995), .A(n6993), .B(n6994), .ZN(
        net220746) );
  AOI22_X4 U4579 ( .A1(n6987), .A2(n6986), .B1(n6989), .B2(n7059), .ZN(n6994)
         );
  OAI222_X4 U4580 ( .A1(n7575), .A2(net225015), .B1(n2732), .B2(n3933), .C1(
        n2700), .C2(n2792), .ZN(regWrData[22]) );
  INV_X1 U4581 ( .A(n7971), .ZN(n6259) );
  NAND2_X4 U4582 ( .A1(n4228), .A2(n2725), .ZN(n4303) );
  INV_X2 U4583 ( .A(n6865), .ZN(n5192) );
  NAND2_X4 U4584 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  NAND3_X2 U4585 ( .A1(n3204), .A2(n7055), .A3(n3424), .ZN(n3374) );
  NAND2_X2 U4586 ( .A1(n2845), .A2(net223245), .ZN(n3417) );
  OAI21_X1 U4587 ( .B1(n6262), .B2(n3940), .A(n6260), .ZN(n6422) );
  NAND2_X1 U4588 ( .A1(n7296), .A2(n2622), .ZN(n6012) );
  AND3_X4 U4589 ( .A1(n6440), .A2(n6441), .A3(n3375), .ZN(n6444) );
  AND2_X2 U4590 ( .A1(n6442), .A2(n7202), .ZN(n3375) );
  INV_X2 U4591 ( .A(n6440), .ZN(n6448) );
  INV_X2 U4592 ( .A(n6441), .ZN(n6447) );
  AND3_X4 U4593 ( .A1(n6440), .A2(n7202), .A3(n6441), .ZN(n5936) );
  INV_X1 U4594 ( .A(n7030), .ZN(n3376) );
  OAI21_X4 U4595 ( .B1(n7017), .B2(n7016), .A(n7015), .ZN(n7018) );
  NAND4_X1 U4596 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n2135)
         );
  NOR2_X1 U4597 ( .A1(n8012), .A2(n3950), .ZN(n6183) );
  NAND2_X4 U4598 ( .A1(n3604), .A2(n3605), .ZN(net229691) );
  INV_X4 U4599 ( .A(n4396), .ZN(n3553) );
  INV_X2 U4600 ( .A(n7513), .ZN(n4396) );
  INV_X1 U4601 ( .A(n3994), .ZN(n3377) );
  INV_X8 U4602 ( .A(n3881), .ZN(n3882) );
  AOI21_X2 U4603 ( .B1(n3743), .B2(n3942), .A(net225084), .ZN(n5275) );
  OAI21_X1 U4604 ( .B1(n6247), .B2(n3940), .A(n3743), .ZN(n6355) );
  INV_X8 U4605 ( .A(n5507), .ZN(n5428) );
  NOR2_X1 U4606 ( .A1(n2612), .A2(n3010), .ZN(n5233) );
  NAND2_X2 U4607 ( .A1(n6721), .A2(n3242), .ZN(n3526) );
  INV_X4 U4608 ( .A(n3262), .ZN(n4747) );
  NAND2_X2 U4609 ( .A1(n2906), .A2(net228552), .ZN(n3379) );
  INV_X4 U4611 ( .A(net228552), .ZN(net230683) );
  NAND2_X2 U4612 ( .A1(n3592), .A2(net228700), .ZN(n3381) );
  NAND2_X2 U4613 ( .A1(n3380), .A2(net228715), .ZN(n3382) );
  NAND2_X2 U4614 ( .A1(n3381), .A2(n3382), .ZN(n6069) );
  INV_X4 U4615 ( .A(n3592), .ZN(n3380) );
  INV_X1 U4616 ( .A(n3242), .ZN(net228700) );
  NAND2_X4 U4617 ( .A1(n6432), .A2(n6013), .ZN(n5980) );
  XNOR2_X2 U4618 ( .A(n4228), .B(n2725), .ZN(n4231) );
  NOR2_X1 U4619 ( .A1(net225084), .A2(n7990), .ZN(n5314) );
  OAI21_X2 U4620 ( .B1(net225084), .B2(n6071), .A(net224859), .ZN(n6072) );
  AOI21_X2 U4621 ( .B1(n5245), .B2(n3942), .A(net225084), .ZN(n5246) );
  NAND2_X4 U4623 ( .A1(net220889), .A2(net221481), .ZN(net221924) );
  NAND2_X4 U4624 ( .A1(n5138), .A2(n5139), .ZN(n3879) );
  NOR2_X4 U4625 ( .A1(n2781), .A2(n3864), .ZN(n5669) );
  NAND2_X4 U4626 ( .A1(n4279), .A2(n4278), .ZN(n4298) );
  NAND2_X4 U4628 ( .A1(n3796), .A2(net224865), .ZN(n3798) );
  NAND2_X2 U4629 ( .A1(net228949), .A2(net220646), .ZN(n7008) );
  INV_X2 U4630 ( .A(net220644), .ZN(net228949) );
  INV_X8 U4631 ( .A(n3458), .ZN(n3459) );
  INV_X8 U4632 ( .A(n7054), .ZN(n6035) );
  NAND2_X4 U4633 ( .A1(n5130), .A2(n5454), .ZN(n3881) );
  INV_X2 U4634 ( .A(n5184), .ZN(n3384) );
  NAND2_X2 U4635 ( .A1(n4524), .A2(n4298), .ZN(n4300) );
  NOR2_X2 U4636 ( .A1(n7662), .A2(net224895), .ZN(\ex_mem/N53 ) );
  INV_X4 U4637 ( .A(n4062), .ZN(n3518) );
  NAND2_X4 U4638 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  INV_X1 U4639 ( .A(n7514), .ZN(n4013) );
  NOR2_X2 U4640 ( .A1(n6552), .A2(n5892), .ZN(n5900) );
  NAND2_X4 U4641 ( .A1(n3654), .A2(n3655), .ZN(n3657) );
  INV_X4 U4642 ( .A(n6897), .ZN(n3386) );
  INV_X1 U4643 ( .A(n5082), .ZN(n4720) );
  NAND3_X1 U4644 ( .A1(n6879), .A2(n6872), .A3(n6880), .ZN(n6877) );
  NAND2_X2 U4645 ( .A1(n3716), .A2(n2620), .ZN(n3537) );
  OAI22_X2 U4646 ( .A1(n7414), .A2(n3912), .B1(n7701), .B2(n3909), .ZN(n5476)
         );
  INV_X4 U4647 ( .A(n8108), .ZN(n4519) );
  INV_X1 U4648 ( .A(iAddr[4]), .ZN(n4456) );
  NAND4_X4 U4649 ( .A1(n6148), .A2(net229271), .A3(n6147), .A4(net220769), 
        .ZN(n7058) );
  NAND3_X1 U4650 ( .A1(n8004), .A2(n3133), .A3(n6046), .ZN(n6047) );
  NOR2_X1 U4651 ( .A1(net33193), .A2(net224897), .ZN(\ex_mem/N141 ) );
  NAND2_X4 U4652 ( .A1(n5839), .A2(n6151), .ZN(n7112) );
  NOR2_X4 U4653 ( .A1(n3901), .A2(n7414), .ZN(n4888) );
  NAND2_X4 U4654 ( .A1(n6042), .A2(n6985), .ZN(net221807) );
  NAND2_X4 U4655 ( .A1(n3897), .A2(n2990), .ZN(n4124) );
  INV_X4 U4656 ( .A(net228080), .ZN(net228081) );
  INV_X2 U4657 ( .A(n2613), .ZN(net220874) );
  INV_X8 U4658 ( .A(n7288), .ZN(n6586) );
  NAND2_X2 U4659 ( .A1(n2906), .A2(net228552), .ZN(n3388) );
  NAND2_X2 U4660 ( .A1(n3378), .A2(n3388), .ZN(n5053) );
  INV_X1 U4661 ( .A(net224737), .ZN(net228552) );
  NOR2_X2 U4662 ( .A1(n5141), .A2(n6370), .ZN(n5051) );
  NAND2_X2 U4663 ( .A1(n4346), .A2(n4349), .ZN(n4179) );
  NOR2_X1 U4664 ( .A1(n6533), .A2(n6343), .ZN(n6344) );
  INV_X1 U4665 ( .A(n6343), .ZN(n5744) );
  NAND2_X1 U4666 ( .A1(n7358), .A2(n6343), .ZN(n5752) );
  NAND2_X4 U4667 ( .A1(n6748), .A2(n3491), .ZN(n3458) );
  NAND3_X2 U4668 ( .A1(n4942), .A2(n3304), .A3(net224993), .ZN(n4890) );
  NOR2_X2 U4669 ( .A1(n6490), .A2(n6489), .ZN(n6493) );
  XNOR2_X2 U4670 ( .A(n6817), .B(net224859), .ZN(n3389) );
  INV_X4 U4671 ( .A(n3389), .ZN(n5554) );
  INV_X4 U4672 ( .A(n7909), .ZN(n6810) );
  AOI21_X1 U4673 ( .B1(net224843), .B2(n8013), .A(net224835), .ZN(n5753) );
  NAND2_X4 U4674 ( .A1(n3643), .A2(memAddr[13]), .ZN(n5415) );
  NOR2_X1 U4675 ( .A1(n5178), .A2(net224901), .ZN(\ex_mem/N121 ) );
  CLKBUF_X3 U4676 ( .A(n6035), .Z(n3532) );
  NAND3_X4 U4677 ( .A1(n4781), .A2(net224991), .A3(\wb/dsize_reg/z2 [4]), .ZN(
        n4992) );
  NAND2_X2 U4678 ( .A1(n3610), .A2(n6779), .ZN(n3392) );
  NAND2_X2 U4679 ( .A1(n3390), .A2(n3391), .ZN(n3393) );
  INV_X4 U4681 ( .A(n3610), .ZN(n3390) );
  INV_X2 U4683 ( .A(n7223), .ZN(n3395) );
  INV_X2 U4684 ( .A(n5912), .ZN(n5045) );
  NAND2_X1 U4685 ( .A1(n5527), .A2(n5522), .ZN(n3396) );
  INV_X4 U4686 ( .A(n3396), .ZN(n3397) );
  NAND2_X4 U4687 ( .A1(n4510), .A2(n7859), .ZN(n4313) );
  XOR2_X2 U4688 ( .A(n5373), .B(net224861), .Z(n3398) );
  NAND2_X4 U4689 ( .A1(n4931), .A2(memAddr[6]), .ZN(n5097) );
  INV_X8 U4690 ( .A(n7857), .ZN(n3399) );
  INV_X16 U4691 ( .A(n3399), .ZN(iAddr[23]) );
  NAND3_X4 U4692 ( .A1(n8000), .A2(n3412), .A3(net224991), .ZN(n5413) );
  XNOR2_X2 U4693 ( .A(n5205), .B(net224865), .ZN(n3401) );
  INV_X4 U4694 ( .A(n3401), .ZN(n3600) );
  NOR3_X4 U4695 ( .A1(n5165), .A2(n5164), .A3(n5166), .ZN(n3402) );
  NAND3_X4 U4696 ( .A1(n5162), .A2(n5163), .A3(n2637), .ZN(n5164) );
  NOR2_X2 U4697 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND2_X1 U4698 ( .A1(n6373), .A2(net221481), .ZN(n6374) );
  NAND2_X4 U4699 ( .A1(net223245), .A2(n2869), .ZN(n5081) );
  OAI21_X2 U4700 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(n6754) );
  NAND2_X4 U4701 ( .A1(n6749), .A2(n3459), .ZN(n6010) );
  NOR2_X1 U4702 ( .A1(n7180), .A2(n3196), .ZN(n7187) );
  NAND2_X2 U4703 ( .A1(n2859), .A2(net229656), .ZN(n3403) );
  OAI21_X1 U4704 ( .B1(n6689), .B2(n6688), .A(n6687), .ZN(n6690) );
  INV_X8 U4705 ( .A(n6688), .ZN(n6683) );
  INV_X4 U4706 ( .A(n5504), .ZN(n3476) );
  NAND2_X4 U4707 ( .A1(n6400), .A2(n5384), .ZN(n5385) );
  INV_X8 U4708 ( .A(n6676), .ZN(n6677) );
  INV_X1 U4709 ( .A(n3846), .ZN(n7060) );
  INV_X2 U4710 ( .A(n5490), .ZN(n5491) );
  NAND2_X4 U4711 ( .A1(n7987), .A2(n5893), .ZN(n5890) );
  INV_X4 U4712 ( .A(net221758), .ZN(net229005) );
  NAND2_X4 U4713 ( .A1(n6866), .A2(n6867), .ZN(n6869) );
  NAND2_X4 U4714 ( .A1(n3425), .A2(n5503), .ZN(n3478) );
  INV_X4 U4715 ( .A(n5508), .ZN(n3439) );
  NAND2_X4 U4717 ( .A1(net225237), .A2(n2979), .ZN(n5387) );
  NAND2_X2 U4718 ( .A1(n5668), .A2(net225047), .ZN(n5671) );
  AOI21_X4 U4719 ( .B1(n6260), .B2(n3942), .A(net225084), .ZN(n5672) );
  NAND4_X4 U4720 ( .A1(n5427), .A2(n5425), .A3(n5426), .A4(n5424), .ZN(n5507)
         );
  NOR2_X4 U4721 ( .A1(n5408), .A2(n5407), .ZN(n5412) );
  NAND2_X4 U4722 ( .A1(n3525), .A2(n3272), .ZN(n3527) );
  NAND2_X2 U4723 ( .A1(n5113), .A2(net230493), .ZN(n3404) );
  NAND2_X2 U4724 ( .A1(n2897), .A2(net230088), .ZN(n3405) );
  NAND2_X4 U4725 ( .A1(n3404), .A2(n3405), .ZN(n5187) );
  INV_X4 U4726 ( .A(net230088), .ZN(net230493) );
  NAND2_X2 U4727 ( .A1(n5111), .A2(n5112), .ZN(n5113) );
  INV_X32 U4728 ( .A(net225017), .ZN(net225015) );
  NOR2_X4 U4729 ( .A1(net225015), .A2(n5387), .ZN(n5379) );
  INV_X8 U4730 ( .A(net225015), .ZN(net225013) );
  INV_X1 U4731 ( .A(net230611), .ZN(net230488) );
  NAND2_X4 U4732 ( .A1(net220894), .A2(n6881), .ZN(n3639) );
  NOR2_X4 U4733 ( .A1(n6899), .A2(n6900), .ZN(n6901) );
  NAND2_X4 U4734 ( .A1(n5088), .A2(n5087), .ZN(n5311) );
  NAND3_X2 U4735 ( .A1(reg31Val_0[7]), .A2(net228359), .A3(net230143), .ZN(
        n5087) );
  NAND3_X1 U4736 ( .A1(n5073), .A2(net224731), .A3(n5072), .ZN(n5077) );
  NAND2_X2 U4737 ( .A1(n3569), .A2(net230181), .ZN(n3492) );
  NAND2_X4 U4738 ( .A1(n3415), .A2(n6936), .ZN(n6937) );
  INV_X1 U4739 ( .A(n5902), .ZN(n3406) );
  NOR2_X2 U4740 ( .A1(n4258), .A2(n4259), .ZN(n4265) );
  INV_X4 U4741 ( .A(n5976), .ZN(n3884) );
  NAND2_X2 U4742 ( .A1(n5967), .A2(n3768), .ZN(n5859) );
  NAND2_X2 U4743 ( .A1(net224865), .A2(n6167), .ZN(n3409) );
  INV_X8 U4745 ( .A(n6829), .ZN(n5893) );
  OAI222_X4 U4746 ( .A1(n3935), .A2(n2950), .B1(n2728), .B2(n3933), .C1(n7546), 
        .C2(n3253), .ZN(regWrData[20]) );
  NAND2_X1 U4747 ( .A1(n3552), .A2(n2778), .ZN(n4399) );
  NAND2_X1 U4748 ( .A1(n7438), .A2(n3247), .ZN(n4120) );
  NAND4_X2 U4749 ( .A1(n5434), .A2(n7970), .A3(n3658), .A4(n5433), .ZN(n3413)
         );
  NAND4_X2 U4750 ( .A1(n5434), .A2(n7970), .A3(n3658), .A4(n5433), .ZN(n6153)
         );
  NAND2_X4 U4751 ( .A1(n6058), .A2(net229239), .ZN(n3659) );
  NAND2_X4 U4752 ( .A1(n4981), .A2(n4990), .ZN(n4985) );
  XOR2_X2 U4753 ( .A(n6047), .B(net224859), .Z(n3789) );
  NAND2_X4 U4755 ( .A1(n6462), .A2(n6126), .ZN(n6935) );
  NAND2_X4 U4756 ( .A1(n5438), .A2(n5437), .ZN(n5098) );
  INV_X1 U4757 ( .A(n2673), .ZN(n4806) );
  NAND2_X4 U4759 ( .A1(n5118), .A2(net225047), .ZN(n5344) );
  NAND3_X2 U4760 ( .A1(n6044), .A2(n6043), .A3(n5647), .ZN(n3416) );
  NAND2_X2 U4761 ( .A1(net228058), .A2(n6644), .ZN(n6650) );
  XNOR2_X2 U4762 ( .A(n6817), .B(net224861), .ZN(n5367) );
  OR2_X4 U4763 ( .A1(n5093), .A2(n7533), .ZN(n3418) );
  NAND2_X4 U4764 ( .A1(n3417), .A2(n3418), .ZN(n4774) );
  OAI21_X4 U4765 ( .B1(n6952), .B2(n6953), .A(n7169), .ZN(n6960) );
  AOI22_X2 U4766 ( .A1(net223245), .A2(n2712), .B1(n3643), .B2(memAddr[24]), 
        .ZN(n4752) );
  NOR2_X4 U4768 ( .A1(n2784), .A2(n3864), .ZN(n6090) );
  INV_X1 U4769 ( .A(iAddr[24]), .ZN(n4512) );
  NAND2_X4 U4770 ( .A1(n5669), .A2(net225047), .ZN(n5670) );
  INV_X2 U4771 ( .A(n3309), .ZN(n6867) );
  XNOR2_X2 U4772 ( .A(n6421), .B(n3226), .ZN(n3567) );
  NAND2_X1 U4773 ( .A1(n6213), .A2(n6212), .ZN(n6218) );
  NAND2_X1 U4774 ( .A1(n6215), .A2(n6213), .ZN(n5248) );
  NAND2_X2 U4775 ( .A1(n2764), .A2(net229782), .ZN(n3420) );
  NAND2_X2 U4776 ( .A1(n5937), .A2(n3421), .ZN(n3422) );
  NAND2_X4 U4777 ( .A1(n3422), .A2(n6464), .ZN(n6468) );
  INV_X4 U4778 ( .A(n6465), .ZN(n3421) );
  INV_X1 U4779 ( .A(net224735), .ZN(net229782) );
  NOR2_X4 U4781 ( .A1(n6468), .A2(n6467), .ZN(n6474) );
  INV_X4 U4782 ( .A(n3494), .ZN(n5143) );
  NOR2_X4 U4783 ( .A1(net225238), .A2(n3651), .ZN(n4765) );
  INV_X1 U4784 ( .A(n6152), .ZN(n3423) );
  INV_X2 U4785 ( .A(n3423), .ZN(n3424) );
  XNOR2_X2 U4786 ( .A(n5497), .B(net228323), .ZN(n3425) );
  INV_X8 U4787 ( .A(n4925), .ZN(n3904) );
  NAND2_X1 U4788 ( .A1(n3916), .A2(n6583), .ZN(n3427) );
  AND3_X4 U4789 ( .A1(n5051), .A2(n5777), .A3(n3215), .ZN(n3871) );
  INV_X8 U4790 ( .A(n5665), .ZN(n5937) );
  INV_X8 U4791 ( .A(regWrData[15]), .ZN(n5481) );
  NAND3_X4 U4793 ( .A1(n4945), .A2(n4944), .A3(n4943), .ZN(regWrData[15]) );
  NAND3_X4 U4794 ( .A1(n3814), .A2(n6884), .A3(n6146), .ZN(n7059) );
  AOI21_X2 U4795 ( .B1(n7061), .B2(n3652), .A(n7059), .ZN(n7063) );
  INV_X8 U4796 ( .A(n7059), .ZN(n6149) );
  INV_X4 U4797 ( .A(n6411), .ZN(n3429) );
  AOI211_X4 U4798 ( .C1(n6400), .C2(n6399), .A(n6398), .B(n6397), .ZN(n6403)
         );
  INV_X8 U4799 ( .A(n6918), .ZN(n6919) );
  NAND2_X1 U4800 ( .A1(n6595), .A2(n3361), .ZN(n6596) );
  INV_X8 U4801 ( .A(n6825), .ZN(n6588) );
  XNOR2_X2 U4802 ( .A(n4362), .B(iAddr[31]), .ZN(n3432) );
  INV_X4 U4803 ( .A(n4541), .ZN(iAddr[29]) );
  OAI22_X2 U4804 ( .A1(n7459), .A2(n7508), .B1(n3139), .B2(n4246), .ZN(n3434)
         );
  OAI221_X1 U4805 ( .B1(n4233), .B2(n4184), .C1(n3150), .C2(n4177), .A(n4187), 
        .ZN(n3435) );
  INV_X2 U4806 ( .A(n7906), .ZN(n4541) );
  NOR2_X4 U4807 ( .A1(n5410), .A2(n3465), .ZN(n5411) );
  NAND2_X4 U4808 ( .A1(n5881), .A2(n3807), .ZN(\ex_mem/N216 ) );
  AOI21_X4 U4809 ( .B1(n3891), .B2(n7201), .A(n5954), .ZN(n5955) );
  NOR2_X2 U4810 ( .A1(net225230), .A2(n7543), .ZN(n3555) );
  NOR2_X1 U4811 ( .A1(n7578), .A2(n3290), .ZN(n5242) );
  NAND2_X2 U4813 ( .A1(n3819), .A2(n3820), .ZN(n6548) );
  NAND3_X1 U4814 ( .A1(n3795), .A2(\wb/dsize_reg/z2 [24]), .A3(net225045), 
        .ZN(n6213) );
  NAND3_X4 U4816 ( .A1(n5159), .A2(n5158), .A3(n3437), .ZN(n5165) );
  INV_X4 U4817 ( .A(n3436), .ZN(n3437) );
  NAND4_X2 U4818 ( .A1(n4323), .A2(n4349), .A3(n4322), .A4(n4321), .ZN(n4324)
         );
  INV_X4 U4819 ( .A(n6950), .ZN(n6953) );
  AND3_X4 U4820 ( .A1(n6068), .A2(n6015), .A3(net225605), .ZN(n3872) );
  OAI21_X4 U4821 ( .B1(n3689), .B2(n6688), .A(n6824), .ZN(n5459) );
  INV_X2 U4822 ( .A(n6895), .ZN(n6896) );
  INV_X8 U4823 ( .A(net220728), .ZN(net220644) );
  NAND2_X2 U4824 ( .A1(n5570), .A2(net224861), .ZN(n3670) );
  NAND2_X2 U4825 ( .A1(n5914), .A2(n2680), .ZN(n3441) );
  NAND2_X4 U4826 ( .A1(n3439), .A2(n3440), .ZN(n3442) );
  NAND2_X4 U4827 ( .A1(n3441), .A2(n3442), .ZN(n5509) );
  OR2_X2 U4828 ( .A1(n4880), .A2(net224999), .ZN(n3443) );
  NAND3_X2 U4829 ( .A1(n3443), .A2(n3444), .A3(n4878), .ZN(n5468) );
  INV_X8 U4830 ( .A(n5509), .ZN(n5911) );
  NOR2_X4 U4831 ( .A1(n6549), .A2(n6552), .ZN(n5899) );
  NOR2_X4 U4832 ( .A1(n8011), .A2(net224871), .ZN(n5319) );
  NAND3_X2 U4834 ( .A1(n4776), .A2(net225237), .A3(net224991), .ZN(n5074) );
  NAND2_X4 U4835 ( .A1(n4991), .A2(n5567), .ZN(n6796) );
  NAND2_X4 U4836 ( .A1(net220885), .A2(n6884), .ZN(n3453) );
  INV_X4 U4837 ( .A(n7342), .ZN(n6913) );
  NOR2_X2 U4838 ( .A1(n5439), .A2(net224745), .ZN(n5442) );
  NAND2_X2 U4839 ( .A1(n5096), .A2(n3901), .ZN(n5439) );
  INV_X4 U4840 ( .A(n3455), .ZN(n3445) );
  OAI22_X4 U4841 ( .A1(n3935), .A2(n4898), .B1(n3252), .B2(n4897), .ZN(n4899)
         );
  INV_X8 U4842 ( .A(n4899), .ZN(n5773) );
  NOR2_X2 U4843 ( .A1(n6990), .A2(net220753), .ZN(n6992) );
  NAND2_X4 U4844 ( .A1(n7941), .A2(n7218), .ZN(n6669) );
  INV_X2 U4845 ( .A(n4868), .ZN(n3505) );
  NAND2_X1 U4846 ( .A1(net224871), .A2(n5330), .ZN(n3447) );
  NAND2_X2 U4847 ( .A1(net224865), .A2(n3446), .ZN(n3448) );
  NAND2_X2 U4848 ( .A1(n3447), .A2(n3448), .ZN(n5339) );
  INV_X4 U4849 ( .A(n5330), .ZN(n3446) );
  OAI21_X4 U4850 ( .B1(net33205), .B2(n3321), .A(net225622), .ZN(n3449) );
  NAND2_X4 U4851 ( .A1(n5339), .A2(n5331), .ZN(n5457) );
  NAND2_X4 U4852 ( .A1(n5891), .A2(n3284), .ZN(n3548) );
  NAND2_X4 U4853 ( .A1(n3451), .A2(n2603), .ZN(n4984) );
  INV_X4 U4854 ( .A(n4983), .ZN(n3450) );
  NAND2_X1 U4855 ( .A1(net220885), .A2(n6884), .ZN(n3452) );
  NAND2_X4 U4856 ( .A1(net220656), .A2(net221881), .ZN(n6884) );
  NAND2_X4 U4857 ( .A1(n3862), .A2(n6191), .ZN(n6197) );
  OAI211_X2 U4858 ( .C1(n3815), .C2(n3261), .A(n6184), .B(n3947), .ZN(n6187)
         );
  NOR2_X2 U4859 ( .A1(n7193), .A2(n6461), .ZN(n5934) );
  NAND3_X2 U4860 ( .A1(n5761), .A2(n5969), .A3(n5760), .ZN(n3454) );
  NAND2_X4 U4861 ( .A1(n6048), .A2(net230493), .ZN(n3456) );
  NAND2_X2 U4862 ( .A1(n2773), .A2(net229522), .ZN(n3457) );
  NAND2_X4 U4863 ( .A1(n3456), .A2(n3457), .ZN(n6066) );
  INV_X1 U4864 ( .A(net224733), .ZN(net229522) );
  INV_X4 U4865 ( .A(n5526), .ZN(n5529) );
  INV_X1 U4866 ( .A(net224735), .ZN(net229784) );
  INV_X8 U4867 ( .A(n5013), .ZN(n5014) );
  XNOR2_X2 U4868 ( .A(n3606), .B(net224865), .ZN(n6039) );
  NAND2_X4 U4869 ( .A1(net223245), .A2(n2743), .ZN(n5034) );
  NOR2_X1 U4870 ( .A1(n4747), .A2(net224899), .ZN(\ex_mem/N122 ) );
  NAND2_X2 U4871 ( .A1(n7965), .A2(n3304), .ZN(n5490) );
  NAND2_X4 U4872 ( .A1(n3463), .A2(n5411), .ZN(n5427) );
  INV_X4 U4873 ( .A(n3462), .ZN(n3463) );
  NOR2_X4 U4874 ( .A1(n2584), .A2(net224743), .ZN(n3464) );
  INV_X4 U4875 ( .A(n3464), .ZN(n3465) );
  INV_X4 U4876 ( .A(net224861), .ZN(net227791) );
  NAND2_X2 U4877 ( .A1(n5323), .A2(n3746), .ZN(n5085) );
  NAND3_X2 U4878 ( .A1(n4302), .A2(n4291), .A3(n4520), .ZN(n4023) );
  NAND2_X2 U4879 ( .A1(n4782), .A2(net225047), .ZN(n4783) );
  BUF_X32 U4880 ( .A(n5145), .Z(n3467) );
  NAND3_X4 U4881 ( .A1(n5495), .A2(n5494), .A3(n5496), .ZN(n5497) );
  NAND2_X1 U4882 ( .A1(net224865), .A2(n5477), .ZN(n5475) );
  OAI211_X1 U4883 ( .C1(n3945), .C2(n6070), .A(net224865), .B(n3133), .ZN(
        n6073) );
  NAND2_X2 U4885 ( .A1(n3469), .A2(n2683), .ZN(n4769) );
  INV_X4 U4886 ( .A(n3468), .ZN(n3469) );
  BUF_X32 U4887 ( .A(n5146), .Z(n3470) );
  NAND2_X4 U4888 ( .A1(n5118), .A2(net225214), .ZN(n5338) );
  INV_X8 U4889 ( .A(n3884), .ZN(n3885) );
  NAND2_X4 U4890 ( .A1(n3471), .A2(n3472), .ZN(n3474) );
  NAND2_X4 U4891 ( .A1(n3473), .A2(n3474), .ZN(n6598) );
  INV_X4 U4892 ( .A(n5453), .ZN(n3471) );
  NOR2_X4 U4893 ( .A1(n5193), .A2(n5192), .ZN(n5195) );
  INV_X1 U4894 ( .A(n5066), .ZN(n3475) );
  NAND2_X4 U4895 ( .A1(n3476), .A2(n3477), .ZN(n3479) );
  NAND2_X4 U4896 ( .A1(n3478), .A2(n3479), .ZN(n6714) );
  INV_X16 U4897 ( .A(n5693), .ZN(n3934) );
  NAND2_X4 U4898 ( .A1(n3785), .A2(net230143), .ZN(n5693) );
  INV_X4 U4899 ( .A(net220315), .ZN(net230231) );
  INV_X8 U4900 ( .A(n3268), .ZN(net220315) );
  AND3_X2 U4901 ( .A1(n5937), .A2(n6944), .A3(n6683), .ZN(n3521) );
  INV_X1 U4902 ( .A(net221165), .ZN(net230225) );
  INV_X2 U4903 ( .A(net230225), .ZN(net230226) );
  NAND2_X2 U4904 ( .A1(n2586), .A2(n5793), .ZN(n3480) );
  NAND2_X4 U4905 ( .A1(n3480), .A2(n3481), .ZN(n6733) );
  INV_X4 U4906 ( .A(n3483), .ZN(n3484) );
  NAND2_X2 U4907 ( .A1(n6713), .A2(n6712), .ZN(n6715) );
  BUF_X8 U4908 ( .A(n3249), .Z(n3539) );
  INV_X8 U4909 ( .A(n2588), .ZN(n3485) );
  NOR2_X2 U4910 ( .A1(net225238), .A2(n2792), .ZN(n4734) );
  NAND3_X4 U4911 ( .A1(n3826), .A2(n3771), .A3(net224993), .ZN(n5220) );
  NAND2_X2 U4912 ( .A1(net224865), .A2(net222155), .ZN(n3486) );
  NAND2_X4 U4913 ( .A1(n3242), .A2(net230199), .ZN(n3487) );
  NAND2_X4 U4914 ( .A1(n3486), .A2(n3487), .ZN(n5842) );
  NAND3_X2 U4915 ( .A1(n3859), .A2(\wb/dsize_reg/z2 [16]), .A3(net225045), 
        .ZN(n6212) );
  NAND2_X2 U4916 ( .A1(net229370), .A2(n5049), .ZN(n3640) );
  NAND2_X2 U4917 ( .A1(net224993), .A2(n5008), .ZN(n3509) );
  NAND2_X1 U4918 ( .A1(net224861), .A2(n6185), .ZN(n3489) );
  NAND2_X4 U4919 ( .A1(net230191), .A2(n3488), .ZN(n3490) );
  INV_X1 U4920 ( .A(net224861), .ZN(net230191) );
  INV_X4 U4921 ( .A(n6185), .ZN(n3488) );
  INV_X2 U4922 ( .A(n5505), .ZN(n3817) );
  NAND2_X4 U4923 ( .A1(n5574), .A2(n5573), .ZN(n3491) );
  INV_X8 U4924 ( .A(n5796), .ZN(n6034) );
  NAND3_X2 U4925 ( .A1(n4882), .A2(n4881), .A3(net224993), .ZN(n4885) );
  NAND2_X2 U4926 ( .A1(n2901), .A2(net227828), .ZN(n3493) );
  INV_X4 U4927 ( .A(net227828), .ZN(net230181) );
  INV_X1 U4928 ( .A(net224737), .ZN(net227828) );
  NAND3_X2 U4929 ( .A1(n4904), .A2(n4905), .A3(n4906), .ZN(n3569) );
  INV_X1 U4930 ( .A(n6790), .ZN(n3724) );
  INV_X1 U4931 ( .A(n3724), .ZN(n3725) );
  NAND2_X4 U4932 ( .A1(n4088), .A2(n4081), .ZN(n4098) );
  XNOR2_X2 U4933 ( .A(n4335), .B(n2920), .ZN(n4087) );
  NAND2_X2 U4934 ( .A1(n8005), .A2(n7021), .ZN(n7015) );
  MUX2_X2 U4935 ( .A(n5203), .B(n2763), .S(net229173), .Z(n3494) );
  AOI21_X2 U4936 ( .B1(n4240), .B2(n7931), .A(n3603), .ZN(n4241) );
  NAND2_X4 U4938 ( .A1(n2613), .A2(n6142), .ZN(n6888) );
  AOI21_X2 U4939 ( .B1(n7181), .B2(n5608), .A(n3242), .ZN(n5609) );
  NAND2_X2 U4940 ( .A1(n2773), .A2(net228345), .ZN(n3498) );
  NAND2_X4 U4941 ( .A1(n3497), .A2(n3498), .ZN(n5198) );
  INV_X1 U4942 ( .A(net224737), .ZN(net228345) );
  INV_X8 U4943 ( .A(net223437), .ZN(net230142) );
  INV_X16 U4944 ( .A(net230144), .ZN(net230145) );
  INV_X1 U4945 ( .A(n3549), .ZN(n6399) );
  NAND4_X4 U4946 ( .A1(n4181), .A2(n4180), .A3(n4323), .A4(n4198), .ZN(n4189)
         );
  NAND2_X4 U4947 ( .A1(n4190), .A2(n4189), .ZN(n4195) );
  MUX2_X2 U4948 ( .A(n4747), .B(n7736), .S(net230157), .Z(n3499) );
  OAI21_X4 U4949 ( .B1(n5077), .B2(n5076), .A(n6811), .ZN(n5366) );
  NAND2_X2 U4950 ( .A1(n5040), .A2(net230130), .ZN(n3500) );
  NAND2_X2 U4951 ( .A1(n2913), .A2(net229958), .ZN(n3501) );
  NAND2_X4 U4952 ( .A1(n3500), .A2(n3501), .ZN(n5041) );
  INV_X1 U4953 ( .A(net229958), .ZN(net230130) );
  INV_X1 U4954 ( .A(net224737), .ZN(net229958) );
  NOR2_X1 U4955 ( .A1(n2576), .A2(n3950), .ZN(n6654) );
  NAND2_X4 U4956 ( .A1(n3503), .A2(n3504), .ZN(n6829) );
  CLKBUF_X3 U4957 ( .A(n6829), .Z(n3683) );
  NAND2_X2 U4958 ( .A1(net223245), .A2(n2748), .ZN(n4986) );
  NAND2_X2 U4959 ( .A1(n2917), .A2(net230103), .ZN(n3506) );
  NAND2_X1 U4960 ( .A1(n5049), .A2(net224733), .ZN(n3507) );
  INV_X1 U4961 ( .A(net224733), .ZN(net230103) );
  OAI21_X1 U4962 ( .B1(n6725), .B2(n3918), .A(n6574), .ZN(n6575) );
  OAI21_X1 U4963 ( .B1(n6725), .B2(n2701), .A(n6724), .ZN(n6726) );
  INV_X1 U4964 ( .A(iAddr[28]), .ZN(n4535) );
  NAND2_X1 U4965 ( .A1(n7176), .A2(n5835), .ZN(n5788) );
  AOI22_X2 U4966 ( .A1(n6661), .A2(n5835), .B1(n5860), .B2(n3955), .ZN(n5728)
         );
  INV_X4 U4967 ( .A(n3509), .ZN(n3510) );
  INV_X2 U4968 ( .A(n6934), .ZN(n3768) );
  OAI221_X4 U4969 ( .B1(n7430), .B2(n4465), .C1(n4133), .C2(n3895), .A(n4132), 
        .ZN(iAddr[4]) );
  NAND2_X4 U4970 ( .A1(net229330), .A2(n6639), .ZN(n6641) );
  INV_X8 U4971 ( .A(n7908), .ZN(n5641) );
  NAND3_X2 U4972 ( .A1(iAddr[9]), .A2(iAddr[12]), .A3(iAddr[13]), .ZN(n4330)
         );
  NAND2_X4 U4974 ( .A1(n3513), .A2(n3514), .ZN(n3689) );
  AOI21_X1 U4976 ( .B1(n6684), .B2(n2838), .A(n2632), .ZN(n6691) );
  AOI21_X1 U4977 ( .B1(net224843), .B2(n2632), .A(net224835), .ZN(n6689) );
  NAND2_X4 U4978 ( .A1(n6685), .A2(n6741), .ZN(n3667) );
  INV_X2 U4979 ( .A(n7341), .ZN(n7343) );
  NAND2_X4 U4980 ( .A1(n8003), .A2(n6915), .ZN(n6918) );
  NAND2_X4 U4981 ( .A1(n2978), .A2(n3515), .ZN(n3516) );
  NAND2_X4 U4982 ( .A1(n3516), .A2(n5446), .ZN(n5448) );
  INV_X4 U4983 ( .A(n5447), .ZN(n3515) );
  NAND3_X2 U4984 ( .A1(n5440), .A2(n5442), .A3(n5441), .ZN(n5447) );
  NOR2_X1 U4985 ( .A1(n6485), .A2(n6342), .ZN(n6346) );
  NAND4_X2 U4986 ( .A1(n5235), .A2(n5441), .A3(n5437), .A4(n2581), .ZN(n5238)
         );
  INV_X4 U4987 ( .A(n3714), .ZN(n3715) );
  INV_X1 U4988 ( .A(n2674), .ZN(n4767) );
  NOR3_X2 U4989 ( .A1(n3905), .A2(n7575), .A3(net225238), .ZN(n4735) );
  NAND2_X4 U4990 ( .A1(n3518), .A2(n4250), .ZN(n3520) );
  NAND2_X4 U4991 ( .A1(n3519), .A2(n3520), .ZN(n4066) );
  NOR2_X2 U4992 ( .A1(n4780), .A2(net224903), .ZN(\ex_mem/N108 ) );
  AOI21_X1 U4993 ( .B1(net224843), .B2(n6814), .A(net224835), .ZN(n6818) );
  AOI21_X2 U4994 ( .B1(n6813), .B2(n2838), .A(n6814), .ZN(n6820) );
  BUF_X32 U4995 ( .A(n6812), .Z(n3696) );
  INV_X8 U4996 ( .A(n4503), .ZN(n4492) );
  NAND2_X4 U4997 ( .A1(n3665), .A2(n3661), .ZN(net221878) );
  XNOR2_X2 U4998 ( .A(n3523), .B(net224859), .ZN(n5582) );
  NAND2_X4 U4999 ( .A1(net221431), .A2(n6639), .ZN(n6115) );
  INV_X8 U5000 ( .A(net220895), .ZN(net220894) );
  INV_X1 U5001 ( .A(n6526), .ZN(n3697) );
  NOR2_X2 U5002 ( .A1(n5600), .A2(n5599), .ZN(n5607) );
  NAND2_X4 U5004 ( .A1(n5405), .A2(n5406), .ZN(n3524) );
  NAND2_X2 U5005 ( .A1(n5405), .A2(n5406), .ZN(n5506) );
  NAND2_X2 U5006 ( .A1(n4802), .A2(n3867), .ZN(n4846) );
  INV_X2 U5007 ( .A(n6335), .ZN(n5787) );
  NAND2_X1 U5008 ( .A1(n7358), .A2(n6335), .ZN(n5827) );
  MUX2_X2 U5009 ( .A(n3750), .B(n2915), .S(net224743), .Z(n3854) );
  NAND2_X2 U5010 ( .A1(n7219), .A2(n6663), .ZN(n3528) );
  NAND2_X1 U5011 ( .A1(n7255), .A2(n7205), .ZN(n3529) );
  NAND2_X4 U5012 ( .A1(n3528), .A2(n3529), .ZN(n7220) );
  NAND2_X1 U5013 ( .A1(n7218), .A2(n7941), .ZN(n7219) );
  INV_X8 U5014 ( .A(n7193), .ZN(n7255) );
  NAND3_X2 U5015 ( .A1(n7256), .A2(n3922), .A3(n3955), .ZN(n7257) );
  INV_X4 U5016 ( .A(n7432), .ZN(n3530) );
  NOR2_X2 U5017 ( .A1(net221874), .A2(n5079), .ZN(n5106) );
  NAND3_X2 U5019 ( .A1(n6403), .A2(n6402), .A3(n3540), .ZN(n6868) );
  INV_X8 U5020 ( .A(net225587), .ZN(net225588) );
  NAND2_X2 U5022 ( .A1(n5451), .A2(n6823), .ZN(n5450) );
  BUF_X8 U5023 ( .A(n6780), .Z(n3610) );
  NAND2_X4 U5024 ( .A1(n3548), .A2(n3615), .ZN(n5796) );
  BUF_X32 U5025 ( .A(n3558), .Z(n3533) );
  NAND2_X4 U5027 ( .A1(n5582), .A2(n3773), .ZN(n6678) );
  INV_X4 U5028 ( .A(n6914), .ZN(n6925) );
  INV_X8 U5029 ( .A(n3524), .ZN(n5429) );
  NAND2_X4 U5030 ( .A1(n5381), .A2(n5380), .ZN(n5395) );
  NOR2_X2 U5031 ( .A1(n2700), .A2(n5386), .ZN(n5377) );
  NAND2_X4 U5033 ( .A1(net224943), .A2(n7556), .ZN(n7884) );
  NAND3_X2 U5034 ( .A1(net228018), .A2(n2760), .A3(net228029), .ZN(n5096) );
  OAI21_X1 U5035 ( .B1(n2694), .B2(net224851), .A(n2838), .ZN(n6719) );
  INV_X1 U5036 ( .A(n2629), .ZN(net229952) );
  INV_X4 U5037 ( .A(n5892), .ZN(n3534) );
  INV_X2 U5038 ( .A(n5891), .ZN(n5892) );
  NOR3_X2 U5039 ( .A1(n3903), .A2(n2951), .A3(n3175), .ZN(n4766) );
  INV_X1 U5040 ( .A(n3285), .ZN(n3535) );
  NAND2_X4 U5041 ( .A1(n3536), .A2(n3709), .ZN(n3538) );
  INV_X4 U5042 ( .A(n6652), .ZN(n3536) );
  NAND2_X4 U5043 ( .A1(n5356), .A2(\wb/dsize_reg/z2 [28]), .ZN(n4834) );
  INV_X1 U5044 ( .A(n6634), .ZN(n3540) );
  INV_X4 U5045 ( .A(n3540), .ZN(n3541) );
  NAND2_X4 U5046 ( .A1(n4837), .A2(n4838), .ZN(n5027) );
  INV_X16 U5047 ( .A(n3910), .ZN(n3912) );
  INV_X4 U5048 ( .A(n5571), .ZN(n5620) );
  INV_X8 U5049 ( .A(net225102), .ZN(net223209) );
  INV_X1 U5050 ( .A(n7947), .ZN(n3543) );
  INV_X4 U5051 ( .A(n3543), .ZN(n3544) );
  NAND2_X4 U5052 ( .A1(net221152), .A2(net221153), .ZN(n6984) );
  NOR2_X2 U5054 ( .A1(n5890), .A2(n5889), .ZN(n5901) );
  NAND2_X4 U5055 ( .A1(n6699), .A2(n6698), .ZN(n6700) );
  NAND2_X4 U5056 ( .A1(n6010), .A2(n3554), .ZN(n6679) );
  NAND2_X1 U5057 ( .A1(n5403), .A2(n5404), .ZN(regWrData[13]) );
  NAND3_X1 U5058 ( .A1(n5667), .A2(n3898), .A3(net225214), .ZN(n4863) );
  BUF_X32 U5059 ( .A(n3825), .Z(n3547) );
  NOR2_X4 U5060 ( .A1(net225238), .A2(n3556), .ZN(n4893) );
  NAND2_X4 U5061 ( .A1(n6124), .A2(n7027), .ZN(n6955) );
  INV_X8 U5062 ( .A(n5231), .ZN(n6124) );
  NAND2_X4 U5063 ( .A1(n3643), .A2(memAddr[1]), .ZN(n4973) );
  NAND2_X4 U5064 ( .A1(n5598), .A2(n6772), .ZN(n6748) );
  AOI22_X4 U5065 ( .A1(n7747), .A2(net224745), .B1(n7993), .B2(net224737), 
        .ZN(n5060) );
  XNOR2_X1 U5066 ( .A(net224869), .B(n2898), .ZN(n6396) );
  INV_X2 U5067 ( .A(n5566), .ZN(n7141) );
  NOR2_X4 U5068 ( .A1(n6038), .A2(n3645), .ZN(n5042) );
  NOR2_X4 U5070 ( .A1(net229307), .A2(net224783), .ZN(n4848) );
  INV_X4 U5071 ( .A(n7553), .ZN(n4802) );
  AND3_X4 U5073 ( .A1(reg31Val_0[29]), .A2(net225237), .A3(net224781), .ZN(
        n3550) );
  NOR2_X4 U5074 ( .A1(n3965), .A2(n3146), .ZN(n3552) );
  AOI21_X2 U5075 ( .B1(n3491), .B2(n6751), .A(n5633), .ZN(n3554) );
  NAND3_X2 U5076 ( .A1(n6215), .A2(n6216), .A3(n6214), .ZN(n5600) );
  NAND2_X4 U5077 ( .A1(net221758), .A2(net225587), .ZN(n3814) );
  INV_X1 U5078 ( .A(n6810), .ZN(n3557) );
  INV_X1 U5079 ( .A(n4519), .ZN(n3790) );
  INV_X1 U5080 ( .A(n3180), .ZN(n4121) );
  NAND3_X2 U5082 ( .A1(n4276), .A2(n4291), .A3(n4290), .ZN(n4228) );
  MUX2_X2 U5083 ( .A(n5183), .B(n2915), .S(n3312), .Z(net221874) );
  NOR2_X4 U5084 ( .A1(n4892), .A2(n4886), .ZN(n3558) );
  NAND2_X4 U5085 ( .A1(n3989), .A2(n7930), .ZN(n4102) );
  NAND3_X1 U5087 ( .A1(n7350), .A2(n7349), .A3(n7348), .ZN(regWrData[24]) );
  OAI22_X4 U5088 ( .A1(n7696), .A2(n3909), .B1(n7421), .B2(n3912), .ZN(n6070)
         );
  NOR2_X1 U5089 ( .A1(net224787), .A2(n2959), .ZN(n4824) );
  NAND2_X4 U5090 ( .A1(n5120), .A2(n5338), .ZN(n5340) );
  NOR2_X2 U5091 ( .A1(n5231), .A2(n3541), .ZN(n3560) );
  OAI211_X4 U5092 ( .C1(n7984), .C2(n5646), .A(n5810), .B(n3652), .ZN(n6044)
         );
  NOR2_X4 U5093 ( .A1(n7334), .A2(n7335), .ZN(n7337) );
  NAND2_X4 U5096 ( .A1(n3562), .A2(n3563), .ZN(n7326) );
  INV_X4 U5097 ( .A(n7066), .ZN(n3561) );
  INV_X2 U5098 ( .A(n5768), .ZN(n3564) );
  INV_X4 U5099 ( .A(n3857), .ZN(n3859) );
  INV_X4 U5100 ( .A(n7183), .ZN(n3565) );
  NAND2_X4 U5102 ( .A1(n4492), .A2(n3138), .ZN(n4495) );
  INV_X8 U5103 ( .A(n4490), .ZN(n4487) );
  OAI21_X4 U5104 ( .B1(net221411), .B2(n6420), .A(n6419), .ZN(n6421) );
  AOI21_X1 U5105 ( .B1(n7045), .B2(n2838), .A(n3165), .ZN(n7051) );
  AOI21_X1 U5106 ( .B1(net224843), .B2(n3165), .A(net224833), .ZN(n7049) );
  NAND2_X1 U5107 ( .A1(n7169), .A2(n5946), .ZN(n5957) );
  AOI21_X1 U5108 ( .B1(n6771), .B2(n2838), .A(n6770), .ZN(n6776) );
  INV_X4 U5109 ( .A(n6898), .ZN(n6904) );
  NOR2_X2 U5110 ( .A1(n6898), .A2(n3648), .ZN(n6916) );
  BUF_X32 U5111 ( .A(n2593), .Z(n3568) );
  INV_X8 U5112 ( .A(n5808), .ZN(n5813) );
  INV_X2 U5113 ( .A(n7931), .ZN(n4257) );
  INV_X8 U5114 ( .A(n5674), .ZN(n6449) );
  NAND2_X2 U5115 ( .A1(net228942), .A2(net220746), .ZN(n3741) );
  NAND3_X2 U5116 ( .A1(n4877), .A2(\wb/dsize_reg/z2 [30]), .A3(net225237), 
        .ZN(n4880) );
  INV_X4 U5117 ( .A(n3295), .ZN(net221153) );
  OAI21_X1 U5118 ( .B1(n4353), .B2(n3169), .A(n4212), .ZN(n4213) );
  NAND4_X2 U5119 ( .A1(n5891), .A2(n7987), .A3(n5555), .A4(n5893), .ZN(n5556)
         );
  INV_X2 U5120 ( .A(n5982), .ZN(n3892) );
  OAI21_X2 U5121 ( .B1(n2940), .B2(n5986), .A(n5985), .ZN(n7240) );
  NAND2_X4 U5122 ( .A1(n3897), .A2(n2991), .ZN(n4114) );
  XNOR2_X2 U5123 ( .A(n7179), .B(net224861), .ZN(n6777) );
  NAND2_X4 U5124 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  INV_X4 U5125 ( .A(n6908), .ZN(n3570) );
  INV_X4 U5126 ( .A(n6929), .ZN(n3571) );
  OAI211_X4 U5127 ( .C1(n7984), .C2(n5646), .A(n5810), .B(n3652), .ZN(n3573)
         );
  INV_X2 U5128 ( .A(n6755), .ZN(n3773) );
  INV_X2 U5130 ( .A(n3874), .ZN(n3877) );
  XNOR2_X2 U5131 ( .A(n5455), .B(n5454), .ZN(n5460) );
  NAND2_X2 U5132 ( .A1(n2901), .A2(net229061), .ZN(n3575) );
  NAND2_X4 U5133 ( .A1(n3574), .A2(n3575), .ZN(n5846) );
  INV_X4 U5134 ( .A(net229061), .ZN(net229719) );
  INV_X4 U5136 ( .A(n3576), .ZN(n3577) );
  NAND2_X1 U5137 ( .A1(n5846), .A2(net224861), .ZN(n3579) );
  NAND2_X2 U5139 ( .A1(n3579), .A2(n3580), .ZN(n5847) );
  INV_X2 U5140 ( .A(n5846), .ZN(n3578) );
  INV_X1 U5141 ( .A(net228159), .ZN(net228341) );
  NAND2_X2 U5142 ( .A1(n3980), .A2(n4148), .ZN(n3581) );
  INV_X4 U5143 ( .A(n3581), .ZN(n3582) );
  NAND2_X2 U5144 ( .A1(n7445), .A2(n3584), .ZN(n3586) );
  NAND2_X2 U5145 ( .A1(n3585), .A2(n3586), .ZN(n3979) );
  INV_X2 U5146 ( .A(n7260), .ZN(n7262) );
  INV_X4 U5147 ( .A(net224855), .ZN(net224853) );
  NAND3_X4 U5148 ( .A1(n3858), .A2(\wb/dsize_reg/z2 [21]), .A3(net225045), 
        .ZN(n5058) );
  INV_X1 U5149 ( .A(n7208), .ZN(n3587) );
  NAND2_X2 U5151 ( .A1(n7169), .A2(n6431), .ZN(n7199) );
  NOR2_X2 U5152 ( .A1(n4845), .A2(net224893), .ZN(\ex_mem/N112 ) );
  INV_X1 U5153 ( .A(n6594), .ZN(n3588) );
  INV_X1 U5154 ( .A(net221479), .ZN(net228150) );
  AOI21_X1 U5155 ( .B1(n3435), .B2(n4021), .A(n4020), .ZN(n3589) );
  NAND2_X4 U5156 ( .A1(n5467), .A2(net221442), .ZN(n5473) );
  OAI21_X1 U5157 ( .B1(n5465), .B2(n5466), .A(n5464), .ZN(n3824) );
  AOI21_X1 U5159 ( .B1(n2838), .B2(n6385), .A(n3309), .ZN(n6386) );
  INV_X8 U5160 ( .A(n5230), .ZN(n5707) );
  NOR3_X4 U5161 ( .A1(n5104), .A2(net220921), .A3(n5103), .ZN(n5105) );
  OAI21_X2 U5162 ( .B1(n5641), .B2(n3941), .A(n5636), .ZN(n6843) );
  XNOR2_X1 U5163 ( .A(n3178), .B(n4394), .ZN(n4395) );
  OAI21_X1 U5164 ( .B1(n6243), .B2(n3940), .A(n6242), .ZN(n6815) );
  NOR2_X2 U5165 ( .A1(n6820), .A2(n6819), .ZN(n6821) );
  INV_X2 U5166 ( .A(n6106), .ZN(regWrData[27]) );
  INV_X4 U5167 ( .A(n7128), .ZN(n7104) );
  NAND2_X2 U5168 ( .A1(n3453), .A2(n7002), .ZN(n7009) );
  NAND2_X1 U5169 ( .A1(n2898), .A2(net228909), .ZN(n3594) );
  NAND2_X4 U5170 ( .A1(n3593), .A2(n3594), .ZN(n6637) );
  INV_X4 U5171 ( .A(net228909), .ZN(net229646) );
  INV_X8 U5172 ( .A(n5260), .ZN(n6583) );
  NAND2_X2 U5173 ( .A1(n6772), .A2(n6432), .ZN(n7203) );
  BUF_X32 U5174 ( .A(n3750), .Z(n3595) );
  NAND3_X2 U5175 ( .A1(n4912), .A2(n4913), .A3(n4914), .ZN(n3750) );
  NOR2_X4 U5176 ( .A1(n5482), .A2(n5483), .ZN(n5484) );
  OAI21_X1 U5177 ( .B1(n3944), .B2(n5635), .A(n5634), .ZN(n5638) );
  NOR2_X4 U5178 ( .A1(n7089), .A2(net228150), .ZN(n7091) );
  INV_X4 U5179 ( .A(n3905), .ZN(n4829) );
  OAI22_X2 U5180 ( .A1(n5521), .A2(n5520), .B1(net224737), .B2(n5519), .ZN(
        n5537) );
  INV_X8 U5182 ( .A(n3596), .ZN(n3597) );
  NOR4_X4 U5183 ( .A1(n7301), .A2(n7299), .A3(n7300), .A4(n7298), .ZN(n7303)
         );
  NAND2_X1 U5185 ( .A1(n2932), .A2(net225434), .ZN(n3599) );
  INV_X1 U5186 ( .A(net225434), .ZN(net229606) );
  INV_X2 U5187 ( .A(n7241), .ZN(n7243) );
  OAI221_X4 U5188 ( .B1(n7694), .B2(n2578), .C1(n3942), .C2(n5705), .A(n5704), 
        .ZN(n6175) );
  NOR2_X1 U5190 ( .A1(n2652), .A2(n5624), .ZN(n4786) );
  NAND2_X1 U5191 ( .A1(n6105), .A2(n5624), .ZN(n5625) );
  NOR3_X2 U5192 ( .A1(n2606), .A2(n7546), .A3(n4865), .ZN(n4901) );
  INV_X8 U5193 ( .A(n5432), .ZN(n3812) );
  NAND2_X4 U5194 ( .A1(reg31Val_0[9]), .A2(net224783), .ZN(n5358) );
  NAND2_X2 U5196 ( .A1(n7169), .A2(n3768), .ZN(n6128) );
  NAND2_X2 U5197 ( .A1(n2859), .A2(net224743), .ZN(n3602) );
  INV_X1 U5199 ( .A(net224743), .ZN(net229596) );
  INV_X8 U5200 ( .A(n5927), .ZN(n7030) );
  AND2_X2 U5201 ( .A1(n3939), .A2(net225082), .ZN(n5317) );
  NOR2_X2 U5202 ( .A1(n7038), .A2(n7037), .ZN(n7043) );
  INV_X4 U5203 ( .A(n4453), .ZN(n4331) );
  INV_X1 U5204 ( .A(n3139), .ZN(n3603) );
  INV_X1 U5205 ( .A(n3542), .ZN(n6252) );
  NOR2_X2 U5206 ( .A1(n5324), .A2(n5323), .ZN(n5328) );
  NAND2_X4 U5207 ( .A1(net220875), .A2(n3484), .ZN(net221431) );
  NAND2_X4 U5208 ( .A1(n5191), .A2(n6381), .ZN(n6865) );
  INV_X1 U5209 ( .A(net224861), .ZN(net229579) );
  INV_X1 U5210 ( .A(net221759), .ZN(net229575) );
  NOR3_X4 U5211 ( .A1(n3374), .A2(n5814), .A3(n7135), .ZN(n7301) );
  NAND4_X4 U5212 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(
        regWrData[14]) );
  INV_X8 U5213 ( .A(regWrData[14]), .ZN(n5110) );
  NAND3_X2 U5214 ( .A1(n4877), .A2(\wb/dsize_reg/z2 [25]), .A3(n3898), .ZN(
        n4773) );
  NAND2_X2 U5215 ( .A1(n5565), .A2(n3401), .ZN(n3607) );
  NAND2_X4 U5216 ( .A1(n3600), .A2(n3286), .ZN(n3608) );
  NAND2_X4 U5217 ( .A1(n3607), .A2(n3608), .ZN(n7140) );
  XNOR2_X2 U5218 ( .A(net220921), .B(n6966), .ZN(net220305) );
  INV_X4 U5219 ( .A(n6966), .ZN(n6943) );
  INV_X1 U5220 ( .A(n3517), .ZN(n4756) );
  NOR2_X1 U5221 ( .A1(n7325), .A2(n3950), .ZN(n7120) );
  INV_X8 U5222 ( .A(n5803), .ZN(n5896) );
  NOR2_X2 U5223 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND3_X2 U5225 ( .A1(n5002), .A2(n5001), .A3(n5000), .ZN(n5543) );
  NAND3_X2 U5226 ( .A1(n6623), .A2(n6624), .A3(n6625), .ZN(n3612) );
  NOR2_X1 U5227 ( .A1(n3950), .A2(n7311), .ZN(n5781) );
  NAND3_X2 U5228 ( .A1(n3826), .A2(\wb/dsize_reg/z2 [27]), .A3(n5014), .ZN(
        n5218) );
  NAND2_X4 U5229 ( .A1(n6704), .A2(n6705), .ZN(n6676) );
  XNOR2_X2 U5230 ( .A(n6681), .B(n6680), .ZN(n6682) );
  NAND2_X1 U5231 ( .A1(net224737), .A2(n5605), .ZN(n5606) );
  INV_X1 U5232 ( .A(n5641), .ZN(regWrData[4]) );
  INV_X4 U5233 ( .A(n3305), .ZN(net220539) );
  NAND2_X4 U5234 ( .A1(n7080), .A2(net220632), .ZN(n3614) );
  NAND3_X1 U5235 ( .A1(n6216), .A2(n6215), .A3(n6214), .ZN(n6217) );
  AOI222_X4 U5236 ( .A1(n7127), .A2(n6728), .B1(n3953), .B2(n7122), .C1(n7126), 
        .C2(n3921), .ZN(n5881) );
  NAND2_X2 U5237 ( .A1(n5971), .A2(n7201), .ZN(n5761) );
  NOR2_X1 U5238 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  OAI21_X2 U5239 ( .B1(n5370), .B2(n5371), .A(n5369), .ZN(n5372) );
  NAND2_X4 U5241 ( .A1(n3617), .A2(n3618), .ZN(n6591) );
  INV_X8 U5242 ( .A(n5550), .ZN(n3616) );
  NAND2_X2 U5243 ( .A1(n2987), .A2(n3929), .ZN(n3620) );
  NAND2_X2 U5244 ( .A1(n3619), .A2(n3620), .ZN(n2176) );
  NAND2_X2 U5245 ( .A1(n6853), .A2(n3953), .ZN(n6854) );
  INV_X2 U5246 ( .A(net229481), .ZN(net229482) );
  NAND2_X2 U5248 ( .A1(n6168), .A2(n3868), .ZN(n3623) );
  NAND2_X4 U5249 ( .A1(n3621), .A2(n3622), .ZN(n3624) );
  NAND2_X1 U5251 ( .A1(n3924), .A2(n6803), .ZN(n6769) );
  INV_X8 U5253 ( .A(n4929), .ZN(n3902) );
  NAND2_X4 U5254 ( .A1(n7058), .A2(n6149), .ZN(n3646) );
  NAND2_X1 U5256 ( .A1(n7731), .A2(net225434), .ZN(n3627) );
  NAND2_X4 U5257 ( .A1(n3626), .A2(n3627), .ZN(n6167) );
  INV_X1 U5258 ( .A(net225434), .ZN(net229454) );
  MUX2_X2 U5259 ( .A(n6382), .B(n2905), .S(net228909), .Z(n5092) );
  AOI21_X1 U5260 ( .B1(n6014), .B2(n2838), .A(n3201), .ZN(n6020) );
  AOI21_X1 U5261 ( .B1(net224843), .B2(n3201), .A(net224835), .ZN(n6018) );
  OR2_X4 U5262 ( .A1(net224731), .A2(n2930), .ZN(n3628) );
  NAND2_X2 U5264 ( .A1(n6621), .A2(n7176), .ZN(n5958) );
  NOR2_X4 U5265 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  OAI21_X2 U5266 ( .B1(n3868), .B2(net230226), .A(n6880), .ZN(n6643) );
  NOR2_X4 U5267 ( .A1(n4314), .A2(n4313), .ZN(n4315) );
  NAND2_X4 U5269 ( .A1(n6209), .A2(n6210), .ZN(n5583) );
  NAND2_X4 U5270 ( .A1(n5966), .A2(n7201), .ZN(n5970) );
  NOR2_X4 U5271 ( .A1(n3386), .A2(n6906), .ZN(n3630) );
  NAND2_X2 U5273 ( .A1(net224865), .A2(n5620), .ZN(n5615) );
  NAND2_X1 U5274 ( .A1(net224865), .A2(n5636), .ZN(n5640) );
  NAND2_X4 U5275 ( .A1(n5099), .A2(net224995), .ZN(n5440) );
  NAND2_X1 U5276 ( .A1(n6485), .A2(net225029), .ZN(n6502) );
  NAND2_X1 U5277 ( .A1(net224913), .A2(n6485), .ZN(n6512) );
  OAI21_X1 U5278 ( .B1(n3945), .B2(n5653), .A(n3133), .ZN(n5654) );
  NOR2_X4 U5279 ( .A1(n3815), .A2(n2636), .ZN(n5951) );
  MUX2_X2 U5280 ( .A(reg31Val_3[1]), .B(reg31Val_0[1]), .S(net224723), .Z(
        n7750) );
  NAND3_X2 U5281 ( .A1(n4119), .A2(n4118), .A3(n4117), .ZN(n4126) );
  NAND3_X2 U5282 ( .A1(net224991), .A2(n5026), .A3(n7969), .ZN(n5029) );
  NOR3_X4 U5283 ( .A1(net220874), .A2(net220875), .A3(n6890), .ZN(n6891) );
  NAND3_X2 U5284 ( .A1(n6739), .A2(n5937), .A3(n6944), .ZN(n6441) );
  BUF_X32 U5285 ( .A(n6870), .Z(n3631) );
  NAND2_X4 U5286 ( .A1(n6390), .A2(net229393), .ZN(n3632) );
  NAND2_X4 U5287 ( .A1(n3632), .A2(n3633), .ZN(n6392) );
  INV_X4 U5288 ( .A(net228407), .ZN(net229393) );
  INV_X1 U5289 ( .A(net224733), .ZN(net228407) );
  NAND3_X4 U5290 ( .A1(n4737), .A2(n4738), .A3(n4739), .ZN(n6058) );
  NAND2_X4 U5291 ( .A1(n4885), .A2(n4884), .ZN(n4886) );
  INV_X4 U5292 ( .A(n3663), .ZN(n3664) );
  INV_X8 U5293 ( .A(n3634), .ZN(n7142) );
  INV_X4 U5294 ( .A(n5489), .ZN(n5487) );
  NAND2_X4 U5295 ( .A1(n3635), .A2(n5902), .ZN(n3637) );
  NAND2_X4 U5296 ( .A1(n3636), .A2(n3637), .ZN(n7283) );
  NAND3_X1 U5297 ( .A1(net228018), .A2(n2760), .A3(net228029), .ZN(n3638) );
  NAND2_X1 U5298 ( .A1(n2917), .A2(net225434), .ZN(n3641) );
  NAND2_X4 U5299 ( .A1(n3640), .A2(n3641), .ZN(n5050) );
  INV_X1 U5300 ( .A(net225434), .ZN(net229370) );
  AOI211_X4 U5301 ( .C1(n6160), .C2(n6159), .A(n3776), .B(n6158), .ZN(n3642)
         );
  INV_X4 U5302 ( .A(n5050), .ZN(n5777) );
  AOI211_X2 U5303 ( .C1(n6160), .C2(n6159), .A(n3776), .B(n6158), .ZN(n6645)
         );
  NAND4_X4 U5304 ( .A1(n6150), .A2(n3846), .A3(n6895), .A4(n6884), .ZN(n6158)
         );
  NAND2_X2 U5305 ( .A1(n6124), .A2(n3540), .ZN(n3699) );
  INV_X16 U5306 ( .A(n4504), .ZN(n4544) );
  INV_X16 U5307 ( .A(n3901), .ZN(n3643) );
  INV_X16 U5308 ( .A(n3901), .ZN(n4931) );
  BUF_X32 U5309 ( .A(n6233), .Z(n3644) );
  INV_X2 U5310 ( .A(n4846), .ZN(n4847) );
  NAND3_X2 U5311 ( .A1(n5996), .A2(n5997), .A3(n3947), .ZN(n5731) );
  NAND2_X4 U5312 ( .A1(n6124), .A2(n6943), .ZN(n5996) );
  INV_X2 U5313 ( .A(net220729), .ZN(net222151) );
  XNOR2_X2 U5314 ( .A(n6754), .B(n3666), .ZN(n7292) );
  NOR3_X4 U5315 ( .A1(n3892), .A2(n7174), .A3(n7173), .ZN(n7197) );
  NAND2_X1 U5316 ( .A1(n7239), .A2(n6495), .ZN(n5790) );
  OAI21_X2 U5317 ( .B1(n5626), .B2(n2595), .A(n5625), .ZN(n5627) );
  INV_X4 U5318 ( .A(net220746), .ZN(net228707) );
  NOR2_X2 U5319 ( .A1(n6896), .A2(n3452), .ZN(n3647) );
  INV_X8 U5320 ( .A(n4259), .ZN(n4261) );
  INV_X1 U5321 ( .A(n6790), .ZN(n3649) );
  NAND2_X1 U5322 ( .A1(n6822), .A2(n3588), .ZN(n6681) );
  NAND3_X2 U5323 ( .A1(net224861), .A2(n5382), .A3(net224737), .ZN(n5394) );
  NAND3_X2 U5324 ( .A1(n5469), .A2(net224861), .A3(n5474), .ZN(n5470) );
  NOR2_X2 U5325 ( .A1(net225230), .A2(n7571), .ZN(n3650) );
  INV_X4 U5326 ( .A(n3650), .ZN(n3651) );
  AOI21_X1 U5327 ( .B1(n4761), .B2(n4760), .A(net224903), .ZN(\ex_mem/N124 )
         );
  NOR2_X2 U5328 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  NAND2_X4 U5329 ( .A1(n4798), .A2(net228029), .ZN(n5006) );
  INV_X4 U5330 ( .A(n3652), .ZN(n3672) );
  INV_X16 U5331 ( .A(net223209), .ZN(net229307) );
  NAND2_X2 U5332 ( .A1(n6143), .A2(net227945), .ZN(net221763) );
  CLKBUF_X3 U5333 ( .A(n6883), .Z(n3701) );
  NAND2_X4 U5334 ( .A1(n4303), .A2(n4302), .ZN(n4221) );
  NAND3_X1 U5335 ( .A1(net220637), .A2(n2604), .A3(n7082), .ZN(n7095) );
  INV_X2 U5336 ( .A(n7080), .ZN(n7081) );
  NAND2_X1 U5337 ( .A1(n3924), .A2(n6728), .ZN(n6577) );
  NAND2_X1 U5338 ( .A1(n3953), .A2(n6728), .ZN(n6729) );
  NAND2_X2 U5339 ( .A1(n5676), .A2(n6462), .ZN(n6445) );
  NAND2_X2 U5340 ( .A1(n6540), .A2(n3924), .ZN(n5766) );
  NAND2_X2 U5341 ( .A1(n7048), .A2(n6064), .ZN(n3656) );
  INV_X2 U5342 ( .A(n7048), .ZN(n3655) );
  INV_X8 U5343 ( .A(n4312), .ZN(n4510) );
  INV_X4 U5344 ( .A(net229270), .ZN(net229271) );
  OAI21_X1 U5346 ( .B1(n4718), .B2(n3941), .A(net229952), .ZN(n6686) );
  AOI21_X1 U5347 ( .B1(n6394), .B2(n6096), .A(n6095), .ZN(n6137) );
  AOI21_X2 U5348 ( .B1(n5264), .B2(n3945), .A(n6101), .ZN(n5265) );
  INV_X1 U5349 ( .A(iAddr[2]), .ZN(n4560) );
  INV_X16 U5350 ( .A(n4465), .ZN(n3897) );
  INV_X1 U5351 ( .A(iAddr[23]), .ZN(n4507) );
  NAND2_X4 U5352 ( .A1(n4141), .A2(n4083), .ZN(n4156) );
  NAND2_X4 U5353 ( .A1(n4098), .A2(n4099), .ZN(n4141) );
  INV_X8 U5354 ( .A(net221818), .ZN(net221759) );
  INV_X2 U5355 ( .A(n5161), .ZN(n5162) );
  INV_X4 U5356 ( .A(n6892), .ZN(n6900) );
  NAND2_X4 U5357 ( .A1(n6253), .A2(n6254), .ZN(n5280) );
  NAND2_X4 U5358 ( .A1(n5709), .A2(memAddr[29]), .ZN(n6253) );
  NAND2_X4 U5360 ( .A1(n5119), .A2(n5338), .ZN(n5332) );
  NAND2_X1 U5362 ( .A1(n2764), .A2(net225434), .ZN(n3660) );
  NAND2_X4 U5363 ( .A1(n3659), .A2(n3660), .ZN(n6059) );
  INV_X1 U5364 ( .A(net225434), .ZN(net229239) );
  NAND3_X1 U5365 ( .A1(net225029), .A2(n3944), .A3(n5798), .ZN(n5433) );
  NAND3_X2 U5366 ( .A1(n6485), .A2(net225029), .A3(n5896), .ZN(n6699) );
  INV_X1 U5367 ( .A(n5903), .ZN(n3662) );
  OAI22_X2 U5368 ( .A1(n7534), .A2(n3912), .B1(n7690), .B2(n3909), .ZN(n5635)
         );
  OAI21_X1 U5369 ( .B1(n3944), .B2(n5514), .A(n3133), .ZN(n5515) );
  OAI21_X4 U5370 ( .B1(n2719), .B2(n3852), .A(n4988), .ZN(n5616) );
  INV_X4 U5371 ( .A(n5014), .ZN(n3852) );
  NAND2_X2 U5372 ( .A1(n4785), .A2(net225047), .ZN(n4988) );
  NAND2_X4 U5373 ( .A1(n6883), .A2(net228941), .ZN(n3665) );
  NAND2_X4 U5374 ( .A1(n2652), .A2(n6105), .ZN(n5621) );
  NAND4_X4 U5375 ( .A1(n5347), .A2(n5345), .A3(n5344), .A4(n5346), .ZN(n5348)
         );
  INV_X1 U5376 ( .A(n5633), .ZN(n3666) );
  NAND3_X4 U5377 ( .A1(n5130), .A2(n3668), .A3(n5206), .ZN(n5104) );
  NAND2_X4 U5378 ( .A1(n7232), .A2(n7224), .ZN(n7235) );
  INV_X2 U5379 ( .A(n6643), .ZN(n6640) );
  NAND2_X4 U5380 ( .A1(n3669), .A2(n3272), .ZN(n3671) );
  NAND2_X4 U5381 ( .A1(n3671), .A2(n3670), .ZN(n5574) );
  INV_X4 U5382 ( .A(n5570), .ZN(n3669) );
  NOR3_X2 U5383 ( .A1(net230741), .A2(n2730), .A3(n3710), .ZN(n6228) );
  NAND2_X4 U5384 ( .A1(n4359), .A2(iAddr[21]), .ZN(n3673) );
  NAND3_X4 U5385 ( .A1(n4500), .A2(n3674), .A3(iAddr[17]), .ZN(n4360) );
  INV_X8 U5386 ( .A(n3673), .ZN(n3674) );
  OAI21_X4 U5387 ( .B1(n4205), .B2(n4206), .A(n4204), .ZN(n3726) );
  NAND3_X2 U5388 ( .A1(n4485), .A2(n4484), .A3(n4483), .ZN(n4359) );
  NAND4_X4 U5389 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(
        iAddr[21]) );
  NAND2_X4 U5391 ( .A1(n6003), .A2(n7242), .ZN(n5679) );
  NAND2_X4 U5392 ( .A1(n5546), .A2(n6840), .ZN(n7288) );
  NOR2_X1 U5393 ( .A1(n6587), .A2(n6586), .ZN(n6590) );
  NAND3_X2 U5394 ( .A1(n5073), .A2(n5072), .A3(n5074), .ZN(n3679) );
  NAND2_X4 U5395 ( .A1(n3680), .A2(n5075), .ZN(n6812) );
  INV_X4 U5396 ( .A(n3679), .ZN(n3680) );
  INV_X16 U5398 ( .A(net230145), .ZN(net225017) );
  NAND2_X4 U5400 ( .A1(n4926), .A2(net225216), .ZN(n4927) );
  INV_X4 U5401 ( .A(n7039), .ZN(n7071) );
  OAI211_X2 U5403 ( .C1(n6965), .C2(n6964), .A(n7224), .B(n3823), .ZN(n6968)
         );
  INV_X2 U5404 ( .A(n6458), .ZN(n6460) );
  AOI21_X1 U5405 ( .B1(n3953), .B2(n7126), .A(n6513), .ZN(n6519) );
  AOI21_X1 U5406 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n7130) );
  OAI221_X4 U5407 ( .B1(n6619), .B2(n7205), .C1(n6618), .C2(n3914), .A(n6617), 
        .ZN(n6809) );
  NAND3_X2 U5408 ( .A1(n5038), .A2(n5490), .A3(n5037), .ZN(n5039) );
  INV_X8 U5409 ( .A(n3815), .ZN(n3816) );
  INV_X1 U5410 ( .A(n4346), .ZN(n3681) );
  INV_X1 U5411 ( .A(n4346), .ZN(n3682) );
  INV_X16 U5412 ( .A(net225001), .ZN(net224999) );
  INV_X8 U5413 ( .A(n5717), .ZN(n5869) );
  NAND3_X2 U5414 ( .A1(net224993), .A2(net224781), .A3(reg31Val_0[4]), .ZN(
        n4996) );
  NOR3_X4 U5415 ( .A1(n5529), .A2(n5528), .A3(net222515), .ZN(n5530) );
  NOR2_X4 U5417 ( .A1(n3684), .A2(net225051), .ZN(n3685) );
  NOR2_X4 U5418 ( .A1(n3685), .A2(n4918), .ZN(n4920) );
  INV_X4 U5419 ( .A(n4919), .ZN(n3684) );
  OAI22_X2 U5420 ( .A1(n7422), .A2(n7996), .B1(n7677), .B2(net225243), .ZN(
        n4918) );
  NAND3_X2 U5421 ( .A1(n4920), .A2(n4921), .A3(n4922), .ZN(n3843) );
  INV_X2 U5422 ( .A(n5498), .ZN(n4960) );
  INV_X1 U5423 ( .A(regWrData[11]), .ZN(n5715) );
  INV_X1 U5424 ( .A(n3294), .ZN(n5510) );
  NOR2_X1 U5425 ( .A1(net224733), .A2(n6396), .ZN(n6397) );
  NOR2_X4 U5426 ( .A1(n6078), .A2(n6077), .ZN(net221864) );
  NOR2_X4 U5427 ( .A1(n5769), .A2(n5770), .ZN(n5774) );
  NOR2_X4 U5428 ( .A1(net221754), .A2(net225588), .ZN(n6148) );
  INV_X8 U5429 ( .A(n6459), .ZN(n5692) );
  AND2_X2 U5430 ( .A1(n4302), .A2(n4291), .ZN(n3686) );
  AND2_X2 U5431 ( .A1(n4290), .A2(n3686), .ZN(n3740) );
  NAND2_X4 U5432 ( .A1(n4529), .A2(n3688), .ZN(n4531) );
  INV_X4 U5433 ( .A(n3687), .ZN(n3688) );
  NAND3_X2 U5434 ( .A1(n4350), .A2(n4349), .A3(n3094), .ZN(n4290) );
  INV_X8 U5435 ( .A(n4531), .ZN(n4543) );
  NOR4_X1 U5436 ( .A1(n4177), .A2(n4260), .A3(n4246), .A4(n4250), .ZN(n4008)
         );
  OAI211_X1 U5437 ( .C1(n5691), .C2(n3907), .A(n5055), .B(n5056), .ZN(n4873)
         );
  INV_X1 U5438 ( .A(n3638), .ZN(n4809) );
  NAND2_X4 U5439 ( .A1(net225017), .A2(n2977), .ZN(n7350) );
  NAND2_X4 U5440 ( .A1(net230143), .A2(net224783), .ZN(n6236) );
  MUX2_X2 U5441 ( .A(n4693), .B(n3047), .S(n3927), .Z(n2015) );
  INV_X4 U5442 ( .A(n5795), .ZN(n3690) );
  NAND2_X4 U5443 ( .A1(n6156), .A2(n6157), .ZN(n6159) );
  INV_X4 U5444 ( .A(n6733), .ZN(n5795) );
  NAND2_X4 U5445 ( .A1(n6357), .A2(net225029), .ZN(n5871) );
  INV_X8 U5446 ( .A(n5871), .ZN(n6040) );
  INV_X8 U5447 ( .A(n5057), .ZN(n5059) );
  NAND2_X4 U5448 ( .A1(n2679), .A2(n5055), .ZN(n5057) );
  NAND4_X2 U5449 ( .A1(n6476), .A2(n6475), .A3(n6474), .A4(n6473), .ZN(n7221)
         );
  MUX2_X2 U5450 ( .A(n3973), .B(reg31Val_0[31]), .S(net224691), .Z(n1915) );
  INV_X4 U5451 ( .A(net224691), .ZN(net224685) );
  NOR2_X2 U5452 ( .A1(n7639), .A2(net224901), .ZN(\ex_mem/N37 ) );
  OAI211_X4 U5453 ( .C1(n7197), .C2(n7267), .A(n7195), .B(n7196), .ZN(n7216)
         );
  NOR2_X1 U5454 ( .A1(net230231), .A2(n3950), .ZN(n7100) );
  NAND2_X4 U5455 ( .A1(n3691), .A2(n3692), .ZN(n3694) );
  NAND2_X4 U5456 ( .A1(n3693), .A2(n3694), .ZN(n6780) );
  INV_X4 U5457 ( .A(n6965), .ZN(n3692) );
  INV_X2 U5458 ( .A(n6669), .ZN(n6670) );
  NAND3_X2 U5459 ( .A1(n6172), .A2(n6171), .A3(n6170), .ZN(n6801) );
  XNOR2_X2 U5462 ( .A(n7439), .B(n3530), .ZN(n3695) );
  NAND3_X1 U5464 ( .A1(n3955), .A2(n6772), .A3(n6432), .ZN(n6433) );
  OAI22_X2 U5466 ( .A1(n2823), .A2(n3950), .B1(n7098), .B2(n2701), .ZN(n6615)
         );
  NOR2_X1 U5467 ( .A1(n3918), .A2(n2695), .ZN(n6614) );
  OAI21_X1 U5468 ( .B1(n2695), .B2(n3923), .A(n7036), .ZN(n7037) );
  OAI21_X2 U5469 ( .B1(n2695), .B2(n3954), .A(n7052), .ZN(n7069) );
  XNOR2_X1 U5471 ( .A(n3449), .B(n2973), .ZN(n5519) );
  AOI21_X1 U5472 ( .B1(n4810), .B2(n5097), .A(net224909), .ZN(\ex_mem/N105 )
         );
  OAI221_X4 U5473 ( .B1(n6412), .B2(n6639), .C1(net229330), .C2(n6412), .A(
        n6413), .ZN(n6414) );
  INV_X1 U5474 ( .A(n4453), .ZN(n4454) );
  NAND2_X1 U5475 ( .A1(iAddr[3]), .A2(iAddr[2]), .ZN(n4455) );
  INV_X1 U5476 ( .A(n4467), .ZN(n4468) );
  NAND3_X4 U5477 ( .A1(n4866), .A2(net224783), .A3(net225251), .ZN(net223338)
         );
  NAND2_X4 U5478 ( .A1(n5709), .A2(memAddr[1]), .ZN(n6209) );
  INV_X4 U5479 ( .A(n7496), .ZN(n4868) );
  NAND2_X4 U5480 ( .A1(n5671), .A2(n5670), .ZN(n6257) );
  XNOR2_X2 U5481 ( .A(n5050), .B(n3272), .ZN(n5778) );
  MUX2_X2 U5482 ( .A(reg31Val_3[0]), .B(reg31Val_0[0]), .S(net224717), .Z(
        n7751) );
  NAND3_X1 U5483 ( .A1(n4524), .A2(n4463), .A3(n3091), .ZN(n4464) );
  XNOR2_X1 U5484 ( .A(n4458), .B(n4463), .ZN(n4459) );
  NAND2_X4 U5485 ( .A1(reg31Val_3[0]), .A2(n4462), .ZN(n4463) );
  NAND3_X4 U5486 ( .A1(n3867), .A2(n3849), .A3(net223209), .ZN(n4715) );
  INV_X8 U5487 ( .A(n4802), .ZN(n3849) );
  INV_X4 U5488 ( .A(n4715), .ZN(n3813) );
  INV_X1 U5489 ( .A(n5304), .ZN(n5129) );
  NOR3_X2 U5490 ( .A1(n6183), .A2(n6182), .A3(n6181), .ZN(n6204) );
  NAND2_X4 U5491 ( .A1(n3702), .A2(net228982), .ZN(n6370) );
  INV_X1 U5492 ( .A(net224737), .ZN(net228981) );
  NOR2_X1 U5494 ( .A1(n2729), .A2(n4772), .ZN(n4714) );
  NAND2_X4 U5495 ( .A1(n6456), .A2(n6455), .ZN(n7222) );
  NAND3_X4 U5496 ( .A1(net228287), .A2(\wb/dsize_reg/z2 [22]), .A3(n3906), 
        .ZN(n3703) );
  INV_X16 U5497 ( .A(n4887), .ZN(n3906) );
  NAND2_X2 U5498 ( .A1(n3303), .A2(n7331), .ZN(n7334) );
  NAND3_X2 U5499 ( .A1(net229330), .A2(n6989), .A3(net228942), .ZN(n6647) );
  NAND2_X2 U5500 ( .A1(n3643), .A2(memAddr[12]), .ZN(n5021) );
  NAND4_X4 U5501 ( .A1(n7349), .A2(n5660), .A3(n7348), .A4(n7350), .ZN(n6045)
         );
  INV_X4 U5502 ( .A(n3453), .ZN(n3719) );
  INV_X4 U5503 ( .A(n5223), .ZN(n7352) );
  OAI22_X2 U5504 ( .A1(n7572), .A2(net225015), .B1(n2733), .B2(n3933), .ZN(
        n5223) );
  OAI21_X4 U5505 ( .B1(n7240), .B2(n3310), .A(n7194), .ZN(n7195) );
  NAND2_X4 U5506 ( .A1(n7931), .A2(n4347), .ZN(n4178) );
  NAND2_X4 U5507 ( .A1(n5094), .A2(n5441), .ZN(n5173) );
  NAND2_X4 U5508 ( .A1(n6069), .A2(n7108), .ZN(net220728) );
  NAND2_X1 U5509 ( .A1(n4534), .A2(n8108), .ZN(n4536) );
  NAND2_X4 U5510 ( .A1(n5059), .A2(n5058), .ZN(n5534) );
  OAI21_X2 U5511 ( .B1(n6076), .B2(n2595), .A(n6074), .ZN(n6077) );
  NAND2_X1 U5512 ( .A1(n7727), .A2(net225434), .ZN(n3705) );
  NAND2_X4 U5513 ( .A1(n3704), .A2(n3705), .ZN(n5486) );
  INV_X1 U5514 ( .A(net225434), .ZN(net228936) );
  NAND3_X4 U5515 ( .A1(n5727), .A2(n5734), .A3(n5726), .ZN(n6495) );
  INV_X4 U5516 ( .A(n6911), .ZN(n7096) );
  NAND3_X4 U5517 ( .A1(n4198), .A2(n4323), .A3(n4197), .ZN(n4199) );
  NAND2_X2 U5518 ( .A1(reg31Val_0[10]), .A2(n3898), .ZN(n5386) );
  NAND2_X4 U5519 ( .A1(n3706), .A2(n3947), .ZN(n6459) );
  NAND2_X4 U5520 ( .A1(n6340), .A2(net225029), .ZN(n6080) );
  NAND2_X4 U5521 ( .A1(n3964), .A2(n4391), .ZN(n3965) );
  NOR4_X4 U5522 ( .A1(n3445), .A2(net225051), .A3(n3290), .A4(n7560), .ZN(
        n5025) );
  NAND2_X4 U5523 ( .A1(net228915), .A2(n3707), .ZN(n3708) );
  INV_X2 U5524 ( .A(net223242), .ZN(net228915) );
  INV_X4 U5525 ( .A(n4928), .ZN(n3707) );
  NAND2_X4 U5526 ( .A1(net228018), .A2(net228597), .ZN(n4865) );
  INV_X8 U5527 ( .A(n7142), .ZN(n7144) );
  OAI211_X4 U5528 ( .C1(n3712), .C2(n5253), .A(n5252), .B(n3947), .ZN(n5984)
         );
  NAND2_X4 U5529 ( .A1(n7009), .A2(n7003), .ZN(n7010) );
  NOR2_X2 U5530 ( .A1(net220354), .A2(n3249), .ZN(n7319) );
  NAND2_X4 U5531 ( .A1(iAddr[24]), .A2(iAddr[23]), .ZN(n4312) );
  BUF_X32 U5532 ( .A(n6875), .Z(n3709) );
  NAND2_X4 U5533 ( .A1(n3882), .A2(n3784), .ZN(n5136) );
  INV_X4 U5534 ( .A(n6445), .ZN(n5677) );
  OAI21_X4 U5535 ( .B1(n6939), .B2(n7225), .A(n7228), .ZN(n6940) );
  AOI211_X1 U5536 ( .C1(n7919), .C2(regWrData[7]), .A(n4720), .B(n3130), .ZN(
        n4721) );
  INV_X4 U5537 ( .A(n5950), .ZN(n5758) );
  OAI221_X4 U5538 ( .B1(n7671), .B2(net224901), .C1(n4040), .C2(n4039), .A(
        n4038), .ZN(iAddr[16]) );
  OAI21_X2 U5539 ( .B1(n4037), .B2(n4173), .A(n4524), .ZN(n4039) );
  INV_X4 U5540 ( .A(net221765), .ZN(net227945) );
  NAND3_X2 U5541 ( .A1(n4784), .A2(n2598), .A3(n3283), .ZN(n3710) );
  OAI22_X4 U5542 ( .A1(n7525), .A2(n3912), .B1(n7687), .B2(n3909), .ZN(n6233)
         );
  INV_X2 U5543 ( .A(n5334), .ZN(n5333) );
  NOR3_X2 U5544 ( .A1(n3905), .A2(n3899), .A3(n7549), .ZN(n4909) );
  NAND2_X4 U5545 ( .A1(n7085), .A2(n2645), .ZN(n7088) );
  NAND2_X4 U5546 ( .A1(n4249), .A2(n3975), .ZN(n4177) );
  BUF_X32 U5547 ( .A(n6548), .Z(n3711) );
  INV_X4 U5548 ( .A(net220640), .ZN(net228869) );
  OAI21_X1 U5549 ( .B1(n4439), .B2(n4472), .A(n4438), .ZN(n4440) );
  XNOR2_X1 U5550 ( .A(iAddr[11]), .B(n7929), .ZN(n4710) );
  OAI211_X4 U5551 ( .C1(n5947), .C2(n5939), .A(n5703), .B(n5734), .ZN(n5860)
         );
  OAI221_X4 U5552 ( .B1(n6619), .B2(n6672), .C1(n6618), .C2(n2703), .A(n5995), 
        .ZN(n6853) );
  AOI21_X2 U5553 ( .B1(n6191), .B2(n7201), .A(n5954), .ZN(n5875) );
  OAI211_X4 U5554 ( .C1(n5950), .C2(n5871), .A(n5870), .B(n3948), .ZN(n6191)
         );
  BUF_X32 U5555 ( .A(net229624), .Z(net228858) );
  AOI22_X1 U5556 ( .A1(n5357), .A2(net224993), .B1(\wb/dsize_reg/z2 [9]), .B2(
        n3934), .ZN(n6239) );
  AOI21_X2 U5557 ( .B1(n5273), .B2(net224993), .A(n5272), .ZN(n6246) );
  NAND3_X2 U5558 ( .A1(net224993), .A2(n3079), .A3(n4829), .ZN(n5526) );
  INV_X8 U5559 ( .A(n5869), .ZN(n3712) );
  BUF_X32 U5560 ( .A(n6138), .Z(n3713) );
  NAND3_X2 U5561 ( .A1(n6655), .A2(n6656), .A3(n3124), .ZN(\ex_mem/N225 ) );
  NAND2_X1 U5562 ( .A1(n3924), .A2(n6801), .ZN(n6657) );
  NOR2_X2 U5563 ( .A1(n6654), .A2(n6653), .ZN(n6656) );
  AOI22_X2 U5564 ( .A1(n3921), .A2(n3166), .B1(n6803), .B2(n7127), .ZN(n6655)
         );
  AOI21_X4 U5565 ( .B1(n7167), .B2(net220535), .A(net220536), .ZN(n7273) );
  INV_X8 U5566 ( .A(n7310), .ZN(n7312) );
  NAND2_X4 U5567 ( .A1(net228094), .A2(net220312), .ZN(n7336) );
  INV_X2 U5568 ( .A(n6610), .ZN(n5834) );
  NOR2_X2 U5569 ( .A1(n3914), .A2(n6610), .ZN(n6611) );
  NAND3_X2 U5570 ( .A1(n4824), .A2(net225237), .A3(net225216), .ZN(n4825) );
  INV_X8 U5571 ( .A(n5583), .ZN(n5589) );
  NAND2_X1 U5572 ( .A1(n7020), .A2(net220714), .ZN(n3717) );
  NAND2_X1 U5573 ( .A1(n3718), .A2(n7112), .ZN(n7022) );
  INV_X4 U5574 ( .A(n3717), .ZN(n3718) );
  OAI21_X1 U5575 ( .B1(n6976), .B2(net220775), .A(n6975), .ZN(n6977) );
  INV_X2 U5576 ( .A(net220775), .ZN(net220780) );
  OAI22_X2 U5577 ( .A1(n7532), .A2(n3912), .B1(n7693), .B2(n3909), .ZN(n5571)
         );
  NAND2_X4 U5578 ( .A1(net228816), .A2(n3719), .ZN(n3720) );
  NAND2_X4 U5579 ( .A1(n6885), .A2(n3720), .ZN(n6920) );
  INV_X4 U5580 ( .A(net225588), .ZN(net220882) );
  NAND2_X2 U5581 ( .A1(net220409), .A2(net228541), .ZN(n3721) );
  NAND2_X4 U5583 ( .A1(net221812), .A2(n6115), .ZN(n6117) );
  NAND2_X2 U5584 ( .A1(net221792), .A2(net230733), .ZN(n7275) );
  OAI22_X2 U5585 ( .A1(n7537), .A2(n3912), .B1(n7697), .B2(n3909), .ZN(n5661)
         );
  NOR2_X4 U5586 ( .A1(net221479), .A2(net220640), .ZN(net228809) );
  INV_X8 U5587 ( .A(n7113), .ZN(n6042) );
  NAND2_X4 U5588 ( .A1(n4208), .A2(n4346), .ZN(n4018) );
  AOI22_X4 U5589 ( .A1(net223245), .A2(n2707), .B1(n4931), .B2(memAddr[30]), 
        .ZN(n4857) );
  INV_X8 U5590 ( .A(n6796), .ZN(n6790) );
  BUF_X8 U5591 ( .A(net225102), .Z(net228697) );
  INV_X1 U5592 ( .A(n7143), .ZN(n7145) );
  INV_X1 U5593 ( .A(n5154), .ZN(n7155) );
  AOI21_X2 U5594 ( .B1(n6852), .B2(n3953), .A(n6767), .ZN(n6768) );
  NAND2_X2 U5595 ( .A1(n4956), .A2(net225047), .ZN(n4957) );
  OAI21_X4 U5596 ( .B1(net230741), .B2(n4958), .A(n4957), .ZN(n5499) );
  INV_X8 U5598 ( .A(n6915), .ZN(n6883) );
  INV_X8 U5599 ( .A(n3751), .ZN(n3948) );
  NAND3_X4 U5600 ( .A1(n5763), .A2(n5764), .A3(n5765), .ZN(n6545) );
  NAND2_X2 U5601 ( .A1(n3955), .A2(n6659), .ZN(n5764) );
  AOI22_X4 U5602 ( .A1(n7176), .A2(n5876), .B1(n7239), .B2(n5762), .ZN(n5763)
         );
  NAND2_X2 U5603 ( .A1(n6877), .A2(n6892), .ZN(n6878) );
  INV_X8 U5604 ( .A(n7171), .ZN(n3949) );
  NAND3_X2 U5605 ( .A1(n6044), .A2(n6043), .A3(n5647), .ZN(n3727) );
  NAND3_X2 U5606 ( .A1(n3573), .A2(n6043), .A3(n5647), .ZN(n6151) );
  INV_X4 U5607 ( .A(n7317), .ZN(n7320) );
  NAND2_X4 U5610 ( .A1(n3730), .A2(n3731), .ZN(n6753) );
  INV_X1 U5613 ( .A(net224787), .ZN(net228276) );
  NOR2_X2 U5614 ( .A1(n7668), .A2(net224895), .ZN(\ex_mem/N46 ) );
  INV_X16 U5615 ( .A(n3949), .ZN(n3856) );
  NAND2_X4 U5616 ( .A1(n6462), .A2(n6772), .ZN(n3874) );
  NAND2_X2 U5617 ( .A1(n6912), .A2(n6926), .ZN(n3841) );
  NOR2_X4 U5618 ( .A1(n3703), .A2(net228735), .ZN(n3733) );
  NOR2_X4 U5619 ( .A1(n3733), .A2(n4736), .ZN(n4737) );
  INV_X1 U5620 ( .A(net224993), .ZN(net228735) );
  NOR2_X4 U5621 ( .A1(net225102), .A2(n3867), .ZN(n3734) );
  NOR2_X4 U5622 ( .A1(n5770), .A2(n3564), .ZN(n5019) );
  INV_X4 U5623 ( .A(n3747), .ZN(n6201) );
  OAI21_X1 U5624 ( .B1(n7292), .B2(n3950), .A(n6763), .ZN(n6764) );
  OAI22_X2 U5625 ( .A1(n6778), .A2(n7179), .B1(net224865), .B2(n7177), .ZN(
        n6779) );
  AOI21_X4 U5626 ( .B1(n5610), .B2(n6777), .A(n5609), .ZN(n5612) );
  NAND3_X2 U5627 ( .A1(n6202), .A2(n6203), .A3(n6204), .ZN(\ex_mem/N224 ) );
  NAND2_X2 U5628 ( .A1(n6852), .A2(n7127), .ZN(n6203) );
  NAND3_X4 U5629 ( .A1(n5033), .A2(n3736), .A3(n5035), .ZN(n5493) );
  INV_X4 U5630 ( .A(n3735), .ZN(n3736) );
  NAND2_X2 U5631 ( .A1(net225588), .A2(n7097), .ZN(n3738) );
  NAND2_X4 U5632 ( .A1(n3737), .A2(net228720), .ZN(n3739) );
  INV_X4 U5633 ( .A(n5493), .ZN(n5038) );
  NAND2_X2 U5634 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  INV_X4 U5635 ( .A(n2583), .ZN(n6931) );
  NAND2_X4 U5636 ( .A1(n3741), .A2(net228710), .ZN(n7331) );
  INV_X1 U5637 ( .A(n6714), .ZN(n6553) );
  NAND2_X4 U5638 ( .A1(n6335), .A2(net225029), .ZN(n5821) );
  NAND2_X1 U5639 ( .A1(n6661), .A2(n7212), .ZN(n6439) );
  AOI22_X2 U5640 ( .A1(n3955), .A2(n7212), .B1(n2681), .B2(n6661), .ZN(n6200)
         );
  INV_X16 U5641 ( .A(net224753), .ZN(net224749) );
  INV_X4 U5642 ( .A(n7088), .ZN(n7089) );
  NOR3_X2 U5643 ( .A1(n4777), .A2(net222840), .A3(n2784), .ZN(n4919) );
  INV_X4 U5644 ( .A(n3765), .ZN(n3742) );
  OAI211_X4 U5645 ( .C1(n4226), .C2(n4227), .A(n4225), .B(n4224), .ZN(
        iAddr[26]) );
  AOI22_X2 U5647 ( .A1(memAddr[12]), .A2(n8014), .B1(n3744), .B2(n5710), .ZN(
        n3743) );
  NAND3_X2 U5648 ( .A1(net221793), .A2(n6119), .A3(net220601), .ZN(net228080)
         );
  NAND2_X4 U5649 ( .A1(net221800), .A2(net221793), .ZN(net221798) );
  NAND2_X4 U5650 ( .A1(n6090), .A2(net224995), .ZN(n6091) );
  NAND2_X4 U5651 ( .A1(n6092), .A2(n6091), .ZN(n6104) );
  INV_X2 U5652 ( .A(n6843), .ZN(n6205) );
  AOI21_X1 U5653 ( .B1(n3951), .B2(n7300), .A(n6743), .ZN(n6744) );
  NOR2_X1 U5654 ( .A1(n6359), .A2(n6843), .ZN(n6360) );
  NAND2_X1 U5655 ( .A1(n7358), .A2(n6843), .ZN(n6844) );
  NAND2_X4 U5656 ( .A1(n6843), .A2(net225029), .ZN(n6845) );
  INV_X2 U5657 ( .A(n4992), .ZN(n4995) );
  INV_X4 U5658 ( .A(net220540), .ZN(net220312) );
  NAND2_X4 U5659 ( .A1(n4055), .A2(n4054), .ZN(n4061) );
  NAND2_X1 U5660 ( .A1(n3902), .A2(\wb/dsize_reg/z2 [18]), .ZN(n4896) );
  NAND2_X1 U5661 ( .A1(reg31Val_0[14]), .A2(n3902), .ZN(n4876) );
  NAND2_X1 U5662 ( .A1(n3902), .A2(n2799), .ZN(n4875) );
  OAI22_X4 U5664 ( .A1(n7205), .A2(n6668), .B1(n6667), .B2(n3914), .ZN(n6675)
         );
  AOI22_X4 U5665 ( .A1(n3955), .A2(n6622), .B1(n6621), .B2(n6661), .ZN(n6623)
         );
  XNOR2_X1 U5666 ( .A(n4387), .B(n2768), .ZN(n4388) );
  XNOR2_X1 U5667 ( .A(n4383), .B(n4382), .ZN(n4384) );
  XOR2_X1 U5668 ( .A(n4404), .B(n7509), .Z(n4405) );
  NOR3_X1 U5669 ( .A1(n6861), .A2(n7190), .A3(net224899), .ZN(n6339) );
  OAI21_X1 U5670 ( .B1(net220310), .B2(n6966), .A(n7193), .ZN(n6967) );
  NAND2_X4 U5671 ( .A1(n6861), .A2(net225029), .ZN(n6966) );
  NAND2_X2 U5672 ( .A1(n6838), .A2(n2592), .ZN(n6710) );
  NAND3_X2 U5673 ( .A1(n3859), .A2(\wb/dsize_reg/z2 [17]), .A3(net224991), 
        .ZN(n5588) );
  NAND2_X4 U5674 ( .A1(n5084), .A2(n3907), .ZN(n3746) );
  NAND2_X4 U5675 ( .A1(n5994), .A2(n5993), .ZN(n3747) );
  INV_X8 U5676 ( .A(n5083), .ZN(n5084) );
  NAND2_X2 U5677 ( .A1(net221153), .A2(net220714), .ZN(n3748) );
  NAND2_X2 U5678 ( .A1(n3749), .A2(n6117), .ZN(n6118) );
  INV_X4 U5679 ( .A(n3748), .ZN(n3749) );
  NAND2_X4 U5681 ( .A1(net220292), .A2(net220293), .ZN(net220409) );
  OAI22_X4 U5682 ( .A1(n5354), .A2(n5353), .B1(n5352), .B2(n5353), .ZN(n5452)
         );
  AOI21_X1 U5683 ( .B1(n7028), .B2(n2838), .A(n7029), .ZN(n7035) );
  AOI21_X1 U5684 ( .B1(net224843), .B2(n7029), .A(net224835), .ZN(n7033) );
  INV_X1 U5685 ( .A(n6751), .ZN(n3754) );
  NAND2_X1 U5686 ( .A1(n4445), .A2(n4467), .ZN(n4446) );
  NOR2_X1 U5687 ( .A1(n4447), .A2(n4453), .ZN(n4449) );
  XNOR2_X1 U5688 ( .A(n4467), .B(iAddr[9]), .ZN(n4555) );
  XNOR2_X1 U5689 ( .A(n4453), .B(iAddr[5]), .ZN(n4553) );
  NAND2_X4 U5690 ( .A1(n4812), .A2(n4719), .ZN(n5082) );
  NAND2_X1 U5691 ( .A1(n3951), .A2(n7335), .ZN(n6483) );
  OAI22_X2 U5692 ( .A1(n7415), .A2(n3901), .B1(n7682), .B2(net225243), .ZN(
        n4902) );
  NOR2_X2 U5693 ( .A1(n7681), .A2(net225243), .ZN(n4729) );
  OAI221_X4 U5695 ( .B1(n4233), .B2(n4184), .C1(n4185), .C2(n4177), .A(n4187), 
        .ZN(n4022) );
  INV_X8 U5696 ( .A(net225096), .ZN(net223346) );
  NAND3_X2 U5697 ( .A1(net220849), .A2(n3205), .A3(net220851), .ZN(n6927) );
  NAND2_X2 U5698 ( .A1(net224859), .A2(n5631), .ZN(n3756) );
  NAND2_X4 U5699 ( .A1(n3755), .A2(net228610), .ZN(n3757) );
  INV_X1 U5701 ( .A(net224859), .ZN(net228610) );
  NAND2_X4 U5702 ( .A1(n5175), .A2(n5174), .ZN(n5371) );
  NAND2_X1 U5704 ( .A1(n5780), .A2(n6373), .ZN(n3760) );
  NAND2_X4 U5705 ( .A1(n3758), .A2(n3759), .ZN(n3761) );
  NAND2_X4 U5706 ( .A1(n3760), .A2(n3761), .ZN(n7311) );
  INV_X4 U5707 ( .A(n5780), .ZN(n3758) );
  INV_X1 U5708 ( .A(n6373), .ZN(n3759) );
  XNOR2_X1 U5709 ( .A(n5551), .B(n5550), .ZN(n3762) );
  NAND2_X2 U5710 ( .A1(n6458), .A2(n5692), .ZN(n3763) );
  OAI22_X4 U5711 ( .A1(n6667), .A2(n6672), .B1(n2703), .B2(n6671), .ZN(n6603)
         );
  NAND2_X4 U5712 ( .A1(n3766), .A2(n3767), .ZN(net228541) );
  NAND2_X4 U5713 ( .A1(n6343), .A2(net225029), .ZN(n5776) );
  NAND2_X4 U5714 ( .A1(n5449), .A2(n6739), .ZN(n6823) );
  NAND2_X2 U5715 ( .A1(n6739), .A2(n6462), .ZN(n5239) );
  XNOR2_X2 U5716 ( .A(n6372), .B(net228150), .ZN(n7285) );
  XNOR2_X2 U5717 ( .A(n6838), .B(n3828), .ZN(n6839) );
  NOR2_X4 U5718 ( .A1(net221924), .A2(n3614), .ZN(n3846) );
  OAI211_X1 U5719 ( .C1(n3907), .C2(n5268), .A(n5022), .B(n5021), .ZN(n4839)
         );
  NAND2_X4 U5721 ( .A1(n5084), .A2(n5309), .ZN(n5323) );
  NAND2_X4 U5722 ( .A1(n5125), .A2(n5124), .ZN(n5324) );
  NAND3_X2 U5723 ( .A1(n4714), .A2(n4713), .A3(net225251), .ZN(n5310) );
  INV_X1 U5724 ( .A(n2694), .ZN(n3764) );
  OAI21_X1 U5725 ( .B1(n6818), .B2(n3557), .A(n6816), .ZN(n6819) );
  NOR2_X1 U5726 ( .A1(n7242), .A2(n3557), .ZN(n5962) );
  NAND2_X2 U5727 ( .A1(net220757), .A2(n3652), .ZN(n6983) );
  NAND2_X4 U5728 ( .A1(n3695), .A2(n4120), .ZN(n4128) );
  NOR2_X2 U5729 ( .A1(n7638), .A2(net224901), .ZN(\ex_mem/N38 ) );
  INV_X4 U5730 ( .A(n7274), .ZN(n3766) );
  INV_X4 U5731 ( .A(n7273), .ZN(n3767) );
  NOR2_X4 U5732 ( .A1(n3249), .A2(n7165), .ZN(n7274) );
  OAI222_X2 U5733 ( .A1(n7574), .A2(net225015), .B1(n2729), .B2(n3933), .C1(
        n3935), .C2(n3080), .ZN(regWrData[23]) );
  MUX2_X2 U5734 ( .A(n5080), .B(n7732), .S(net227817), .Z(n3770) );
  INV_X1 U5736 ( .A(n6741), .ZN(n6735) );
  NAND2_X2 U5737 ( .A1(n5007), .A2(n5011), .ZN(n3844) );
  NAND2_X1 U5738 ( .A1(reg31Val_0[3]), .A2(net224783), .ZN(n5011) );
  INV_X8 U5739 ( .A(n5012), .ZN(n5007) );
  INV_X8 U5740 ( .A(n6461), .ZN(n6944) );
  NOR2_X1 U5741 ( .A1(n7939), .A2(net220775), .ZN(n5935) );
  NOR2_X1 U5742 ( .A1(n7939), .A2(n6125), .ZN(n6126) );
  NOR2_X1 U5743 ( .A1(n7939), .A2(n3309), .ZN(n6424) );
  NAND2_X4 U5744 ( .A1(n3960), .A2(n4382), .ZN(n3961) );
  INV_X8 U5745 ( .A(n3968), .ZN(n4409) );
  NOR3_X4 U5746 ( .A1(n4772), .A2(net228697), .A3(net224783), .ZN(n4877) );
  NOR2_X4 U5747 ( .A1(n4775), .A2(n4774), .ZN(n5075) );
  INV_X1 U5748 ( .A(n3595), .ZN(n4915) );
  NAND2_X2 U5749 ( .A1(n4751), .A2(net228287), .ZN(n4753) );
  NOR2_X2 U5750 ( .A1(n2730), .A2(n3899), .ZN(n4751) );
  INV_X1 U5752 ( .A(n7861), .ZN(n4491) );
  MUX2_X2 U5753 ( .A(n5301), .B(n2896), .S(net230088), .Z(n7183) );
  INV_X8 U5754 ( .A(n5341), .ZN(n5347) );
  OAI211_X1 U5755 ( .C1(n5284), .C2(n3907), .A(n4986), .B(n4987), .ZN(n4787)
         );
  NAND2_X2 U5756 ( .A1(n7086), .A2(net228869), .ZN(n7087) );
  NAND3_X2 U5757 ( .A1(\wb/dsize_reg/z2 [19]), .A2(net228018), .A3(net228597), 
        .ZN(net223345) );
  OAI21_X1 U5758 ( .B1(n4537), .B2(n4532), .A(n4533), .ZN(n4516) );
  INV_X4 U5759 ( .A(net224871), .ZN(net224869) );
  INV_X8 U5760 ( .A(net224861), .ZN(net227884) );
  INV_X2 U5761 ( .A(net224861), .ZN(net228323) );
  INV_X8 U5762 ( .A(net220720), .ZN(net220714) );
  NOR2_X4 U5763 ( .A1(n3772), .A2(n3864), .ZN(n3771) );
  NAND2_X4 U5764 ( .A1(n5574), .A2(n5573), .ZN(n6750) );
  INV_X8 U5765 ( .A(n5359), .ZN(n4856) );
  NAND2_X4 U5767 ( .A1(n5415), .A2(n5414), .ZN(n5409) );
  NAND2_X2 U5768 ( .A1(n5961), .A2(n3816), .ZN(n6427) );
  NAND2_X2 U5769 ( .A1(n4993), .A2(n4996), .ZN(n3777) );
  NAND3_X4 U5770 ( .A1(n5002), .A2(n4992), .A3(n3778), .ZN(n7908) );
  INV_X4 U5771 ( .A(n3777), .ZN(n3778) );
  OR2_X2 U5772 ( .A1(n5641), .A2(n2595), .ZN(n3779) );
  OR2_X2 U5773 ( .A1(n7908), .A2(n5640), .ZN(n3780) );
  NAND3_X4 U5774 ( .A1(n3779), .A2(n3780), .A3(n5639), .ZN(n5643) );
  NAND3_X2 U5775 ( .A1(net224991), .A2(n3122), .A3(n3904), .ZN(n4993) );
  NAND2_X4 U5776 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND3_X2 U5777 ( .A1(n3885), .A2(n5707), .A3(n6406), .ZN(n5855) );
  NAND3_X2 U5778 ( .A1(n3885), .A2(n3373), .A3(n7150), .ZN(n6950) );
  NAND3_X2 U5779 ( .A1(n3373), .A2(n3885), .A3(net221494), .ZN(n6184) );
  NAND3_X4 U5780 ( .A1(n5945), .A2(n7935), .A3(n5944), .ZN(n6621) );
  INV_X8 U5782 ( .A(n5541), .ZN(n5463) );
  INV_X1 U5783 ( .A(n3207), .ZN(n3781) );
  NAND3_X4 U5784 ( .A1(n4272), .A2(n4273), .A3(n4271), .ZN(iAddr[30]) );
  NOR2_X2 U5785 ( .A1(net220640), .A2(n7081), .ZN(n7082) );
  OAI21_X2 U5786 ( .B1(net220640), .B2(net221477), .A(n6374), .ZN(n6375) );
  NAND2_X4 U5787 ( .A1(n4973), .A2(n3907), .ZN(n4977) );
  NAND4_X2 U5788 ( .A1(n5586), .A2(n5584), .A3(net224737), .A4(n5587), .ZN(
        n5596) );
  NOR3_X2 U5789 ( .A1(n5417), .A2(n3920), .A3(n3936), .ZN(n5420) );
  INV_X16 U5790 ( .A(n3920), .ZN(n6400) );
  NAND2_X2 U5791 ( .A1(n4867), .A2(n3505), .ZN(n6261) );
  NAND3_X1 U5792 ( .A1(n5586), .A2(n5587), .A3(n5584), .ZN(n4790) );
  INV_X4 U5793 ( .A(n5063), .ZN(n5068) );
  NAND2_X4 U5794 ( .A1(regWrData[7]), .A2(n3787), .ZN(n3788) );
  NAND2_X4 U5795 ( .A1(n5322), .A2(n3788), .ZN(n6486) );
  XNOR2_X2 U5796 ( .A(n3789), .B(n7029), .ZN(net221813) );
  OAI21_X1 U5797 ( .B1(n3207), .B2(net224851), .A(n2838), .ZN(n7107) );
  NAND2_X2 U5798 ( .A1(n5707), .A2(n5976), .ZN(n5665) );
  NAND2_X4 U5799 ( .A1(n5081), .A2(n5082), .ZN(n5083) );
  NAND2_X2 U5800 ( .A1(n7244), .A2(n7246), .ZN(n3791) );
  NAND3_X4 U5801 ( .A1(n7245), .A2(n7247), .A3(n3792), .ZN(n7249) );
  INV_X4 U5802 ( .A(n3791), .ZN(n3792) );
  INV_X4 U5803 ( .A(n6425), .ZN(n7245) );
  NAND2_X4 U5804 ( .A1(n7242), .A2(n7201), .ZN(n7244) );
  NAND2_X2 U5805 ( .A1(n3793), .A2(n4980), .ZN(n4981) );
  NAND3_X1 U5806 ( .A1(n4979), .A2(net224737), .A3(net225047), .ZN(n4980) );
  NAND2_X1 U5807 ( .A1(n5347), .A2(n5334), .ZN(n5121) );
  NAND3_X1 U5809 ( .A1(\wb/dsize_reg/z2 [24]), .A2(net224995), .A3(n5343), 
        .ZN(n5346) );
  NAND3_X2 U5810 ( .A1(\wb/dsize_reg/z2 [24]), .A2(net224991), .A3(n5343), 
        .ZN(n5334) );
  NAND3_X2 U5811 ( .A1(n5213), .A2(n5211), .A3(n5212), .ZN(n3794) );
  NAND3_X2 U5812 ( .A1(n5212), .A2(n5211), .A3(n5213), .ZN(n5933) );
  OAI21_X1 U5813 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4505) );
  INV_X2 U5814 ( .A(n4116), .ZN(n4118) );
  NOR2_X2 U5815 ( .A1(n3995), .A2(n4116), .ZN(n3992) );
  NOR2_X4 U5816 ( .A1(n4715), .A2(net228359), .ZN(n3795) );
  INV_X8 U5817 ( .A(n6261), .ZN(n3939) );
  NAND2_X2 U5818 ( .A1(n3301), .A2(net224861), .ZN(n3797) );
  NAND2_X4 U5819 ( .A1(n3797), .A2(n3798), .ZN(n5430) );
  NAND2_X2 U5820 ( .A1(net228326), .A2(n7725), .ZN(n3799) );
  NAND2_X4 U5821 ( .A1(n5032), .A2(n3799), .ZN(n6570) );
  INV_X1 U5822 ( .A(net224731), .ZN(net228326) );
  NAND2_X4 U5823 ( .A1(n2609), .A2(net230611), .ZN(n3801) );
  NAND2_X4 U5824 ( .A1(n3800), .A2(n3801), .ZN(n7310) );
  NAND4_X4 U5825 ( .A1(n5031), .A2(n5030), .A3(n5028), .A4(n5029), .ZN(n5032)
         );
  INV_X2 U5826 ( .A(n3301), .ZN(n3818) );
  AOI22_X2 U5827 ( .A1(n7123), .A2(n6521), .B1(n3951), .B2(n7310), .ZN(n6377)
         );
  NAND4_X1 U5828 ( .A1(n6640), .A2(n6641), .A3(n6915), .A4(net221163), .ZN(
        n6651) );
  NAND3_X1 U5829 ( .A1(net225237), .A2(reg31Val_0[24]), .A3(net224781), .ZN(
        n4750) );
  NOR3_X2 U5830 ( .A1(net225230), .A2(n3860), .A3(n7562), .ZN(n4822) );
  INV_X1 U5831 ( .A(n6524), .ZN(n5903) );
  NAND2_X2 U5832 ( .A1(n5935), .A2(n6462), .ZN(n6440) );
  NOR2_X4 U5834 ( .A1(n5046), .A2(n3803), .ZN(n5229) );
  OAI21_X1 U5835 ( .B1(n3944), .B2(n6054), .A(n3133), .ZN(n6055) );
  NOR2_X1 U5836 ( .A1(n6050), .A2(n6054), .ZN(n6057) );
  NAND3_X2 U5837 ( .A1(n6378), .A2(n6377), .A3(n6379), .ZN(n3804) );
  INV_X4 U5838 ( .A(n3804), .ZN(n3805) );
  INV_X2 U5839 ( .A(n3350), .ZN(net228280) );
  INV_X16 U5840 ( .A(net224789), .ZN(net224785) );
  NAND3_X2 U5841 ( .A1(n5882), .A2(n5883), .A3(n5884), .ZN(n3806) );
  INV_X4 U5842 ( .A(n3806), .ZN(n3807) );
  AOI21_X1 U5843 ( .B1(n6040), .B2(n5831), .A(n5830), .ZN(n5884) );
  NOR2_X2 U5844 ( .A1(n5850), .A2(n5849), .ZN(n5882) );
  OAI21_X1 U5845 ( .B1(n6635), .B2(n3541), .A(n6633), .ZN(n6636) );
  NOR2_X1 U5846 ( .A1(n7939), .A2(n3541), .ZN(n6463) );
  NAND3_X2 U5847 ( .A1(n6626), .A2(n6627), .A3(n3123), .ZN(\ex_mem/N204 ) );
  NAND2_X2 U5848 ( .A1(n3612), .A2(n3924), .ZN(n3809) );
  OAI21_X2 U5849 ( .B1(net224833), .B2(n6585), .A(n6584), .ZN(n6628) );
  AOI21_X1 U5850 ( .B1(n6583), .B2(n6582), .A(n6581), .ZN(n6629) );
  INV_X8 U5851 ( .A(net220646), .ZN(net221758) );
  INV_X8 U5852 ( .A(n3170), .ZN(n5993) );
  AOI21_X1 U5853 ( .B1(n5779), .B2(n4971), .A(n4970), .ZN(n5743) );
  NAND2_X4 U5855 ( .A1(n6522), .A2(n5949), .ZN(n7172) );
  NAND2_X4 U5856 ( .A1(net220865), .A2(n6897), .ZN(n6905) );
  INV_X1 U5857 ( .A(n5218), .ZN(n3810) );
  INV_X2 U5858 ( .A(n3810), .ZN(n3811) );
  NAND3_X2 U5859 ( .A1(net33205), .A2(n3069), .A3(n2704), .ZN(net220517) );
  NAND2_X4 U5860 ( .A1(n7306), .A2(n7305), .ZN(n7307) );
  NAND3_X2 U5861 ( .A1(\wb/dsize_reg/z2 [1]), .A2(n4856), .A3(net225214), .ZN(
        n5584) );
  NAND2_X4 U5862 ( .A1(n4331), .A2(iAddr[6]), .ZN(n4332) );
  OAI211_X4 U5863 ( .C1(n4108), .C2(n3895), .A(n4107), .B(n4106), .ZN(iAddr[6]) );
  INV_X1 U5864 ( .A(n4978), .ZN(n4979) );
  NOR2_X1 U5865 ( .A1(n7557), .A2(n3290), .ZN(n5668) );
  NAND2_X2 U5866 ( .A1(n5941), .A2(n6462), .ZN(n6470) );
  INV_X8 U5867 ( .A(n6933), .ZN(n6934) );
  OAI211_X4 U5868 ( .C1(n3914), .C2(n3151), .A(n6099), .B(n6170), .ZN(n6835)
         );
  NOR2_X2 U5869 ( .A1(n7743), .A2(net224897), .ZN(\ex_mem/N140 ) );
  NAND2_X2 U5870 ( .A1(n6583), .A2(n5972), .ZN(n5987) );
  AOI21_X2 U5871 ( .B1(n5732), .B2(n5967), .A(n5954), .ZN(n5261) );
  OAI21_X1 U5872 ( .B1(n4817), .B2(n4816), .A(net224915), .ZN(n4818) );
  INV_X1 U5873 ( .A(n7232), .ZN(n3822) );
  INV_X2 U5874 ( .A(n3822), .ZN(n3823) );
  INV_X2 U5875 ( .A(n6032), .ZN(n6037) );
  INV_X8 U5876 ( .A(n4171), .ZN(n4173) );
  INV_X8 U5877 ( .A(n6947), .ZN(n6432) );
  NAND2_X4 U5878 ( .A1(n5044), .A2(n5469), .ZN(n5912) );
  NAND2_X2 U5879 ( .A1(n6838), .A2(n2842), .ZN(n7296) );
  INV_X4 U5882 ( .A(net228148), .ZN(net228149) );
  INV_X2 U5883 ( .A(n4266), .ZN(n4268) );
  OAI21_X1 U5884 ( .B1(n4233), .B2(n4200), .A(n4187), .ZN(n4192) );
  INV_X8 U5885 ( .A(n4233), .ZN(n4249) );
  NAND2_X1 U5886 ( .A1(n7127), .A2(n6540), .ZN(n5923) );
  OAI221_X4 U5887 ( .B1(n5461), .B2(n5462), .C1(n5459), .C2(n5460), .A(n5458), 
        .ZN(n5465) );
  NAND3_X2 U5888 ( .A1(reg31Val_0[17]), .A2(net224781), .A3(net224991), .ZN(
        n5650) );
  NAND3_X2 U5889 ( .A1(reg31Val_0[1]), .A2(net224781), .A3(net225045), .ZN(
        n5587) );
  NAND3_X2 U5890 ( .A1(net224781), .A2(reg31Val_0[15]), .A3(net224991), .ZN(
        n4944) );
  NAND3_X2 U5891 ( .A1(reg31Val_0[28]), .A2(net225237), .A3(net224781), .ZN(
        n4928) );
  NOR3_X1 U5892 ( .A1(net223209), .A2(n7564), .A3(net228276), .ZN(n4956) );
  INV_X2 U5894 ( .A(n3434), .ZN(n4255) );
  NOR2_X2 U5895 ( .A1(n4865), .A2(n2729), .ZN(n4740) );
  NOR2_X4 U5896 ( .A1(n5577), .A2(n5576), .ZN(n5581) );
  OAI22_X2 U5897 ( .A1(n7530), .A2(n3912), .B1(n7691), .B2(n3909), .ZN(n5578)
         );
  NOR2_X2 U5898 ( .A1(n3901), .A2(n7540), .ZN(n4730) );
  INV_X8 U5899 ( .A(n6075), .ZN(n6105) );
  OAI221_X4 U5900 ( .B1(n7702), .B2(n2578), .C1(n3942), .C2(n5110), .A(n5109), 
        .ZN(n6348) );
  NAND3_X2 U5901 ( .A1(n5347), .A2(n5344), .A3(n5120), .ZN(n5331) );
  NAND2_X4 U5902 ( .A1(net225520), .A2(net228018), .ZN(n4887) );
  OAI21_X1 U5903 ( .B1(net224833), .B2(n5817), .A(n5816), .ZN(n5818) );
  NAND2_X4 U5904 ( .A1(n4149), .A2(n4085), .ZN(n4335) );
  INV_X8 U5905 ( .A(n4467), .ZN(n4341) );
  NAND2_X4 U5906 ( .A1(n5007), .A2(net225238), .ZN(n3826) );
  INV_X8 U5907 ( .A(n5539), .ZN(n5551) );
  OAI211_X4 U5908 ( .C1(n5538), .C2(n5537), .A(n5536), .B(n5535), .ZN(n5539)
         );
  BUF_X32 U5910 ( .A(n5204), .Z(n3827) );
  AOI22_X4 U5911 ( .A1(n4727), .A2(net225047), .B1(n2634), .B2(net225047), 
        .ZN(n5152) );
  INV_X1 U5912 ( .A(n2842), .ZN(n3828) );
  NAND2_X2 U5914 ( .A1(n7044), .A2(n5869), .ZN(n5988) );
  NAND3_X2 U5915 ( .A1(n3916), .A2(n5869), .A3(n2759), .ZN(n5870) );
  INV_X4 U5916 ( .A(net228093), .ZN(net228094) );
  NAND2_X2 U5917 ( .A1(n6392), .A2(n6391), .ZN(n3831) );
  NAND2_X4 U5918 ( .A1(n3829), .A2(n3830), .ZN(n3832) );
  NAND2_X4 U5919 ( .A1(n3831), .A2(n3832), .ZN(n6870) );
  NAND2_X4 U5921 ( .A1(n3833), .A2(n3834), .ZN(n3836) );
  NAND2_X4 U5922 ( .A1(n3836), .A2(n3835), .ZN(n5337) );
  INV_X4 U5923 ( .A(n5329), .ZN(n3834) );
  NOR2_X1 U5924 ( .A1(net229037), .A2(n6120), .ZN(n6119) );
  NOR2_X1 U5925 ( .A1(net224955), .A2(n6333), .ZN(\id_ex/N38 ) );
  INV_X1 U5926 ( .A(net228029), .ZN(net228074) );
  NOR2_X2 U5928 ( .A1(n4288), .A2(n4522), .ZN(n4289) );
  NOR2_X2 U5929 ( .A1(net228697), .A2(net224783), .ZN(n4713) );
  XNOR2_X2 U5930 ( .A(n5307), .B(net224865), .ZN(n3838) );
  NOR3_X2 U5931 ( .A1(n6984), .A2(n3672), .A3(n2645), .ZN(n6981) );
  NAND2_X4 U5932 ( .A1(n6406), .A2(n6405), .ZN(n6880) );
  NAND2_X4 U5933 ( .A1(n4544), .A2(n4510), .ZN(n4513) );
  AOI21_X4 U5934 ( .B1(n3223), .B2(n3985), .A(n4138), .ZN(n3986) );
  NAND3_X2 U5935 ( .A1(n4823), .A2(net228074), .A3(n4856), .ZN(n4826) );
  INV_X1 U5937 ( .A(n7960), .ZN(n3839) );
  INV_X1 U5938 ( .A(n3475), .ZN(n4760) );
  OAI22_X1 U5939 ( .A1(n2699), .A2(n7938), .B1(n2700), .B2(n5417), .ZN(n4841)
         );
  NOR2_X2 U5940 ( .A1(n2699), .A2(n5383), .ZN(n5378) );
  INV_X1 U5941 ( .A(n3698), .ZN(n6527) );
  NAND2_X4 U5942 ( .A1(n5020), .A2(n5771), .ZN(n5751) );
  INV_X8 U5943 ( .A(n6758), .ZN(n6755) );
  NAND2_X4 U5944 ( .A1(n5526), .A2(n5522), .ZN(n5548) );
  INV_X2 U5945 ( .A(n5522), .ZN(n5525) );
  OAI211_X2 U5947 ( .C1(n7057), .C2(n3482), .A(n7055), .B(n3532), .ZN(n7064)
         );
  NAND3_X2 U5948 ( .A1(n5087), .A2(n5088), .A3(n5308), .ZN(n4716) );
  NAND2_X4 U5949 ( .A1(n4389), .A2(n4011), .ZN(n4392) );
  NAND2_X4 U5950 ( .A1(n4385), .A2(n2775), .ZN(n4387) );
  NOR3_X1 U5951 ( .A1(n4320), .A2(n4250), .A3(n3169), .ZN(n4251) );
  NOR2_X2 U5952 ( .A1(n6525), .A2(n5904), .ZN(n5909) );
  INV_X8 U5953 ( .A(n7014), .ZN(n7006) );
  NAND3_X4 U5954 ( .A1(n7006), .A2(n7910), .A3(n7005), .ZN(n7019) );
  OAI21_X2 U5955 ( .B1(n7014), .B2(n7013), .A(n7012), .ZN(n7021) );
  NAND2_X4 U5956 ( .A1(n7010), .A2(net228159), .ZN(n7014) );
  NAND2_X2 U5957 ( .A1(net223346), .A2(net225091), .ZN(n4929) );
  NOR3_X2 U5958 ( .A1(n3082), .A2(net224787), .A3(net225238), .ZN(n4894) );
  INV_X8 U5959 ( .A(net223348), .ZN(net228018) );
  NAND3_X4 U5960 ( .A1(n7241), .A2(n3947), .A3(n5239), .ZN(n5960) );
  NOR2_X1 U5961 ( .A1(n7293), .A2(n3950), .ZN(n6781) );
  INV_X1 U5962 ( .A(n3566), .ZN(n7184) );
  XNOR2_X2 U5963 ( .A(n7177), .B(n3242), .ZN(n7290) );
  NAND3_X2 U5964 ( .A1(n7001), .A2(n3571), .A3(n3842), .ZN(n7341) );
  INV_X4 U5965 ( .A(n3841), .ZN(n3842) );
  NOR2_X2 U5966 ( .A1(n6910), .A2(n6927), .ZN(n6912) );
  NAND2_X4 U5967 ( .A1(n6920), .A2(n6886), .ZN(n6926) );
  NAND2_X4 U5969 ( .A1(n5719), .A2(n5718), .ZN(n5835) );
  OAI22_X1 U5971 ( .A1(n7522), .A2(n3912), .B1(n7706), .B2(n3909), .ZN(n5398)
         );
  OAI22_X1 U5972 ( .A1(n7541), .A2(n3912), .B1(n7700), .B2(n3909), .ZN(n5563)
         );
  OAI22_X1 U5973 ( .A1(n7705), .A2(n3909), .B1(n7528), .B2(n3912), .ZN(n5713)
         );
  OAI22_X1 U5974 ( .A1(n7523), .A2(n3911), .B1(n7703), .B2(n3909), .ZN(n5402)
         );
  NAND2_X2 U5975 ( .A1(n4868), .A2(n7476), .ZN(n5685) );
  NAND2_X4 U5976 ( .A1(n5972), .A2(n6788), .ZN(n5977) );
  INV_X8 U5977 ( .A(n4332), .ZN(n4442) );
  OAI211_X4 U5978 ( .C1(n4115), .C2(n3896), .A(n4114), .B(n4113), .ZN(iAddr[2]) );
  INV_X1 U5979 ( .A(n7248), .ZN(n3847) );
  INV_X2 U5980 ( .A(net33276), .ZN(net35542) );
  INV_X4 U5981 ( .A(net228479), .ZN(net227982) );
  NAND3_X1 U5982 ( .A1(net224787), .A2(n2619), .A3(\wb/dsize_reg/z2 [17]), 
        .ZN(n4937) );
  INV_X16 U5983 ( .A(net224785), .ZN(net224783) );
  NOR2_X2 U5984 ( .A1(n7098), .A2(n3918), .ZN(n6832) );
  NOR2_X2 U5985 ( .A1(n7098), .A2(n3923), .ZN(n7068) );
  NAND2_X1 U5986 ( .A1(n6424), .A2(n5972), .ZN(n6430) );
  OAI21_X4 U5987 ( .B1(n2940), .B2(n5986), .A(n5985), .ZN(n3850) );
  AOI21_X1 U5989 ( .B1(n6638), .B2(n3428), .A(n6636), .ZN(n6658) );
  AOI21_X1 U5990 ( .B1(net224843), .B2(n2628), .A(net224835), .ZN(n6635) );
  NOR2_X2 U5991 ( .A1(n3869), .A2(net224895), .ZN(\ex_mem/N128 ) );
  INV_X16 U5992 ( .A(n3919), .ZN(n3920) );
  INV_X4 U5993 ( .A(net228809), .ZN(net220849) );
  OAI21_X1 U5994 ( .B1(net224745), .B2(n3179), .A(n6381), .ZN(n6384) );
  INV_X8 U5995 ( .A(n4770), .ZN(n5002) );
  NAND3_X2 U5996 ( .A1(n4804), .A2(n4803), .A3(net225251), .ZN(n5437) );
  NOR2_X2 U5998 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  OAI211_X4 U5999 ( .C1(n7920), .C2(n7201), .A(n6443), .B(n5936), .ZN(n6129)
         );
  NAND3_X4 U6000 ( .A1(n6450), .A2(n3874), .A3(n3947), .ZN(n6003) );
  INV_X1 U6002 ( .A(net220895), .ZN(net221765) );
  NAND3_X1 U6003 ( .A1(n5034), .A2(n5490), .A3(n5035), .ZN(n4817) );
  BUF_X32 U6004 ( .A(n5006), .Z(n3853) );
  NAND3_X2 U6005 ( .A1(net229330), .A2(net220865), .A3(n2910), .ZN(n6417) );
  NAND3_X2 U6006 ( .A1(n2910), .A2(net229330), .A3(n3701), .ZN(n6415) );
  NAND2_X4 U6007 ( .A1(n6414), .A2(n6415), .ZN(net221424) );
  NAND2_X4 U6008 ( .A1(n2653), .A2(n6748), .ZN(n6799) );
  NAND2_X4 U6009 ( .A1(n4156), .A2(n4134), .ZN(n4149) );
  NAND3_X2 U6010 ( .A1(n4041), .A2(n4102), .A3(n4069), .ZN(n3997) );
  NAND3_X2 U6011 ( .A1(n4068), .A2(n4069), .A3(n4070), .ZN(n4071) );
  OAI21_X1 U6012 ( .B1(n7466), .B2(n7501), .A(n4270), .ZN(n4030) );
  NAND2_X1 U6013 ( .A1(n7127), .A2(n7968), .ZN(n7042) );
  INV_X16 U6014 ( .A(n3904), .ZN(n3905) );
  INV_X2 U6015 ( .A(net221491), .ZN(net223329) );
  NOR3_X1 U6016 ( .A1(n6356), .A2(n6355), .A3(net221491), .ZN(n6363) );
  NAND2_X1 U6017 ( .A1(n7358), .A2(net221491), .ZN(net221490) );
  NOR2_X2 U6018 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  NAND2_X1 U6019 ( .A1(n7201), .A2(n5984), .ZN(n5262) );
  NAND2_X4 U6020 ( .A1(n5984), .A2(n3862), .ZN(n5985) );
  NAND3_X2 U6021 ( .A1(n5467), .A2(net224731), .A3(n5043), .ZN(n5044) );
  OAI21_X1 U6022 ( .B1(n3818), .B2(net224851), .A(n2838), .ZN(n6567) );
  NAND2_X4 U6023 ( .A1(net229628), .A2(net225601), .ZN(n6882) );
  XNOR2_X1 U6024 ( .A(n4427), .B(n2771), .ZN(n4428) );
  XNOR2_X1 U6025 ( .A(n4392), .B(n4391), .ZN(n4393) );
  XNOR2_X1 U6026 ( .A(n2986), .B(n4396), .ZN(n4397) );
  OAI21_X1 U6027 ( .B1(n7111), .B2(n3781), .A(n7109), .ZN(n7121) );
  NAND2_X4 U6028 ( .A1(n5148), .A2(n5147), .ZN(n7110) );
  NAND2_X4 U6029 ( .A1(n5976), .A2(n5707), .ZN(n5231) );
  NAND2_X4 U6031 ( .A1(n4769), .A2(n4768), .ZN(n4770) );
  INV_X16 U6032 ( .A(n5706), .ZN(n3908) );
  NAND2_X4 U6033 ( .A1(n5026), .A2(net225047), .ZN(n5268) );
  NAND2_X4 U6034 ( .A1(n5274), .A2(n5275), .ZN(n6185) );
  NAND2_X4 U6035 ( .A1(n4814), .A2(net225047), .ZN(n5033) );
  NAND2_X4 U6036 ( .A1(n5006), .A2(n5005), .ZN(n5012) );
  AOI21_X1 U6037 ( .B1(n3946), .B2(regWrData[0]), .A(n2647), .ZN(n6299) );
  NOR2_X1 U6038 ( .A1(n5064), .A2(n5063), .ZN(n4761) );
  OAI211_X4 U6039 ( .C1(n6034), .C2(n6033), .A(n6032), .B(n6985), .ZN(n5512)
         );
  NAND3_X2 U6040 ( .A1(n4848), .A2(n4847), .A3(\wb/dsize_reg/z2 [26]), .ZN(
        n4849) );
  AOI21_X1 U6041 ( .B1(n4799), .B2(n3853), .A(net224903), .ZN(\ex_mem/N102 )
         );
  INV_X1 U6042 ( .A(n3827), .ZN(n4728) );
  NAND3_X2 U6043 ( .A1(n6414), .A2(n6415), .A3(n6417), .ZN(n6416) );
  NAND2_X4 U6044 ( .A1(n5153), .A2(n5152), .ZN(n5204) );
  OAI211_X2 U6046 ( .C1(n6459), .C2(n6460), .A(n3862), .B(n7242), .ZN(n6475)
         );
  NAND2_X4 U6047 ( .A1(n5039), .A2(n5492), .ZN(n6721) );
  NAND2_X4 U6048 ( .A1(n3654), .A2(n7044), .ZN(net220885) );
  NAND3_X4 U6049 ( .A1(n5955), .A2(n5957), .A3(n5956), .ZN(n6622) );
  XNOR2_X1 U6050 ( .A(n3141), .B(n4413), .ZN(n4414) );
  NAND2_X2 U6051 ( .A1(n3988), .A2(n3999), .ZN(n4053) );
  INV_X8 U6052 ( .A(n3999), .ZN(n4046) );
  NAND2_X4 U6053 ( .A1(n4544), .A2(n4515), .ZN(n4518) );
  OAI21_X2 U6054 ( .B1(n3815), .B2(n5990), .A(n7202), .ZN(n5991) );
  NAND2_X4 U6055 ( .A1(n6733), .A2(n5893), .ZN(n6489) );
  NAND3_X2 U6056 ( .A1(n2615), .A2(n3222), .A3(n6825), .ZN(n5888) );
  NAND2_X4 U6057 ( .A1(n5047), .A2(n5048), .ZN(n5049) );
  INV_X8 U6058 ( .A(n4358), .ZN(n4500) );
  XNOR2_X2 U6059 ( .A(n7440), .B(n7431), .ZN(n3993) );
  NAND2_X1 U6060 ( .A1(n6568), .A2(n6462), .ZN(n5276) );
  NAND2_X4 U6061 ( .A1(net221929), .A2(n7020), .ZN(n7113) );
  AOI211_X1 U6062 ( .C1(n7919), .C2(regWrData[4]), .A(n4997), .B(n4998), .ZN(
        n4771) );
  AOI22_X4 U6063 ( .A1(n4766), .A2(net224993), .B1(n4765), .B2(net224993), 
        .ZN(n5114) );
  MUX2_X2 U6064 ( .A(n3569), .B(n2901), .S(net227828), .Z(n6038) );
  NAND2_X4 U6065 ( .A1(n5649), .A2(n7150), .ZN(n7080) );
  NAND3_X2 U6066 ( .A1(n6212), .A2(n6213), .A3(n5298), .ZN(n5599) );
  NAND3_X1 U6067 ( .A1(n3361), .A2(n5451), .A3(n3588), .ZN(n6827) );
  NAND3_X1 U6068 ( .A1(n3762), .A2(n6705), .A3(n3222), .ZN(n6592) );
  INV_X8 U6069 ( .A(n6823), .ZN(n6594) );
  AOI21_X1 U6070 ( .B1(n3467), .B2(n3470), .A(net224903), .ZN(\ex_mem/N120 )
         );
  NAND2_X4 U6071 ( .A1(n7227), .A2(n7226), .ZN(n5858) );
  NAND2_X4 U6072 ( .A1(n5895), .A2(n5894), .ZN(n6549) );
  NAND2_X4 U6073 ( .A1(n3127), .A2(n4722), .ZN(n4723) );
  NAND3_X2 U6074 ( .A1(n4912), .A2(n4913), .A3(n4914), .ZN(n5183) );
  NAND2_X4 U6075 ( .A1(n3394), .A2(net228942), .ZN(n6906) );
  OAI211_X4 U6076 ( .C1(n6905), .C2(n3359), .A(n6904), .B(n6903), .ZN(n6914)
         );
  INV_X8 U6077 ( .A(n4356), .ZN(n4355) );
  NOR3_X1 U6078 ( .A1(n4232), .A2(n4318), .A3(n3169), .ZN(n4007) );
  NAND3_X4 U6079 ( .A1(n4486), .A2(n4344), .A3(iAddr[16]), .ZN(n4345) );
  NAND2_X4 U6080 ( .A1(n3990), .A2(n4458), .ZN(n4117) );
  NAND2_X4 U6081 ( .A1(n3867), .A2(n4802), .ZN(n4772) );
  OAI21_X1 U6082 ( .B1(n6370), .B2(net224851), .A(n2838), .ZN(net221492) );
  NAND2_X4 U6083 ( .A1(n6124), .A2(net220780), .ZN(n7241) );
  NAND2_X2 U6084 ( .A1(n7331), .A2(n7325), .ZN(n7277) );
  INV_X8 U6085 ( .A(n6591), .ZN(n7297) );
  NAND2_X4 U6086 ( .A1(n6586), .A2(n7297), .ZN(n6704) );
  NOR2_X1 U6087 ( .A1(net224955), .A2(n6321), .ZN(\id_ex/N40 ) );
  NAND3_X4 U6088 ( .A1(n5393), .A2(n5395), .A3(n5394), .ZN(n5803) );
  NOR3_X4 U6089 ( .A1(n5392), .A2(n5391), .A3(n5390), .ZN(n5393) );
  INV_X8 U6090 ( .A(net35037), .ZN(net224789) );
  INV_X32 U6091 ( .A(net225049), .ZN(net225045) );
  OAI21_X1 U6093 ( .B1(net224833), .B2(n4972), .A(net222371), .ZN(n5742) );
  OAI21_X1 U6094 ( .B1(net222371), .B2(net224851), .A(n2838), .ZN(n4971) );
  NAND2_X4 U6095 ( .A1(n3795), .A2(net230143), .ZN(n5013) );
  NAND2_X4 U6096 ( .A1(n6679), .A2(n2599), .ZN(n6838) );
  NAND2_X4 U6097 ( .A1(n6045), .A2(n6046), .ZN(n5927) );
  NAND2_X4 U6099 ( .A1(n3643), .A2(memAddr[2]), .ZN(n4987) );
  INV_X16 U6100 ( .A(n3906), .ZN(n3907) );
  INV_X16 U6101 ( .A(net223262), .ZN(net225237) );
  INV_X1 U6102 ( .A(n3907), .ZN(n3946) );
  NOR3_X1 U6103 ( .A1(n7059), .A2(n7060), .A3(n3776), .ZN(n7065) );
  NAND2_X4 U6104 ( .A1(net223348), .A2(net225096), .ZN(n5296) );
  AOI21_X4 U6105 ( .B1(n7233), .B2(n7232), .A(n3923), .ZN(n7234) );
  INV_X8 U6106 ( .A(n5513), .ZN(n5839) );
  INV_X1 U6107 ( .A(n5577), .ZN(n4797) );
  INV_X8 U6108 ( .A(n5296), .ZN(n3900) );
  INV_X8 U6109 ( .A(n6932), .ZN(n3861) );
  INV_X16 U6110 ( .A(n3861), .ZN(n3862) );
  NAND4_X4 U6111 ( .A1(n3573), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(
        net221416) );
  OAI21_X1 U6112 ( .B1(n6571), .B2(n3301), .A(n6569), .ZN(n6572) );
  NAND3_X4 U6113 ( .A1(n2598), .A2(n4784), .A3(net224787), .ZN(n5256) );
  INV_X8 U6114 ( .A(n7212), .ZN(n7252) );
  NAND4_X4 U6115 ( .A1(n6199), .A2(n6197), .A3(n6198), .A4(n6196), .ZN(n7212)
         );
  NAND2_X1 U6116 ( .A1(n7019), .A2(net220714), .ZN(n7023) );
  INV_X8 U6117 ( .A(n6089), .ZN(n3863) );
  NAND2_X4 U6118 ( .A1(n3785), .A2(net230143), .ZN(n3865) );
  INV_X4 U6119 ( .A(n7552), .ZN(n3866) );
  INV_X16 U6120 ( .A(n3866), .ZN(n3867) );
  OAI222_X2 U6122 ( .A1(n6236), .A2(n2937), .B1(n2735), .B2(n2699), .C1(
        net35052), .C2(n3252), .ZN(regWrData[19]) );
  INV_X1 U6123 ( .A(n3713), .ZN(n4923) );
  NAND3_X2 U6124 ( .A1(n6731), .A2(n6732), .A3(n3690), .ZN(n6822) );
  OAI211_X1 U6125 ( .C1(n6594), .C2(n3690), .A(n6593), .B(n6592), .ZN(n6595)
         );
  NAND2_X4 U6126 ( .A1(n6113), .A2(n6114), .ZN(n6141) );
  NOR3_X2 U6127 ( .A1(n3864), .A2(n2737), .A3(n3899), .ZN(n4726) );
  OAI211_X4 U6128 ( .C1(n3712), .C2(n5871), .A(n2678), .B(n3856), .ZN(n6933)
         );
  NOR2_X1 U6129 ( .A1(net228087), .A2(net224871), .ZN(n5321) );
  NAND2_X1 U6130 ( .A1(n7358), .A2(n3568), .ZN(n5913) );
  NOR2_X1 U6131 ( .A1(n6349), .A2(n3568), .ZN(n6353) );
  INV_X1 U6132 ( .A(n3568), .ZN(n5885) );
  NOR2_X1 U6133 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  NAND3_X2 U6134 ( .A1(n6152), .A2(n5813), .A3(n3413), .ZN(n6154) );
  INV_X8 U6137 ( .A(n5256), .ZN(n5356) );
  NAND2_X4 U6138 ( .A1(n3295), .A2(net220885), .ZN(n7002) );
  NOR2_X4 U6139 ( .A1(n3849), .A2(net225102), .ZN(n4784) );
  NAND2_X4 U6140 ( .A1(n5365), .A2(n6810), .ZN(n6706) );
  NAND2_X4 U6141 ( .A1(n5007), .A2(net225238), .ZN(n5015) );
  OAI21_X1 U6142 ( .B1(iAddr[16]), .B2(n3136), .A(n4482), .ZN(n4481) );
  INV_X2 U6143 ( .A(n4481), .ZN(n4706) );
  XNOR2_X1 U6144 ( .A(iAddr[17]), .B(n4482), .ZN(n4705) );
  INV_X8 U6145 ( .A(n6902), .ZN(n3868) );
  INV_X8 U6146 ( .A(n6872), .ZN(n6902) );
  NAND2_X4 U6147 ( .A1(n6974), .A2(net225029), .ZN(net220775) );
  NAND3_X2 U6148 ( .A1(net227982), .A2(n3646), .A3(net220663), .ZN(n6161) );
  NAND2_X4 U6149 ( .A1(n5363), .A2(n5364), .ZN(n6817) );
  OAI21_X1 U6150 ( .B1(net224833), .B2(n6097), .A(n3485), .ZN(n6136) );
  OAI21_X1 U6151 ( .B1(n3485), .B2(net224851), .A(n2838), .ZN(n6096) );
  XNOR2_X1 U6152 ( .A(n3485), .B(net224865), .ZN(n6393) );
  NAND3_X2 U6154 ( .A1(n5263), .A2(n5262), .A3(n5261), .ZN(n6616) );
  OAI211_X4 U6155 ( .C1(n4264), .C2(n4265), .A(n4263), .B(n4262), .ZN(
        iAddr[24]) );
  NOR3_X2 U6156 ( .A1(net225226), .A2(n2736), .A3(net230622), .ZN(n4731) );
  INV_X32 U6157 ( .A(net225243), .ZN(net223245) );
  BUF_X32 U6158 ( .A(n5080), .Z(n3869) );
  NAND4_X4 U6159 ( .A1(n5737), .A2(n5736), .A3(n5739), .A4(n5738), .ZN(n7133)
         );
  INV_X8 U6160 ( .A(n5108), .ZN(n5976) );
  INV_X1 U6161 ( .A(net228858), .ZN(net223337) );
  NAND2_X4 U6162 ( .A1(n5228), .A2(n5229), .ZN(n5230) );
  NAND2_X2 U6163 ( .A1(n4740), .A2(n4856), .ZN(n4742) );
  AND2_X2 U6164 ( .A1(n7073), .A2(n7997), .ZN(n3873) );
  NAND3_X2 U6165 ( .A1(n5145), .A2(n5146), .A3(net224731), .ZN(n5148) );
  NAND2_X1 U6166 ( .A1(n3725), .A2(n3722), .ZN(n6467) );
  NAND2_X1 U6167 ( .A1(n5048), .A2(n7924), .ZN(n4966) );
  BUF_X32 U6168 ( .A(n3732), .Z(n3875) );
  NAND4_X4 U6169 ( .A1(n5877), .A2(n5880), .A3(n5878), .A4(n5879), .ZN(n7126)
         );
  NAND4_X2 U6170 ( .A1(n4276), .A2(n4290), .A3(n4293), .A4(n4277), .ZN(n4278)
         );
  OAI22_X4 U6171 ( .A1(n7458), .A2(n7509), .B1(n4325), .B2(n4247), .ZN(n4239)
         );
  AOI21_X4 U6172 ( .B1(n4022), .B2(n4021), .A(n4020), .ZN(n4325) );
  OAI211_X4 U6173 ( .C1(n4286), .C2(n3895), .A(n4285), .B(n4284), .ZN(n7906)
         );
  BUF_X32 U6174 ( .A(n6174), .Z(n3876) );
  NAND2_X4 U6175 ( .A1(n5663), .A2(n5662), .ZN(n6946) );
  INV_X4 U6176 ( .A(n3751), .ZN(n3888) );
  NAND2_X4 U6177 ( .A1(n5137), .A2(n3880), .ZN(n5140) );
  NAND2_X4 U6178 ( .A1(n5129), .A2(n5128), .ZN(n5454) );
  XNOR2_X1 U6179 ( .A(n7508), .B(n2863), .ZN(n4406) );
  XNOR2_X1 U6180 ( .A(n7419), .B(n4423), .ZN(n4424) );
  XNOR2_X1 U6181 ( .A(n7431), .B(n4451), .ZN(n4452) );
  NAND2_X1 U6182 ( .A1(n4423), .A2(n4415), .ZN(n4425) );
  NAND2_X4 U6184 ( .A1(n5102), .A2(n5443), .ZN(n6741) );
  NOR2_X4 U6186 ( .A1(n3525), .A2(n3796), .ZN(n5207) );
  INV_X4 U6187 ( .A(n5041), .ZN(n6174) );
  NAND2_X2 U6189 ( .A1(n2790), .A2(n2696), .ZN(n6517) );
  NAND2_X4 U6190 ( .A1(n5863), .A2(n7941), .ZN(n6602) );
  INV_X2 U6191 ( .A(n7198), .ZN(n7200) );
  NAND2_X4 U6192 ( .A1(n7861), .A2(n3726), .ZN(n4358) );
  NAND2_X4 U6193 ( .A1(n3967), .A2(n2770), .ZN(n3968) );
  NAND2_X4 U6194 ( .A1(n5241), .A2(n5240), .ZN(n5876) );
  AOI21_X2 U6195 ( .B1(n6944), .B2(n6431), .A(n5708), .ZN(n5241) );
  NAND3_X2 U6196 ( .A1(n5989), .A2(n3916), .A3(n5886), .ZN(n5674) );
  NAND3_X2 U6198 ( .A1(n2683), .A2(\wb/dsize_reg/z2 [29]), .A3(net224991), 
        .ZN(n5522) );
  NAND4_X1 U6199 ( .A1(n3121), .A2(net228697), .A3(net224993), .A4(n7921), 
        .ZN(n4936) );
  NAND3_X2 U6200 ( .A1(n2683), .A2(\wb/dsize_reg/z2 [25]), .A3(net225216), 
        .ZN(n5585) );
  OAI222_X2 U6202 ( .A1(n7571), .A2(net225015), .B1(n2731), .B2(n3933), .C1(
        n3935), .C2(n2951), .ZN(regWrData[31]) );
  NAND3_X1 U6203 ( .A1(n3661), .A2(n6888), .A3(n3665), .ZN(n6143) );
  NAND2_X4 U6204 ( .A1(n5368), .A2(n5440), .ZN(n5172) );
  AOI22_X4 U6205 ( .A1(net223245), .A2(n2709), .B1(n3643), .B2(memAddr[28]), 
        .ZN(n4932) );
  NAND2_X4 U6206 ( .A1(n5692), .A2(n6458), .ZN(n5833) );
  NAND2_X4 U6207 ( .A1(n7046), .A2(net225029), .ZN(n7048) );
  NAND2_X4 U6208 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X4 U6209 ( .A1(n4891), .A2(n4890), .ZN(n4892) );
  INV_X2 U6210 ( .A(n5323), .ZN(n5126) );
  NAND3_X1 U6211 ( .A1(n5310), .A2(n5309), .A3(n5308), .ZN(n5316) );
  INV_X2 U6212 ( .A(net220319), .ZN(net221792) );
  AOI21_X1 U6213 ( .B1(n5043), .B2(n2600), .A(net224903), .ZN(\ex_mem/N113 )
         );
  INV_X2 U6214 ( .A(n5912), .ZN(n5918) );
  AOI21_X1 U6215 ( .B1(net224843), .B2(n5912), .A(net224835), .ZN(n5915) );
  OAI21_X1 U6216 ( .B1(n7033), .B2(n7032), .A(n7031), .ZN(n7034) );
  NAND2_X4 U6217 ( .A1(n7030), .A2(net225029), .ZN(n7032) );
  AOI211_X4 U6218 ( .C1(n4889), .C2(net225214), .A(net223300), .B(n4888), .ZN(
        n4891) );
  NOR2_X1 U6219 ( .A1(net229071), .A2(n2949), .ZN(n4823) );
  NOR3_X1 U6220 ( .A1(net228029), .A2(n7561), .A3(net223348), .ZN(n4830) );
  INV_X2 U6221 ( .A(n3696), .ZN(n4780) );
  OAI21_X1 U6222 ( .B1(net224745), .B2(n3696), .A(n6811), .ZN(n6814) );
  INV_X8 U6223 ( .A(n6706), .ZN(n6702) );
  INV_X4 U6224 ( .A(net225053), .ZN(net225051) );
  NAND2_X1 U6225 ( .A1(n3454), .A2(n7239), .ZN(n6666) );
  NAND3_X2 U6226 ( .A1(n6664), .A2(n6665), .A3(n6666), .ZN(n7040) );
  NAND3_X2 U6227 ( .A1(n5196), .A2(n3355), .A3(n5197), .ZN(n5201) );
  OAI21_X1 U6228 ( .B1(n6530), .B2(n3698), .A(n3629), .ZN(n5908) );
  NAND2_X4 U6229 ( .A1(n5431), .A2(n6526), .ZN(n5432) );
  INV_X16 U6230 ( .A(n5297), .ZN(n3898) );
  NAND3_X2 U6231 ( .A1(n6961), .A2(n6960), .A3(n6959), .ZN(n6962) );
  NAND2_X4 U6232 ( .A1(n6876), .A2(n6879), .ZN(n6892) );
  NAND2_X4 U6233 ( .A1(n6879), .A2(n6880), .ZN(n6889) );
  NAND2_X4 U6234 ( .A1(n6871), .A2(n6874), .ZN(n6879) );
  NAND2_X4 U6235 ( .A1(n6870), .A2(n6869), .ZN(n6874) );
  MUX2_X2 U6236 ( .A(n5372), .B(n7746), .S(net225434), .Z(n5794) );
  AOI21_X1 U6237 ( .B1(net224953), .B2(n2915), .A(n4633), .ZN(n4631) );
  AOI21_X1 U6238 ( .B1(net224955), .B2(n2928), .A(n4633), .ZN(n4629) );
  AOI21_X1 U6239 ( .B1(net224953), .B2(n2913), .A(n4633), .ZN(n4627) );
  AOI21_X1 U6240 ( .B1(net224953), .B2(n2898), .A(n4633), .ZN(n4625) );
  AOI21_X1 U6241 ( .B1(net224953), .B2(n2905), .A(n4633), .ZN(n4623) );
  AOI21_X1 U6242 ( .B1(net224953), .B2(n2923), .A(n4633), .ZN(n4621) );
  OAI21_X1 U6243 ( .B1(n3566), .B2(net224851), .A(n2838), .ZN(n7178) );
  NAND2_X1 U6244 ( .A1(n5302), .A2(n3566), .ZN(n7192) );
  NAND2_X1 U6245 ( .A1(n5723), .A2(n3566), .ZN(n7213) );
  NOR2_X1 U6246 ( .A1(net224859), .A2(n3566), .ZN(n6778) );
  NAND2_X4 U6247 ( .A1(n6067), .A2(n7027), .ZN(n6915) );
  NAND2_X4 U6248 ( .A1(n4361), .A2(n4544), .ZN(n4362) );
  NAND4_X4 U6249 ( .A1(n4053), .A2(n4051), .A3(n4052), .A4(n4060), .ZN(n4349)
         );
  OAI211_X4 U6250 ( .C1(n4244), .C2(n3895), .A(n4243), .B(n4242), .ZN(n7857)
         );
  NAND2_X1 U6251 ( .A1(n4953), .A2(net225047), .ZN(n4955) );
  NAND2_X1 U6252 ( .A1(n5667), .A2(net225047), .ZN(n6258) );
  XNOR2_X1 U6253 ( .A(n7512), .B(n3552), .ZN(n4398) );
  NOR2_X1 U6254 ( .A1(n7511), .A2(n7512), .ZN(n3966) );
  NOR3_X1 U6255 ( .A1(n4320), .A2(n3169), .A3(n4319), .ZN(n4321) );
  OAI21_X1 U6256 ( .B1(n4319), .B2(n3150), .A(n4184), .ZN(n4186) );
  NOR2_X1 U6257 ( .A1(n4319), .A2(n4207), .ZN(n4197) );
  NOR2_X1 U6258 ( .A1(n4245), .A2(n4319), .ZN(n4253) );
  NOR2_X1 U6259 ( .A1(n4250), .A2(n4319), .ZN(n4235) );
  NOR2_X2 U6260 ( .A1(n6615), .A2(n6614), .ZN(n6627) );
  INV_X8 U6261 ( .A(net221648), .ZN(net225003) );
  OAI211_X4 U6262 ( .C1(n4231), .C2(n3896), .A(n4230), .B(n4229), .ZN(n7859)
         );
  INV_X2 U6263 ( .A(n7134), .ZN(n5924) );
  NAND2_X1 U6264 ( .A1(n7358), .A2(n7134), .ZN(n7163) );
  NOR2_X1 U6265 ( .A1(n6335), .A2(n7134), .ZN(n6336) );
  NOR2_X1 U6266 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  NAND3_X1 U6267 ( .A1(n3352), .A2(net228869), .A3(n3653), .ZN(n6988) );
  NOR2_X1 U6268 ( .A1(n7242), .A2(n7156), .ZN(n5251) );
  NAND2_X4 U6269 ( .A1(n7134), .A2(net225029), .ZN(n7156) );
  NAND2_X4 U6270 ( .A1(n6348), .A2(net225029), .ZN(n5914) );
  INV_X16 U6271 ( .A(n5167), .ZN(n5972) );
  NAND2_X4 U6272 ( .A1(net225013), .A2(n2976), .ZN(n6031) );
  NAND2_X4 U6273 ( .A1(net221802), .A2(n6118), .ZN(net221793) );
  NAND2_X4 U6274 ( .A1(n5796), .A2(n5797), .ZN(n6156) );
  NAND3_X1 U6275 ( .A1(n3407), .A2(n2594), .A3(n5036), .ZN(n4816) );
  OAI21_X1 U6276 ( .B1(n6722), .B2(n3764), .A(n6720), .ZN(n6723) );
  NAND4_X2 U6277 ( .A1(n6558), .A2(n6698), .A3(n5906), .A4(n5905), .ZN(n6528)
         );
  NAND2_X1 U6278 ( .A1(n6698), .A2(n3615), .ZN(n6491) );
  NAND3_X4 U6279 ( .A1(n3534), .A2(n5888), .A3(n5792), .ZN(n6698) );
  NAND2_X4 U6280 ( .A1(n7272), .A2(n7271), .ZN(net220293) );
  NAND3_X2 U6281 ( .A1(n5981), .A2(n5980), .A3(n5979), .ZN(n7175) );
  NAND2_X4 U6282 ( .A1(n3734), .A2(n3283), .ZN(net222840) );
  NAND2_X4 U6283 ( .A1(net220644), .A2(net225587), .ZN(n6895) );
  INV_X4 U6284 ( .A(n6941), .ZN(n6942) );
  NAND2_X4 U6285 ( .A1(n6683), .A2(n3838), .ZN(n6825) );
  AOI22_X4 U6286 ( .A1(n4733), .A2(net225214), .B1(n4732), .B2(net225214), 
        .ZN(n5146) );
  NAND2_X1 U6287 ( .A1(net223346), .A2(net225091), .ZN(n4777) );
  NAND3_X1 U6288 ( .A1(n7607), .A2(net225091), .A3(net225096), .ZN(n5005) );
  OAI211_X4 U6289 ( .C1(n5724), .C2(n5947), .A(n5734), .B(n5664), .ZN(n6514)
         );
  NAND2_X4 U6290 ( .A1(n3921), .A2(n7220), .ZN(n7237) );
  XNOR2_X1 U6291 ( .A(n7297), .B(n6012), .ZN(n6022) );
  OAI22_X1 U6292 ( .A1(n2842), .A2(n7289), .B1(n7297), .B2(n2622), .ZN(n7291)
         );
  NAND2_X1 U6293 ( .A1(n7288), .A2(n7297), .ZN(n7289) );
  NAND4_X1 U6294 ( .A1(net225622), .A2(net225605), .A3(n7719), .A4(n7254), 
        .ZN(n5730) );
  NAND2_X1 U6295 ( .A1(net225622), .A2(n3069), .ZN(n5658) );
  NAND2_X4 U6296 ( .A1(n4509), .A2(n4508), .ZN(n4504) );
  INV_X8 U6297 ( .A(n4360), .ZN(n4509) );
  NAND2_X4 U6298 ( .A1(n3984), .A2(n3982), .ZN(n4142) );
  OAI211_X4 U6299 ( .C1(n4219), .C2(n3895), .A(n4218), .B(n4217), .ZN(n7861)
         );
  NAND3_X2 U6300 ( .A1(n6485), .A2(n5896), .A3(n3133), .ZN(n5431) );
  NAND3_X1 U6302 ( .A1(n7859), .A2(iAddr[23]), .A3(iAddr[24]), .ZN(n4514) );
  NAND2_X1 U6303 ( .A1(n7859), .A2(iAddr[24]), .ZN(n4532) );
  NAND2_X1 U6304 ( .A1(n3681), .A2(n4165), .ZN(n4170) );
  AOI21_X1 U6305 ( .B1(n3682), .B2(n4348), .A(n4167), .ZN(n4168) );
  NOR2_X1 U6306 ( .A1(n4166), .A2(n3682), .ZN(n4167) );
  NOR3_X1 U6307 ( .A1(n3682), .A2(n4247), .A3(n4246), .ZN(n4252) );
  NOR3_X1 U6308 ( .A1(n3681), .A2(n3169), .A3(n4233), .ZN(n4234) );
  INV_X2 U6309 ( .A(n2585), .ZN(n5925) );
  NOR3_X1 U6310 ( .A1(n6350), .A2(n6815), .A3(n2585), .ZN(n6352) );
  OAI21_X1 U6311 ( .B1(n7076), .B2(net220651), .A(n7075), .ZN(n7077) );
  NAND2_X1 U6312 ( .A1(n7358), .A2(n2585), .ZN(n7075) );
  NAND2_X1 U6313 ( .A1(reg31Val_0[9]), .A2(n3937), .ZN(n6241) );
  NOR2_X1 U6314 ( .A1(n7242), .A2(net220651), .ZN(n5961) );
  NAND2_X1 U6315 ( .A1(net220651), .A2(n3269), .ZN(n6145) );
  INV_X2 U6316 ( .A(net220651), .ZN(net220656) );
  NAND2_X4 U6317 ( .A1(n7074), .A2(net225029), .ZN(net220651) );
  NAND3_X1 U6318 ( .A1(reg31Val_0[27]), .A2(n3937), .A3(n6105), .ZN(n6111) );
  INV_X8 U6319 ( .A(n5807), .ZN(n7057) );
  NAND2_X1 U6320 ( .A1(n6621), .A2(n7239), .ZN(n6133) );
  NOR3_X2 U6321 ( .A1(n7344), .A2(n7343), .A3(n2602), .ZN(net220297) );
  NAND2_X4 U6322 ( .A1(n6888), .A2(net221766), .ZN(net220895) );
  NAND2_X4 U6323 ( .A1(n6140), .A2(n6394), .ZN(net221165) );
  NAND3_X2 U6324 ( .A1(n4341), .A2(iAddr[9]), .A3(iAddr[10]), .ZN(n4472) );
  AOI21_X1 U6325 ( .B1(n4042), .B2(n4102), .A(n2668), .ZN(n3998) );
  NOR2_X2 U6326 ( .A1(n7429), .A2(n7428), .ZN(n3956) );
  NAND2_X4 U6327 ( .A1(n5839), .A2(n3727), .ZN(n6911) );
  NAND2_X4 U6328 ( .A1(n3197), .A2(n5487), .ZN(n7143) );
  NAND2_X4 U6329 ( .A1(n5488), .A2(n7143), .ZN(n7053) );
  OAI21_X1 U6330 ( .B1(net224833), .B2(n5832), .A(n2633), .ZN(n5883) );
  OAI21_X1 U6331 ( .B1(n2633), .B2(net224851), .A(n2838), .ZN(n5831) );
  NAND2_X4 U6332 ( .A1(n6039), .A2(n6040), .ZN(net221818) );
  NAND2_X4 U6333 ( .A1(n5778), .A2(n5779), .ZN(net220632) );
  NOR2_X2 U6334 ( .A1(n3821), .A2(net220753), .ZN(n6982) );
  NAND2_X4 U6335 ( .A1(n5207), .A2(n6174), .ZN(n5161) );
  NAND2_X4 U6336 ( .A1(n5189), .A2(n5190), .ZN(n6382) );
  NAND2_X4 U6337 ( .A1(n5728), .A2(n5729), .ZN(n6540) );
  NAND4_X4 U6338 ( .A1(n4342), .A2(n4339), .A3(n4341), .A4(n4340), .ZN(n4343)
         );
  NAND3_X2 U6339 ( .A1(n4437), .A2(n4436), .A3(n4435), .ZN(iAddr[11]) );
  NAND2_X4 U6340 ( .A1(n4487), .A2(iAddr[18]), .ZN(n4503) );
  NAND2_X1 U6341 ( .A1(n6246), .A2(n7945), .ZN(regWrData[12]) );
  NAND3_X2 U6342 ( .A1(n6245), .A2(n3743), .A3(n6246), .ZN(n5274) );
  NAND2_X4 U6344 ( .A1(n3734), .A2(net224787), .ZN(n5359) );
  OAI211_X4 U6345 ( .C1(n2972), .C2(n7205), .A(n6434), .B(n6433), .ZN(n7248)
         );
  OAI211_X4 U6346 ( .C1(n7252), .C2(n3914), .A(n7250), .B(n7251), .ZN(n7270)
         );
  NAND2_X4 U6347 ( .A1(n7248), .A2(n7249), .ZN(n7250) );
  NAND3_X2 U6348 ( .A1(n5761), .A2(n7935), .A3(n5760), .ZN(n6659) );
  INV_X1 U6349 ( .A(n3711), .ZN(n6563) );
  NAND2_X4 U6350 ( .A1(n3164), .A2(n3163), .ZN(n4407) );
  NAND2_X4 U6351 ( .A1(n4409), .A2(n2776), .ZN(n4427) );
  NAND2_X4 U6352 ( .A1(n6558), .A2(n5812), .ZN(n7055) );
  INV_X8 U6353 ( .A(n5568), .ZN(n4991) );
  OAI211_X1 U6354 ( .C1(net220307), .C2(n7166), .A(net33205), .B(n2839), .ZN(
        net220537) );
  NOR2_X1 U6355 ( .A1(net225622), .A2(net33205), .ZN(n4968) );
  NOR2_X1 U6356 ( .A1(net225083), .A2(net33205), .ZN(n5170) );
  NAND3_X2 U6357 ( .A1(n7283), .A2(n7282), .A3(n2682), .ZN(n7286) );
  INV_X2 U6358 ( .A(n6549), .ZN(n6701) );
  NAND2_X4 U6359 ( .A1(n5842), .A2(net221494), .ZN(net220889) );
  NAND2_X4 U6360 ( .A1(n5663), .A2(n3402), .ZN(n5167) );
  NAND3_X4 U6361 ( .A1(n7271), .A2(n7238), .A3(n7237), .ZN(net220292) );
  NAND2_X4 U6363 ( .A1(n7112), .A2(n3653), .ZN(n6372) );
  NAND3_X2 U6364 ( .A1(n5997), .A2(n3947), .A3(n5996), .ZN(n7256) );
  NAND2_X4 U6365 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  INV_X8 U6367 ( .A(n5645), .ZN(n5810) );
  NAND2_X4 U6368 ( .A1(n5861), .A2(n5862), .ZN(n6728) );
  AOI22_X4 U6369 ( .A1(n7176), .A2(n3172), .B1(n6661), .B2(n6620), .ZN(n5861)
         );
  INV_X8 U6370 ( .A(n5140), .ZN(n5663) );
  NAND2_X4 U6371 ( .A1(n5897), .A2(n5907), .ZN(n5541) );
  NAND2_X4 U6372 ( .A1(n5401), .A2(n5400), .ZN(n5897) );
  NAND2_X4 U6373 ( .A1(n5428), .A2(n5429), .ZN(n5907) );
  NOR3_X4 U6374 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(n7316) );
  NAND3_X2 U6375 ( .A1(net220403), .A2(n7275), .A3(net229367), .ZN(n7276) );
  XNOR2_X2 U6376 ( .A(n7116), .B(n7910), .ZN(n7117) );
  AOI22_X4 U6377 ( .A1(n6651), .A2(n6650), .B1(n6649), .B2(n6648), .ZN(n6652)
         );
  NAND2_X4 U6378 ( .A1(n6913), .A2(n7341), .ZN(net220540) );
  NAND2_X4 U6379 ( .A1(n5430), .A2(n6568), .ZN(n6526) );
  AOI21_X1 U6380 ( .B1(n6973), .B2(n2838), .A(n7997), .ZN(n6978) );
  AOI21_X1 U6381 ( .B1(net224843), .B2(n7997), .A(net224833), .ZN(n6976) );
  INV_X4 U6382 ( .A(net35036), .ZN(net225101) );
  OAI221_X4 U6383 ( .B1(n6201), .B2(n6672), .C1(n6619), .C2(n2703), .A(n6200), 
        .ZN(n6803) );
  NAND2_X1 U6384 ( .A1(n5967), .A2(n6431), .ZN(n5968) );
  NAND3_X2 U6385 ( .A1(n6431), .A2(n7169), .A3(n3955), .ZN(n6434) );
  NAND3_X1 U6386 ( .A1(n7181), .A2(n5662), .A3(n5663), .ZN(n5997) );
  NOR2_X2 U6387 ( .A1(net220539), .A2(net220540), .ZN(n7167) );
  OAI21_X1 U6388 ( .B1(n7145), .B2(n7144), .A(n3652), .ZN(n7146) );
  NAND2_X1 U6389 ( .A1(n7144), .A2(n3672), .ZN(n7135) );
  NAND2_X4 U6390 ( .A1(n5809), .A2(n3652), .ZN(n6043) );
  OAI211_X4 U6391 ( .C1(n3689), .C2(n6688), .A(n5337), .B(n5451), .ZN(n5891)
         );
  NAND2_X4 U6392 ( .A1(n5707), .A2(n5976), .ZN(n6466) );
  INV_X16 U6393 ( .A(net225216), .ZN(net223242) );
  NAND3_X2 U6394 ( .A1(n6623), .A2(n6624), .A3(n6625), .ZN(n7039) );
  NAND2_X4 U6395 ( .A1(n3794), .A2(n7255), .ZN(n7171) );
  INV_X2 U6396 ( .A(n7112), .ZN(n7114) );
  NAND2_X4 U6397 ( .A1(n6155), .A2(n3413), .ZN(n6032) );
  NAND2_X4 U6398 ( .A1(n5435), .A2(n6153), .ZN(n6033) );
  INV_X8 U6399 ( .A(n6395), .ZN(n3919) );
  MUX2_X2 U6400 ( .A(n3247), .B(reg31Val_0[2]), .S(net224725), .Z(n1979) );
  XNOR2_X1 U6401 ( .A(n4431), .B(n2769), .ZN(n4432) );
  XNOR2_X1 U6402 ( .A(n4407), .B(n2770), .ZN(n4408) );
  XNOR2_X1 U6403 ( .A(n4411), .B(n2921), .ZN(n4412) );
  NOR2_X1 U6404 ( .A1(n3247), .A2(n3531), .ZN(n4451) );
  NOR3_X1 U6405 ( .A1(n4401), .A2(n7511), .A3(n7512), .ZN(n4402) );
  XOR2_X1 U6406 ( .A(n3247), .B(n3531), .Z(n4457) );
  XNOR2_X1 U6407 ( .A(n7438), .B(n3247), .ZN(n4111) );
  NAND2_X4 U6408 ( .A1(n6175), .A2(net225029), .ZN(n6188) );
  NAND2_X4 U6409 ( .A1(n5170), .A2(n6861), .ZN(n7193) );
  NAND2_X4 U6410 ( .A1(n5708), .A2(n3862), .ZN(n5969) );
  INV_X8 U6411 ( .A(n5734), .ZN(n5708) );
  NAND2_X4 U6412 ( .A1(n7242), .A2(n7255), .ZN(n5734) );
  INV_X16 U6413 ( .A(n6946), .ZN(n6462) );
  NAND2_X4 U6415 ( .A1(n7115), .A2(net221759), .ZN(net220646) );
  NAND2_X4 U6416 ( .A1(n3630), .A2(n3233), .ZN(n6929) );
  NAND2_X4 U6417 ( .A1(net220312), .A2(net220313), .ZN(n7318) );
  NAND2_X4 U6418 ( .A1(n5317), .A2(n3449), .ZN(n6075) );
  NAND4_X4 U6419 ( .A1(n7314), .A2(n7313), .A3(n7312), .A4(n7311), .ZN(n7317)
         );
  NAND2_X4 U6420 ( .A1(n2671), .A2(net224787), .ZN(n6089) );
  NAND2_X4 U6421 ( .A1(n5463), .A2(n3812), .ZN(n7056) );
  NAND2_X4 U6422 ( .A1(n6911), .A2(n7020), .ZN(n7001) );
  NAND2_X4 U6423 ( .A1(n5975), .A2(n5976), .ZN(n5717) );
  NAND3_X2 U6424 ( .A1(n5105), .A2(n5106), .A3(n5107), .ZN(n5108) );
  OAI211_X4 U6425 ( .C1(n5983), .C2(n7201), .A(n5982), .B(n7170), .ZN(n7253)
         );
  OAI21_X1 U6426 ( .B1(net229367), .B2(n3950), .A(n6082), .ZN(n6083) );
  NAND2_X4 U6427 ( .A1(n4254), .A2(n4258), .ZN(n4276) );
  OAI22_X4 U6428 ( .A1(n7459), .A2(n7508), .B1(n3139), .B2(n4246), .ZN(n4254)
         );
  XNOR2_X1 U6429 ( .A(n3174), .B(n4418), .ZN(n4419) );
  NAND2_X1 U6430 ( .A1(n4151), .A2(n3438), .ZN(n4159) );
  NAND2_X1 U6432 ( .A1(n3438), .A2(n4152), .ZN(n4155) );
  XNOR2_X1 U6433 ( .A(n7445), .B(n3174), .ZN(n4084) );
  NAND3_X2 U6434 ( .A1(n4153), .A2(n4152), .A3(n4083), .ZN(n4139) );
  NOR2_X2 U6435 ( .A1(n7445), .A2(n7426), .ZN(n4067) );
  NAND2_X4 U6436 ( .A1(net224925), .A2(n2941), .ZN(n4465) );
  NAND2_X4 U6437 ( .A1(n4633), .A2(n4632), .ZN(n4652) );
  INV_X32 U6438 ( .A(n3898), .ZN(n3899) );
  NAND2_X4 U6439 ( .A1(net223346), .A2(net225091), .ZN(n5297) );
  INV_X32 U6440 ( .A(net225237), .ZN(net225238) );
  INV_X32 U6441 ( .A(n3900), .ZN(n3901) );
  NAND2_X4 U6442 ( .A1(net224785), .A2(net225102), .ZN(n4925) );
  INV_X32 U6443 ( .A(n3908), .ZN(n3909) );
  NAND2_X4 U6444 ( .A1(n7496), .A2(n7476), .ZN(n5706) );
  INV_X8 U6445 ( .A(n5685), .ZN(n3910) );
  INV_X16 U6446 ( .A(n3910), .ZN(n3911) );
  INV_X16 U6447 ( .A(n3911), .ZN(n5709) );
  INV_X32 U6448 ( .A(n3915), .ZN(n3916) );
  INV_X32 U6449 ( .A(n3916), .ZN(n7242) );
  NAND2_X4 U6450 ( .A1(n6790), .A2(n6965), .ZN(n7205) );
  INV_X8 U6451 ( .A(n7244), .ZN(n7169) );
  NAND2_X4 U6452 ( .A1(n3724), .A2(n6965), .ZN(n6672) );
  NAND2_X4 U6453 ( .A1(n5934), .A2(n5933), .ZN(n7202) );
  INV_X32 U6454 ( .A(net225049), .ZN(net225047) );
  INV_X32 U6455 ( .A(net225053), .ZN(net225049) );
  INV_X32 U6456 ( .A(net224997), .ZN(net224993) );
  INV_X32 U6459 ( .A(net224953), .ZN(net224943) );
  INV_X32 U6460 ( .A(net224937), .ZN(net224955) );
  INV_X32 U6461 ( .A(n3949), .ZN(n3947) );
  INV_X32 U6462 ( .A(net224865), .ZN(net224861) );
  INV_X32 U6463 ( .A(net224741), .ZN(net224735) );
  INV_X32 U6464 ( .A(net224741), .ZN(net224737) );
  INV_X32 U6466 ( .A(net224749), .ZN(net224745) );
  INV_X4 U6468 ( .A(n4383), .ZN(n3960) );
  INV_X4 U6470 ( .A(n4387), .ZN(n3962) );
  INV_X4 U6472 ( .A(n4392), .ZN(n3964) );
  INV_X4 U6473 ( .A(n4407), .ZN(n3967) );
  INV_X4 U6474 ( .A(n4427), .ZN(n3969) );
  XNOR2_X2 U6475 ( .A(n3972), .B(n7400), .ZN(n3973) );
  XNOR2_X2 U6476 ( .A(\mem/addImm/mux_map1/M3/z2[31] ), .B(n7400), .ZN(n4031)
         );
  XNOR2_X2 U6477 ( .A(n7466), .B(n7501), .ZN(n4267) );
  INV_X4 U6478 ( .A(n4267), .ZN(n4029) );
  XNOR2_X2 U6479 ( .A(n7456), .B(n7511), .ZN(n4233) );
  XNOR2_X2 U6480 ( .A(n7455), .B(n7512), .ZN(n4319) );
  INV_X4 U6481 ( .A(n4319), .ZN(n3975) );
  XNOR2_X2 U6482 ( .A(n7460), .B(n7507), .ZN(n4260) );
  XNOR2_X2 U6483 ( .A(n7459), .B(n7508), .ZN(n4246) );
  XNOR2_X2 U6484 ( .A(n7451), .B(n7516), .ZN(n4250) );
  XNOR2_X2 U6485 ( .A(n7458), .B(n7509), .ZN(n4247) );
  INV_X4 U6486 ( .A(n4247), .ZN(n4329) );
  XNOR2_X2 U6487 ( .A(n7457), .B(n7510), .ZN(n4188) );
  NAND2_X2 U6488 ( .A1(n4329), .A2(n4021), .ZN(n4232) );
  XNOR2_X2 U6489 ( .A(n7452), .B(n7515), .ZN(n4037) );
  INV_X4 U6490 ( .A(n7452), .ZN(n3976) );
  NAND2_X2 U6491 ( .A1(n4391), .A2(n3976), .ZN(n4165) );
  NAND2_X2 U6492 ( .A1(n4037), .A2(n4165), .ZN(n4348) );
  XNOR2_X2 U6493 ( .A(n7453), .B(n7514), .ZN(n4248) );
  NAND2_X2 U6494 ( .A1(n4348), .A2(n4346), .ZN(n4318) );
  XNOR2_X2 U6495 ( .A(n7454), .B(n7513), .ZN(n4356) );
  XNOR2_X2 U6496 ( .A(n7447), .B(n7519), .ZN(n3977) );
  INV_X4 U6497 ( .A(n3977), .ZN(n4337) );
  NAND2_X2 U6498 ( .A1(n2744), .A2(n2996), .ZN(n4083) );
  NAND2_X2 U6499 ( .A1(n4382), .A2(n2997), .ZN(n3983) );
  NAND2_X2 U6500 ( .A1(n4417), .A2(n2998), .ZN(n4081) );
  NAND2_X2 U6501 ( .A1(n3983), .A2(n4081), .ZN(n3978) );
  INV_X4 U6502 ( .A(n3978), .ZN(n4000) );
  XNOR2_X2 U6503 ( .A(n7449), .B(n7518), .ZN(n4047) );
  XNOR2_X2 U6504 ( .A(n7448), .B(n7425), .ZN(n4151) );
  INV_X4 U6505 ( .A(n4151), .ZN(n3982) );
  XNOR2_X2 U6506 ( .A(n7444), .B(n7427), .ZN(n4082) );
  INV_X4 U6507 ( .A(n3983), .ZN(n4138) );
  OAI21_X4 U6508 ( .B1(n3987), .B2(n4142), .A(n3986), .ZN(n3999) );
  XNOR2_X2 U6509 ( .A(n7441), .B(n7419), .ZN(n4042) );
  XNOR2_X2 U6510 ( .A(n7442), .B(n7429), .ZN(n4045) );
  NAND2_X2 U6511 ( .A1(n2793), .A2(n2999), .ZN(n4069) );
  INV_X4 U6513 ( .A(n4463), .ZN(n3990) );
  NAND2_X2 U6514 ( .A1(reg31Val_3[1]), .A2(n3093), .ZN(n4119) );
  INV_X4 U6515 ( .A(n3993), .ZN(n4131) );
  OAI21_X4 U6516 ( .B1(n4110), .B2(n4072), .A(n3161), .ZN(n4041) );
  INV_X4 U6517 ( .A(n4070), .ZN(n3996) );
  AOI21_X4 U6518 ( .B1(n3997), .B2(n3998), .A(n3996), .ZN(n4051) );
  NAND2_X2 U6519 ( .A1(n2775), .A2(n3000), .ZN(n4052) );
  NAND2_X2 U6520 ( .A1(n2768), .A2(n3001), .ZN(n4060) );
  INV_X4 U6521 ( .A(n4047), .ZN(n4144) );
  XNOR2_X2 U6522 ( .A(n7443), .B(n7428), .ZN(n4075) );
  INV_X4 U6523 ( .A(n4075), .ZN(n4090) );
  NAND2_X2 U6524 ( .A1(n4144), .A2(n4090), .ZN(n4003) );
  OAI21_X4 U6525 ( .B1(n4046), .B2(n4003), .A(n4052), .ZN(n4005) );
  XNOR2_X2 U6526 ( .A(n7450), .B(n7517), .ZN(n4049) );
  INV_X4 U6527 ( .A(n4049), .ZN(n4004) );
  OAI21_X4 U6528 ( .B1(n4006), .B2(n4005), .A(n4004), .ZN(n4050) );
  INV_X4 U6529 ( .A(n4260), .ZN(n4258) );
  NAND2_X2 U6530 ( .A1(n2778), .A2(n3002), .ZN(n4184) );
  NAND2_X2 U6534 ( .A1(n4013), .A2(n4012), .ZN(n4209) );
  INV_X4 U6535 ( .A(n4209), .ZN(n4016) );
  INV_X4 U6536 ( .A(n7454), .ZN(n4014) );
  NAND2_X2 U6537 ( .A1(n4396), .A2(n4014), .ZN(n4212) );
  INV_X4 U6538 ( .A(n4212), .ZN(n4015) );
  AOI21_X4 U6539 ( .B1(n4016), .B2(n4355), .A(n4015), .ZN(n4017) );
  OAI21_X4 U6540 ( .B1(n4019), .B2(n4018), .A(n4017), .ZN(n4183) );
  NAND2_X2 U6541 ( .A1(n2762), .A2(n3097), .ZN(n4187) );
  INV_X4 U6542 ( .A(n4188), .ZN(n4021) );
  NAND2_X2 U6543 ( .A1(n2769), .A2(n3003), .ZN(n4025) );
  NAND2_X2 U6544 ( .A1(n2774), .A2(n3004), .ZN(n4293) );
  NAND2_X2 U6545 ( .A1(n4025), .A2(n4293), .ZN(n4024) );
  NAND2_X2 U6546 ( .A1(n2776), .A2(n3005), .ZN(n4302) );
  NAND2_X2 U6547 ( .A1(n2770), .A2(n3006), .ZN(n4291) );
  NAND2_X2 U6548 ( .A1(n2771), .A2(n3007), .ZN(n4520) );
  NAND2_X2 U6549 ( .A1(n4520), .A2(n4302), .ZN(n4275) );
  XNOR2_X2 U6550 ( .A(n7463), .B(n7504), .ZN(n4523) );
  INV_X4 U6551 ( .A(n4523), .ZN(n4521) );
  XNOR2_X2 U6552 ( .A(n7462), .B(n7505), .ZN(n4222) );
  NAND2_X2 U6553 ( .A1(n4222), .A2(n4520), .ZN(n4304) );
  OAI211_X2 U6554 ( .C1(n2725), .C2(n4275), .A(n4521), .B(n4304), .ZN(n4287)
         );
  XNOR2_X2 U6555 ( .A(n7464), .B(n7503), .ZN(n4292) );
  INV_X4 U6556 ( .A(n4025), .ZN(n4280) );
  XNOR2_X2 U6557 ( .A(n7465), .B(n7502), .ZN(n4282) );
  INV_X4 U6558 ( .A(n4282), .ZN(n4026) );
  OAI21_X4 U6559 ( .B1(n4028), .B2(n4027), .A(n2994), .ZN(n4266) );
  XNOR2_X2 U6560 ( .A(n4031), .B(n4030), .ZN(n4035) );
  INV_X4 U6561 ( .A(n4250), .ZN(n4347) );
  OAI21_X4 U6562 ( .B1(n4178), .B2(n4238), .A(n4036), .ZN(n4171) );
  NAND2_X2 U6563 ( .A1(n3897), .A2(n3098), .ZN(n4038) );
  NAND2_X2 U6564 ( .A1(net224915), .A2(n3043), .ZN(n4059) );
  NAND2_X2 U6565 ( .A1(n4069), .A2(n4041), .ZN(n4093) );
  INV_X4 U6566 ( .A(n4042), .ZN(n4094) );
  INV_X4 U6567 ( .A(n4102), .ZN(n4043) );
  OAI211_X2 U6569 ( .C1(n4057), .C2(n4056), .A(n2684), .B(n4524), .ZN(n4058)
         );
  OAI21_X4 U6570 ( .B1(n4066), .B2(n3895), .A(n4065), .ZN(iAddr[15]) );
  INV_X4 U6571 ( .A(n4071), .ZN(n4074) );
  NAND3_X2 U6572 ( .A1(n4074), .A2(n4117), .A3(n4073), .ZN(n4080) );
  NAND2_X2 U6573 ( .A1(n4074), .A2(n3224), .ZN(n4079) );
  AOI21_X4 U6574 ( .B1(n4077), .B2(n4076), .A(n4075), .ZN(n4078) );
  NAND3_X4 U6575 ( .A1(n4080), .A2(n4079), .A3(n4078), .ZN(n4088) );
  INV_X4 U6576 ( .A(n4082), .ZN(n4099) );
  INV_X4 U6577 ( .A(n4084), .ZN(n4134) );
  NAND2_X2 U6578 ( .A1(net224915), .A2(n3063), .ZN(n4086) );
  NAND2_X2 U6579 ( .A1(net224919), .A2(n3058), .ZN(n4092) );
  OAI211_X2 U6580 ( .C1(n4090), .C2(n4089), .A(n4088), .B(n4524), .ZN(n4091)
         );
  NAND2_X2 U6581 ( .A1(n3897), .A2(n3099), .ZN(n4097) );
  OAI211_X2 U6582 ( .C1(n4094), .C2(n4093), .A(n4524), .B(n4103), .ZN(n4096)
         );
  NAND2_X2 U6583 ( .A1(net224915), .A2(n3055), .ZN(n4095) );
  XNOR2_X2 U6584 ( .A(n4099), .B(n4098), .ZN(n4101) );
  NAND2_X2 U6585 ( .A1(n3897), .A2(n3100), .ZN(n4100) );
  OAI221_X2 U6586 ( .B1(n7673), .B2(net224909), .C1(n3895), .C2(n4101), .A(
        n4100), .ZN(iAddr[8]) );
  XNOR2_X2 U6587 ( .A(n4105), .B(n4104), .ZN(n4108) );
  NAND2_X2 U6588 ( .A1(n3897), .A2(n3101), .ZN(n4107) );
  NAND2_X2 U6589 ( .A1(net224915), .A2(n3059), .ZN(n4106) );
  INV_X4 U6590 ( .A(n4119), .ZN(n4109) );
  XNOR2_X2 U6591 ( .A(n4112), .B(n4111), .ZN(n4115) );
  NAND2_X2 U6592 ( .A1(net224913), .A2(n3062), .ZN(n4113) );
  NAND2_X2 U6593 ( .A1(net224913), .A2(n3061), .ZN(n4123) );
  INV_X4 U6594 ( .A(n4126), .ZN(n4129) );
  XNOR2_X2 U6595 ( .A(n4131), .B(n4130), .ZN(n4133) );
  NAND2_X2 U6596 ( .A1(net224913), .A2(n3060), .ZN(n4132) );
  NAND2_X2 U6597 ( .A1(n3897), .A2(n3102), .ZN(n4137) );
  NAND2_X2 U6598 ( .A1(net224915), .A2(n3057), .ZN(n4135) );
  XNOR2_X2 U6599 ( .A(n4144), .B(n4143), .ZN(n4147) );
  NAND2_X2 U6600 ( .A1(n3897), .A2(n3103), .ZN(n4146) );
  NAND2_X2 U6601 ( .A1(net224919), .A2(n3065), .ZN(n4145) );
  NAND2_X2 U6602 ( .A1(n3897), .A2(n3104), .ZN(n4163) );
  OAI21_X4 U6603 ( .B1(n4160), .B2(n4159), .A(n4158), .ZN(n4162) );
  NAND2_X2 U6604 ( .A1(net224919), .A2(n3056), .ZN(n4161) );
  NAND3_X4 U6605 ( .A1(n4163), .A2(n4162), .A3(n4161), .ZN(iAddr[12]) );
  NAND2_X2 U6606 ( .A1(n3897), .A2(n3105), .ZN(n4176) );
  NAND2_X2 U6607 ( .A1(n4346), .A2(n4164), .ZN(n4172) );
  INV_X4 U6608 ( .A(n4165), .ZN(n4166) );
  OAI221_X2 U6609 ( .B1(n4173), .B2(n4172), .C1(n4171), .C2(n4170), .A(n4169), 
        .ZN(n4175) );
  NAND2_X2 U6610 ( .A1(net224919), .A2(n3066), .ZN(n4174) );
  INV_X4 U6611 ( .A(n4177), .ZN(n4181) );
  NAND2_X2 U6612 ( .A1(n4355), .A2(n4348), .ZN(n4207) );
  INV_X4 U6613 ( .A(n4207), .ZN(n4180) );
  INV_X4 U6614 ( .A(n4179), .ZN(n4198) );
  NAND2_X2 U6616 ( .A1(n4182), .A2(n2942), .ZN(n4196) );
  INV_X4 U6617 ( .A(n4186), .ZN(n4200) );
  NAND2_X2 U6618 ( .A1(net224915), .A2(n3084), .ZN(n4193) );
  NOR2_X4 U6620 ( .A1(n4257), .A2(n4207), .ZN(n4214) );
  INV_X4 U6621 ( .A(n4211), .ZN(n4353) );
  AOI21_X4 U6622 ( .B1(n4214), .B2(n4215), .A(n4213), .ZN(n4216) );
  XNOR2_X2 U6623 ( .A(n4216), .B(n4319), .ZN(n4219) );
  NAND2_X2 U6624 ( .A1(n3897), .A2(n3106), .ZN(n4218) );
  NAND2_X2 U6625 ( .A1(net224919), .A2(n3044), .ZN(n4217) );
  INV_X4 U6626 ( .A(n4222), .ZN(n4220) );
  NOR2_X4 U6627 ( .A1(n4221), .A2(n4220), .ZN(n4227) );
  OAI21_X4 U6628 ( .B1(n4223), .B2(n4222), .A(n4524), .ZN(n4226) );
  NAND2_X2 U6629 ( .A1(n3897), .A2(n3107), .ZN(n4225) );
  NAND2_X2 U6630 ( .A1(net224913), .A2(n3068), .ZN(n4224) );
  NAND2_X2 U6631 ( .A1(n3897), .A2(n3108), .ZN(n4230) );
  NAND2_X2 U6632 ( .A1(net224915), .A2(n3045), .ZN(n4229) );
  INV_X4 U6633 ( .A(n4232), .ZN(n4236) );
  NAND4_X2 U6634 ( .A1(n4236), .A2(n4348), .A3(n4235), .A4(n4234), .ZN(n4237)
         );
  NOR2_X4 U6635 ( .A1(n4238), .A2(n4237), .ZN(n4240) );
  XNOR2_X2 U6636 ( .A(n4241), .B(n4246), .ZN(n4244) );
  NAND2_X2 U6637 ( .A1(n3897), .A2(n3109), .ZN(n4243) );
  NAND2_X2 U6638 ( .A1(net224915), .A2(n3046), .ZN(n4242) );
  INV_X4 U6639 ( .A(n4348), .ZN(n4245) );
  NAND2_X2 U6640 ( .A1(n4021), .A2(n4249), .ZN(n4320) );
  NAND4_X2 U6641 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4349), .ZN(n4256)
         );
  OAI21_X4 U6642 ( .B1(n4256), .B2(n4257), .A(n4255), .ZN(n4259) );
  OAI21_X4 U6643 ( .B1(n4261), .B2(n4260), .A(n4524), .ZN(n4264) );
  NAND2_X2 U6644 ( .A1(n3897), .A2(n3110), .ZN(n4263) );
  NAND2_X2 U6645 ( .A1(net224915), .A2(n3054), .ZN(n4262) );
  NAND2_X2 U6646 ( .A1(n3897), .A2(n3111), .ZN(n4273) );
  NAND2_X2 U6647 ( .A1(n4268), .A2(n4267), .ZN(n4269) );
  NAND3_X2 U6648 ( .A1(n4524), .A2(n4270), .A3(n4269), .ZN(n4272) );
  NAND2_X2 U6649 ( .A1(net224919), .A2(n3047), .ZN(n4271) );
  INV_X4 U6650 ( .A(n4291), .ZN(n4274) );
  NOR2_X4 U6651 ( .A1(n4275), .A2(n4274), .ZN(n4277) );
  INV_X4 U6652 ( .A(n4298), .ZN(n4281) );
  NOR2_X4 U6653 ( .A1(n4281), .A2(n4280), .ZN(n4283) );
  XNOR2_X2 U6654 ( .A(n4283), .B(n4282), .ZN(n4286) );
  NAND2_X2 U6655 ( .A1(n3897), .A2(n3112), .ZN(n4285) );
  NAND2_X2 U6656 ( .A1(net224915), .A2(n3048), .ZN(n4284) );
  INV_X4 U6657 ( .A(n4287), .ZN(n4297) );
  INV_X4 U6658 ( .A(n4520), .ZN(n4522) );
  INV_X4 U6659 ( .A(n4292), .ZN(n4295) );
  INV_X4 U6660 ( .A(n4293), .ZN(n4294) );
  NAND2_X2 U6661 ( .A1(net224919), .A2(n3049), .ZN(n4299) );
  NAND3_X2 U6662 ( .A1(n4303), .A2(n4302), .A3(n4520), .ZN(n4305) );
  XNOR2_X2 U6663 ( .A(n4306), .B(n4523), .ZN(n4310) );
  NAND2_X2 U6664 ( .A1(n3897), .A2(n3113), .ZN(n4525) );
  INV_X4 U6665 ( .A(n4525), .ZN(n4308) );
  NAND2_X2 U6666 ( .A1(net224915), .A2(n3050), .ZN(n4526) );
  INV_X4 U6667 ( .A(n4526), .ZN(n4307) );
  OAI21_X4 U6668 ( .B1(n4310), .B2(n3895), .A(n4309), .ZN(n8108) );
  NAND2_X2 U6669 ( .A1(n7646), .A2(n4666), .ZN(\hazard_detect/eq_83/A[1] ) );
  NAND2_X2 U6670 ( .A1(n7648), .A2(n4666), .ZN(\hazard_detect/eq_83/A[3] ) );
  NAND2_X2 U6671 ( .A1(n7649), .A2(n4666), .ZN(\hazard_detect/eq_83/A[4] ) );
  INV_X4 U6672 ( .A(iAddr[30]), .ZN(n4314) );
  NOR3_X4 U6673 ( .A1(n4317), .A2(n4519), .A3(n4316), .ZN(n4361) );
  NAND2_X2 U6674 ( .A1(net224919), .A2(n3051), .ZN(n4497) );
  NAND2_X2 U6675 ( .A1(n3897), .A2(n3114), .ZN(n4499) );
  INV_X4 U6676 ( .A(n4318), .ZN(n4322) );
  NAND3_X4 U6677 ( .A1(n4498), .A2(n4499), .A3(n4497), .ZN(n4344) );
  NOR2_X4 U6678 ( .A1(n4330), .A2(n4470), .ZN(n4342) );
  INV_X4 U6679 ( .A(iAddr[8]), .ZN(n4443) );
  INV_X4 U6680 ( .A(iAddr[5]), .ZN(n4447) );
  NOR2_X4 U6681 ( .A1(n4443), .A2(n4447), .ZN(n4333) );
  NAND3_X4 U6682 ( .A1(n4333), .A2(n4442), .A3(iAddr[7]), .ZN(n4467) );
  NAND2_X2 U6683 ( .A1(net224919), .A2(n3064), .ZN(n4435) );
  NAND2_X2 U6684 ( .A1(n3897), .A2(n3115), .ZN(n4437) );
  XNOR2_X2 U6685 ( .A(n4336), .B(n3546), .ZN(n4338) );
  NOR2_X4 U6686 ( .A1(n4477), .A2(n4480), .ZN(n4339) );
  NAND2_X2 U6687 ( .A1(net224915), .A2(n3067), .ZN(n4483) );
  NAND2_X2 U6688 ( .A1(n3897), .A2(n3116), .ZN(n4484) );
  AND3_X2 U6689 ( .A1(n4348), .A2(n4347), .A3(n4346), .ZN(n4351) );
  NAND2_X2 U6690 ( .A1(n4353), .A2(n4352), .ZN(n4354) );
  INV_X4 U6691 ( .A(n4354), .ZN(n4357) );
  OAI221_X2 U6692 ( .B1(n4357), .B2(n3169), .C1(n4354), .C2(n4355), .A(n4524), 
        .ZN(n4485) );
  INV_X4 U6693 ( .A(\hazard_detect/eq_83/A[0] ), .ZN(n6291) );
  XNOR2_X2 U6694 ( .A(rd_2[0]), .B(n6291), .ZN(n4367) );
  INV_X4 U6695 ( .A(\hazard_detect/eq_83/A[1] ), .ZN(n4613) );
  XNOR2_X2 U6696 ( .A(rd_2[1]), .B(n4613), .ZN(n4366) );
  NAND2_X2 U6697 ( .A1(valid_2), .A2(n4365), .ZN(n4373) );
  NOR3_X2 U6698 ( .A1(n4367), .A2(n4366), .A3(n4373), .ZN(n4372) );
  INV_X4 U6699 ( .A(\hazard_detect/eq_83/A[4] ), .ZN(n4607) );
  XNOR2_X2 U6700 ( .A(rd_2[4]), .B(n4607), .ZN(n4370) );
  INV_X4 U6701 ( .A(\hazard_detect/eq_83/A[3] ), .ZN(n4609) );
  XNOR2_X2 U6702 ( .A(rd_2[3]), .B(n4609), .ZN(n4369) );
  INV_X4 U6703 ( .A(\hazard_detect/eq_83/A[2] ), .ZN(n4611) );
  XNOR2_X2 U6704 ( .A(rd_2[2]), .B(n4611), .ZN(n4368) );
  NOR3_X2 U6705 ( .A1(n4370), .A2(n4369), .A3(n4368), .ZN(n4371) );
  NAND2_X2 U6706 ( .A1(n4372), .A2(n4371), .ZN(n6321) );
  INV_X4 U6707 ( .A(n6321), .ZN(n4381) );
  XOR2_X2 U6708 ( .A(rs1[0]), .B(rd_2[0]), .Z(n4374) );
  XNOR2_X2 U6709 ( .A(rs1[1]), .B(rd_2[1]), .ZN(n4379) );
  XOR2_X2 U6710 ( .A(rs1[4]), .B(rd_2[4]), .Z(n4377) );
  XOR2_X2 U6711 ( .A(rs1[2]), .B(rd_2[2]), .Z(n4376) );
  XOR2_X2 U6712 ( .A(rs1[3]), .B(rd_2[3]), .Z(n4375) );
  INV_X4 U6713 ( .A(n6333), .ZN(n6280) );
  OAI21_X4 U6714 ( .B1(n4381), .B2(n6280), .A(n2922), .ZN(n4549) );
  NAND2_X2 U6715 ( .A1(n7493), .A2(n7494), .ZN(n6271) );
  NOR2_X4 U6716 ( .A1(n4711), .A2(n3040), .ZN(n4546) );
  MUX2_X2 U6717 ( .A(reg31Val_0[12]), .B(n4384), .S(net224681), .Z(n1919) );
  XNOR2_X2 U6718 ( .A(n7518), .B(n4385), .ZN(n4386) );
  MUX2_X2 U6719 ( .A(reg31Val_0[13]), .B(n4386), .S(net224681), .Z(n1920) );
  MUX2_X2 U6720 ( .A(reg31Val_0[14]), .B(n4388), .S(net224681), .Z(n1926) );
  MUX2_X2 U6721 ( .A(reg31Val_0[15]), .B(n4390), .S(net224681), .Z(n1927) );
  MUX2_X2 U6722 ( .A(reg31Val_0[16]), .B(n4393), .S(net224681), .Z(n1928) );
  MUX2_X2 U6723 ( .A(reg31Val_0[17]), .B(n4395), .S(net224681), .Z(n1929) );
  MUX2_X2 U6724 ( .A(reg31Val_0[18]), .B(n4397), .S(net224681), .Z(n1930) );
  MUX2_X2 U6725 ( .A(reg31Val_0[19]), .B(n4398), .S(net224681), .Z(n1931) );
  XNOR2_X2 U6726 ( .A(n4399), .B(n2762), .ZN(n4400) );
  MUX2_X2 U6727 ( .A(reg31Val_0[20]), .B(n4400), .S(net224681), .Z(n1932) );
  XNOR2_X2 U6728 ( .A(n4402), .B(n7510), .ZN(n4403) );
  MUX2_X2 U6729 ( .A(reg31Val_0[21]), .B(n4403), .S(net224681), .Z(n1933) );
  MUX2_X2 U6730 ( .A(reg31Val_0[22]), .B(n4405), .S(net224683), .Z(n1934) );
  MUX2_X2 U6731 ( .A(reg31Val_0[23]), .B(n4406), .S(net224683), .Z(n1935) );
  MUX2_X2 U6732 ( .A(reg31Val_0[24]), .B(n4408), .S(net224683), .Z(n1936) );
  XNOR2_X2 U6733 ( .A(n7506), .B(n4409), .ZN(n4410) );
  MUX2_X2 U6734 ( .A(reg31Val_0[25]), .B(n4410), .S(net224683), .Z(n1937) );
  MUX2_X2 U6735 ( .A(reg31Val_0[10]), .B(n4412), .S(net224683), .Z(n1938) );
  MUX2_X2 U6736 ( .A(reg31Val_0[11]), .B(n4414), .S(net224683), .Z(n1939) );
  INV_X4 U6737 ( .A(n4425), .ZN(n4416) );
  NAND2_X2 U6738 ( .A1(n2980), .A2(n4417), .ZN(n4421) );
  MUX2_X2 U6739 ( .A(reg31Val_0[9]), .B(n4419), .S(net224683), .Z(n1940) );
  MUX2_X2 U6740 ( .A(reg31Val_0[7]), .B(n4420), .S(net224683), .Z(n1941) );
  XNOR2_X2 U6741 ( .A(n4421), .B(n2744), .ZN(n4422) );
  MUX2_X2 U6742 ( .A(reg31Val_0[8]), .B(n4422), .S(net224683), .Z(n1942) );
  MUX2_X2 U6743 ( .A(reg31Val_0[5]), .B(n4424), .S(net224683), .Z(n1943) );
  XNOR2_X2 U6744 ( .A(n4425), .B(n2741), .ZN(n4426) );
  MUX2_X2 U6745 ( .A(reg31Val_0[6]), .B(n4426), .S(net224683), .Z(n1944) );
  MUX2_X2 U6746 ( .A(n3055), .B(n4553), .S(n3926), .Z(n1947) );
  MUX2_X2 U6747 ( .A(reg31Val_0[26]), .B(n4428), .S(net224683), .Z(n1950) );
  XNOR2_X2 U6748 ( .A(n7504), .B(n4429), .ZN(n4430) );
  MUX2_X2 U6749 ( .A(reg31Val_0[27]), .B(n4430), .S(net224683), .Z(n1952) );
  MUX2_X2 U6750 ( .A(reg31Val_0[28]), .B(n4432), .S(net224683), .Z(n1954) );
  MUX2_X2 U6751 ( .A(reg31Val_0[29]), .B(n4434), .S(net224685), .Z(n1955) );
  INV_X4 U6752 ( .A(iAddr[11]), .ZN(n4439) );
  INV_X4 U6753 ( .A(iAddr[12]), .ZN(n4438) );
  INV_X4 U6754 ( .A(n4441), .ZN(n4554) );
  MUX2_X2 U6755 ( .A(n3056), .B(n4554), .S(n3926), .Z(n1958) );
  MUX2_X2 U6756 ( .A(n3057), .B(n4555), .S(n3926), .Z(n1961) );
  INV_X4 U6757 ( .A(iAddr[7]), .ZN(n4444) );
  INV_X4 U6758 ( .A(n4446), .ZN(n4556) );
  MUX2_X2 U6759 ( .A(n3131), .B(n4556), .S(n3926), .Z(n1964) );
  XNOR2_X2 U6760 ( .A(n4448), .B(iAddr[7]), .ZN(n4557) );
  MUX2_X2 U6761 ( .A(n3058), .B(n4557), .S(n3926), .Z(n1967) );
  INV_X4 U6762 ( .A(n4450), .ZN(n4558) );
  MUX2_X2 U6763 ( .A(n3059), .B(n4558), .S(n3926), .Z(n1970) );
  MUX2_X2 U6764 ( .A(reg31Val_0[4]), .B(n4452), .S(net224685), .Z(n1971) );
  MUX2_X2 U6765 ( .A(n3060), .B(n4559), .S(n4546), .Z(n1974) );
  MUX2_X2 U6766 ( .A(reg31Val_0[3]), .B(n4457), .S(net224685), .Z(n1975) );
  MUX2_X2 U6767 ( .A(n3061), .B(n2739), .S(n3925), .Z(n1978) );
  MUX2_X2 U6768 ( .A(n3062), .B(n4560), .S(n4546), .Z(n7866) );
  NAND2_X2 U6769 ( .A1(n4524), .A2(n4459), .ZN(n4460) );
  NAND2_X2 U6770 ( .A1(n4546), .A2(n4561), .ZN(n4461) );
  NAND2_X2 U6771 ( .A1(n3926), .A2(n4563), .ZN(n4466) );
  MUX2_X2 U6772 ( .A(net223209), .B(n2969), .S(net224685), .Z(n7757) );
  MUX2_X2 U6773 ( .A(net224783), .B(link_3), .S(net224685), .Z(n1992) );
  NAND2_X2 U6774 ( .A1(iAddr[9]), .A2(n4468), .ZN(n4471) );
  MUX2_X2 U6775 ( .A(n3063), .B(n4712), .S(n4546), .Z(n1996) );
  MUX2_X2 U6776 ( .A(n3064), .B(n4710), .S(n3925), .Z(n1997) );
  MUX2_X2 U6777 ( .A(n3065), .B(n4709), .S(n3925), .Z(n1998) );
  INV_X4 U6778 ( .A(n4473), .ZN(n4474) );
  NAND2_X2 U6779 ( .A1(n4474), .A2(iAddr[13]), .ZN(n4478) );
  INV_X4 U6780 ( .A(n4478), .ZN(n4475) );
  INV_X4 U6781 ( .A(n4479), .ZN(n4476) );
  XNOR2_X2 U6782 ( .A(n4476), .B(n7915), .ZN(n4707) );
  MUX2_X2 U6783 ( .A(n3129), .B(n4706), .S(n3925), .Z(n2001) );
  MUX2_X2 U6784 ( .A(n3066), .B(n4705), .S(n3925), .Z(n2002) );
  NAND3_X4 U6785 ( .A1(n4486), .A2(iAddr[17]), .A3(iAddr[16]), .ZN(n4490) );
  INV_X4 U6786 ( .A(iAddr[18]), .ZN(n4489) );
  MUX2_X2 U6787 ( .A(n3067), .B(n4704), .S(n3925), .Z(n2003) );
  XNOR2_X2 U6788 ( .A(n7926), .B(n4491), .ZN(n4703) );
  INV_X4 U6789 ( .A(n4494), .ZN(n4702) );
  INV_X4 U6790 ( .A(iAddr[22]), .ZN(n4501) );
  INV_X4 U6791 ( .A(n4506), .ZN(n4700) );
  XNOR2_X2 U6792 ( .A(n4544), .B(n4507), .ZN(n4699) );
  NOR2_X4 U6793 ( .A1(n4533), .A2(n4514), .ZN(n4515) );
  INV_X4 U6794 ( .A(n4517), .ZN(n4696) );
  INV_X4 U6796 ( .A(n4539), .ZN(n4694) );
  XNOR2_X2 U6797 ( .A(n4545), .B(iAddr[30]), .ZN(n4693) );
  MUX2_X2 U6798 ( .A(n2843), .B(dSize[1]), .S(net224685), .Z(n2121) );
  MUX2_X2 U6799 ( .A(dSize[1]), .B(n2824), .S(n2740), .Z(n2122) );
  MUX2_X2 U6800 ( .A(n4802), .B(dSize[0]), .S(net224685), .Z(n2124) );
  MUX2_X2 U6801 ( .A(dSize[0]), .B(n2825), .S(n2740), .Z(n2125) );
  MUX2_X2 U6802 ( .A(net229988), .B(fp_3), .S(net224685), .Z(n2128) );
  MUX2_X2 U6803 ( .A(instruction[0]), .B(n2766), .S(n3929), .Z(n2139) );
  MUX2_X2 U6804 ( .A(instruction[2]), .B(n2765), .S(n3932), .Z(n2141) );
  MUX2_X2 U6805 ( .A(instruction[4]), .B(n2870), .S(n3932), .Z(n2143) );
  NAND2_X2 U6806 ( .A1(net224943), .A2(n7554), .ZN(\id_ex/N4 ) );
  NAND2_X2 U6807 ( .A1(n7579), .A2(net224915), .ZN(\ex_mem/N242 ) );
  NAND2_X2 U6808 ( .A1(n7713), .A2(n2849), .ZN(n4550) );
  NAND3_X2 U6809 ( .A1(n7628), .A2(op0_1), .A3(n2911), .ZN(n4551) );
  INV_X4 U6810 ( .A(n4667), .ZN(n4632) );
  NAND2_X2 U6811 ( .A1(n4632), .A2(n2919), .ZN(n6309) );
  NAND2_X2 U6812 ( .A1(net224967), .A2(n7555), .ZN(n7886) );
  MUX2_X2 U6813 ( .A(n2800), .B(n3012), .S(net224937), .Z(n1916) );
  MUX2_X2 U6814 ( .A(n3432), .B(n3012), .S(n3932), .Z(n1917) );
  MUX2_X2 U6815 ( .A(n2801), .B(n2721), .S(net224943), .Z(n1945) );
  MUX2_X2 U6816 ( .A(n4553), .B(n2721), .S(n3932), .Z(n1946) );
  MUX2_X2 U6817 ( .A(n2802), .B(n3013), .S(net224943), .Z(n1956) );
  MUX2_X2 U6818 ( .A(n4554), .B(n3013), .S(n3932), .Z(n1957) );
  MUX2_X2 U6819 ( .A(n3032), .B(n2826), .S(net224937), .Z(n1959) );
  MUX2_X2 U6820 ( .A(n4555), .B(n2826), .S(n3932), .Z(n1960) );
  MUX2_X2 U6821 ( .A(n2803), .B(n3014), .S(net224943), .Z(n1962) );
  MUX2_X2 U6822 ( .A(n4556), .B(n3014), .S(n3932), .Z(n1963) );
  MUX2_X2 U6823 ( .A(n2804), .B(n3015), .S(net224943), .Z(n1965) );
  MUX2_X2 U6824 ( .A(n4557), .B(n3015), .S(n3932), .Z(n1966) );
  MUX2_X2 U6825 ( .A(n2805), .B(n3016), .S(net224937), .Z(n1968) );
  MUX2_X2 U6826 ( .A(n4558), .B(n3016), .S(n3932), .Z(n1969) );
  MUX2_X2 U6827 ( .A(n2806), .B(n2722), .S(net224937), .Z(n1972) );
  MUX2_X2 U6828 ( .A(n4559), .B(n2722), .S(n3931), .Z(n1973) );
  MUX2_X2 U6829 ( .A(n2834), .B(n2705), .S(net224937), .Z(n1976) );
  MUX2_X2 U6830 ( .A(n2739), .B(n2705), .S(n3931), .Z(n1977) );
  MUX2_X2 U6831 ( .A(n3033), .B(n2827), .S(net224937), .Z(n1980) );
  MUX2_X2 U6832 ( .A(n4560), .B(n2827), .S(n3931), .Z(n1981) );
  MUX2_X2 U6833 ( .A(n2807), .B(n3017), .S(net224937), .Z(n7873) );
  INV_X4 U6834 ( .A(n4561), .ZN(n4562) );
  MUX2_X2 U6835 ( .A(iAddr[1]), .B(n3017), .S(n3931), .Z(n7862) );
  MUX2_X2 U6836 ( .A(n3034), .B(n2828), .S(net224937), .Z(n7874) );
  INV_X4 U6837 ( .A(n4563), .ZN(n4564) );
  MUX2_X2 U6838 ( .A(iAddr[0]), .B(n2828), .S(n3931), .Z(n7863) );
  NAND2_X2 U6839 ( .A1(op0_1), .A2(n4692), .ZN(n4684) );
  INV_X4 U6840 ( .A(n4684), .ZN(n4566) );
  NAND2_X2 U6841 ( .A1(n4615), .A2(n4632), .ZN(n4567) );
  MUX2_X2 U6842 ( .A(n2786), .B(n4567), .S(net224939), .Z(n4568) );
  INV_X4 U6843 ( .A(n6319), .ZN(n4604) );
  NAND2_X2 U6844 ( .A1(net224937), .A2(n2855), .ZN(n4669) );
  INV_X4 U6845 ( .A(n4669), .ZN(n7377) );
  INV_X4 U6846 ( .A(n4572), .ZN(n4573) );
  NAND2_X2 U6847 ( .A1(n7377), .A2(n4573), .ZN(n4576) );
  NAND2_X2 U6848 ( .A1(n2795), .A2(n7713), .ZN(n4671) );
  INV_X4 U6849 ( .A(n4671), .ZN(n4574) );
  NAND2_X2 U6850 ( .A1(net224947), .A2(n2847), .ZN(n4656) );
  INV_X4 U6851 ( .A(n4656), .ZN(n7378) );
  NAND4_X2 U6852 ( .A1(n4577), .A2(n4687), .A3(n4576), .A4(n4575), .ZN(n2016)
         );
  MUX2_X2 U6853 ( .A(n4579), .B(n4592), .S(n7712), .Z(n4590) );
  INV_X4 U6854 ( .A(n4672), .ZN(n4582) );
  NAND2_X2 U6855 ( .A1(n2944), .A2(n2766), .ZN(n4580) );
  MUX2_X2 U6856 ( .A(net225605), .B(n4580), .S(net224937), .Z(n4589) );
  INV_X4 U6857 ( .A(n7886), .ZN(n6303) );
  NAND3_X2 U6858 ( .A1(n2757), .A2(n4660), .A3(n4692), .ZN(n4587) );
  INV_X4 U6859 ( .A(n4663), .ZN(n4585) );
  NAND2_X2 U6860 ( .A1(n4596), .A2(n4585), .ZN(n4586) );
  NAND3_X2 U6861 ( .A1(n4590), .A2(n4589), .A3(n4588), .ZN(n2017) );
  NAND2_X2 U6862 ( .A1(n4591), .A2(n2765), .ZN(n4686) );
  NAND3_X2 U6863 ( .A1(n4593), .A2(n4686), .A3(n4592), .ZN(n4594) );
  NAND2_X2 U6864 ( .A1(n4594), .A2(n2766), .ZN(n4602) );
  NAND2_X2 U6865 ( .A1(n4597), .A2(n2757), .ZN(n4598) );
  INV_X4 U6866 ( .A(\id_ex/N4 ), .ZN(n6302) );
  NAND2_X2 U6867 ( .A1(n2944), .A2(n6302), .ZN(n4681) );
  NAND2_X2 U6868 ( .A1(n4598), .A2(n4681), .ZN(n4599) );
  NAND4_X2 U6869 ( .A1(n4602), .A2(n4601), .A3(net223781), .A4(n4600), .ZN(
        n2018) );
  MUX2_X2 U6870 ( .A(n2890), .B(busB[31]), .S(net224937), .Z(n7813) );
  MUX2_X2 U6871 ( .A(n2707), .B(busB[30]), .S(net224937), .Z(n7814) );
  MUX2_X2 U6872 ( .A(n2708), .B(busB[29]), .S(net224937), .Z(n7815) );
  MUX2_X2 U6873 ( .A(n2709), .B(busB[28]), .S(net224937), .Z(n7816) );
  MUX2_X2 U6874 ( .A(n2873), .B(busB[27]), .S(net224937), .Z(n7817) );
  MUX2_X2 U6875 ( .A(n2874), .B(busB[26]), .S(net224937), .Z(n7818) );
  MUX2_X2 U6876 ( .A(n2891), .B(busB[25]), .S(net224937), .Z(n7819) );
  MUX2_X2 U6877 ( .A(n2712), .B(busB[24]), .S(net224937), .Z(n7820) );
  MUX2_X2 U6878 ( .A(n2710), .B(busB[23]), .S(net224937), .Z(n7821) );
  MUX2_X2 U6879 ( .A(n2875), .B(busB[22]), .S(net224937), .Z(n7822) );
  MUX2_X2 U6880 ( .A(n2888), .B(busB[21]), .S(net224937), .Z(n7823) );
  MUX2_X2 U6881 ( .A(n2876), .B(busB[20]), .S(net224939), .Z(n7824) );
  MUX2_X2 U6882 ( .A(n2862), .B(busB[19]), .S(net224939), .Z(n7825) );
  MUX2_X2 U6883 ( .A(n2877), .B(busB[18]), .S(net224939), .Z(n7826) );
  MUX2_X2 U6884 ( .A(n2844), .B(busB[17]), .S(net224939), .Z(n7827) );
  MUX2_X2 U6885 ( .A(n2889), .B(busB[16]), .S(net224939), .Z(n7828) );
  MUX2_X2 U6886 ( .A(net35542), .B(busB[15]), .S(net224939), .Z(n7829) );
  MUX2_X2 U6887 ( .A(n2713), .B(busB[14]), .S(net224939), .Z(n7830) );
  MUX2_X2 U6888 ( .A(n2742), .B(busB[13]), .S(net224939), .Z(n7831) );
  MUX2_X2 U6889 ( .A(n2746), .B(busB[12]), .S(net224939), .Z(n7832) );
  MUX2_X2 U6890 ( .A(n2743), .B(busB[11]), .S(net224939), .Z(n7833) );
  MUX2_X2 U6891 ( .A(n2711), .B(busB[10]), .S(net224939), .Z(n7834) );
  MUX2_X2 U6892 ( .A(n2845), .B(busB[9]), .S(net224939), .Z(n7835) );
  MUX2_X2 U6893 ( .A(n7606), .B(busB[8]), .S(net224939), .Z(n7836) );
  MUX2_X2 U6894 ( .A(n2869), .B(busB[7]), .S(net224939), .Z(n7837) );
  MUX2_X2 U6895 ( .A(n2760), .B(busB[6]), .S(net224939), .Z(n7838) );
  MUX2_X2 U6896 ( .A(n2745), .B(busB[5]), .S(net224939), .Z(n7839) );
  MUX2_X2 U6897 ( .A(n2747), .B(busB[4]), .S(net224939), .Z(n7840) );
  MUX2_X2 U6898 ( .A(n7607), .B(busB[3]), .S(net224939), .Z(n7841) );
  MUX2_X2 U6899 ( .A(n2748), .B(busB[2]), .S(net224939), .Z(n7842) );
  MUX2_X2 U6900 ( .A(n2749), .B(busB[1]), .S(net224939), .Z(n7843) );
  MUX2_X2 U6901 ( .A(n2878), .B(busB[0]), .S(net224939), .Z(n7844) );
  MUX2_X2 U6902 ( .A(n2714), .B(busA[31]), .S(net224937), .Z(n7781) );
  MUX2_X2 U6903 ( .A(n2864), .B(busA[30]), .S(net224937), .Z(n7782) );
  MUX2_X2 U6904 ( .A(n2750), .B(busA[29]), .S(net224937), .Z(n7783) );
  MUX2_X2 U6905 ( .A(n2860), .B(busA[28]), .S(net224937), .Z(n7784) );
  MUX2_X2 U6906 ( .A(n2872), .B(busA[27]), .S(net224937), .Z(n7785) );
  MUX2_X2 U6907 ( .A(n2866), .B(busA[26]), .S(net224937), .Z(n7786) );
  MUX2_X2 U6908 ( .A(n2751), .B(busA[25]), .S(net224937), .Z(n7787) );
  MUX2_X2 U6909 ( .A(n2879), .B(busA[24]), .S(net224937), .Z(n7788) );
  MUX2_X2 U6910 ( .A(n2715), .B(busA[23]), .S(net224937), .Z(n7789) );
  MUX2_X2 U6911 ( .A(n2716), .B(busA[22]), .S(net224937), .Z(n7790) );
  MUX2_X2 U6912 ( .A(n7603), .B(busA[21]), .S(net224937), .Z(n7791) );
  MUX2_X2 U6913 ( .A(n2717), .B(busA[20]), .S(net224937), .Z(n7792) );
  MUX2_X2 U6914 ( .A(n2718), .B(busA[19]), .S(net224937), .Z(n7793) );
  MUX2_X2 U6915 ( .A(n2752), .B(busA[18]), .S(net224937), .Z(n7794) );
  MUX2_X2 U6916 ( .A(n2880), .B(busA[17]), .S(net224937), .Z(n7795) );
  MUX2_X2 U6917 ( .A(n2892), .B(busA[16]), .S(net224937), .Z(n7796) );
  MUX2_X2 U6918 ( .A(n2881), .B(busA[15]), .S(net224937), .Z(n7797) );
  MUX2_X2 U6919 ( .A(n2861), .B(busA[14]), .S(net224937), .Z(n7798) );
  MUX2_X2 U6920 ( .A(n2893), .B(busA[13]), .S(net224937), .Z(n7799) );
  MUX2_X2 U6921 ( .A(n3744), .B(busA[12]), .S(net224937), .Z(n7800) );
  MUX2_X2 U6922 ( .A(n2895), .B(busA[11]), .S(net224937), .Z(n7801) );
  MUX2_X2 U6923 ( .A(n2894), .B(busA[10]), .S(net224943), .Z(n7802) );
  MUX2_X2 U6924 ( .A(n2882), .B(busA[9]), .S(net224943), .Z(n7803) );
  MUX2_X2 U6925 ( .A(n2865), .B(busA[8]), .S(net224943), .Z(n7804) );
  MUX2_X2 U6926 ( .A(n7605), .B(busA[7]), .S(net224943), .Z(n7805) );
  MUX2_X2 U6927 ( .A(n2753), .B(busA[6]), .S(net224943), .Z(n7806) );
  MUX2_X2 U6928 ( .A(n2883), .B(busA[5]), .S(net224943), .Z(n7807) );
  MUX2_X2 U6929 ( .A(n2884), .B(busA[4]), .S(net224943), .Z(n7808) );
  MUX2_X2 U6930 ( .A(n2885), .B(busA[3]), .S(net224943), .Z(n7809) );
  MUX2_X2 U6931 ( .A(n2886), .B(busA[2]), .S(net224943), .Z(n7810) );
  MUX2_X2 U6932 ( .A(n2754), .B(busA[1]), .S(net224943), .Z(n7811) );
  MUX2_X2 U6933 ( .A(n2755), .B(busA[0]), .S(net224943), .Z(n7812) );
  NAND2_X2 U6934 ( .A1(n4604), .A2(n4603), .ZN(n4690) );
  NAND2_X2 U6935 ( .A1(n2724), .A2(n2849), .ZN(n4605) );
  NAND2_X2 U6936 ( .A1(net224943), .A2(n2939), .ZN(n4614) );
  NAND2_X2 U6937 ( .A1(rd_2[4]), .A2(net224957), .ZN(n4606) );
  OAI221_X2 U6938 ( .B1(n4607), .B2(n4691), .C1(n4690), .C2(n4614), .A(n4606), 
        .ZN(n2083) );
  NAND2_X2 U6939 ( .A1(net224937), .A2(n2955), .ZN(n6330) );
  NAND2_X2 U6940 ( .A1(rd_2[3]), .A2(net224957), .ZN(n4608) );
  OAI221_X2 U6941 ( .B1(n4609), .B2(n4691), .C1(n4690), .C2(n6330), .A(n4608), 
        .ZN(n2084) );
  NAND2_X2 U6942 ( .A1(net224937), .A2(n2956), .ZN(n6329) );
  NAND2_X2 U6943 ( .A1(rd_2[2]), .A2(net224957), .ZN(n4610) );
  OAI221_X2 U6944 ( .B1(n4611), .B2(n4691), .C1(n4690), .C2(n6329), .A(n4610), 
        .ZN(n2086) );
  NAND2_X2 U6945 ( .A1(net224937), .A2(n2957), .ZN(n6328) );
  NAND2_X2 U6946 ( .A1(rd_2[1]), .A2(net224957), .ZN(n4612) );
  OAI221_X2 U6947 ( .B1(n4613), .B2(n4691), .C1(n4690), .C2(n6328), .A(n4612), 
        .ZN(n2088) );
  INV_X4 U6948 ( .A(n4614), .ZN(n7376) );
  NAND2_X2 U6949 ( .A1(n7376), .A2(n4657), .ZN(n4655) );
  NAND2_X2 U6950 ( .A1(op0_1), .A2(n7708), .ZN(n4616) );
  INV_X4 U6951 ( .A(n4617), .ZN(n4670) );
  NOR3_X4 U6952 ( .A1(n4655), .A2(n4619), .A3(n4618), .ZN(n4633) );
  NAND2_X2 U6953 ( .A1(n2702), .A2(n2939), .ZN(n4620) );
  NAND2_X2 U6954 ( .A1(n4621), .A2(n4620), .ZN(n2089) );
  NAND2_X2 U6955 ( .A1(n2702), .A2(n2955), .ZN(n4622) );
  NAND2_X2 U6956 ( .A1(n4623), .A2(n4622), .ZN(n2090) );
  NAND2_X2 U6957 ( .A1(n2702), .A2(n2956), .ZN(n4624) );
  NAND2_X2 U6958 ( .A1(n4625), .A2(n4624), .ZN(n2091) );
  NAND2_X2 U6959 ( .A1(n2702), .A2(n2957), .ZN(n4626) );
  NAND2_X2 U6960 ( .A1(n4627), .A2(n4626), .ZN(n2092) );
  NAND2_X2 U6961 ( .A1(n2702), .A2(n2958), .ZN(n4628) );
  NAND2_X2 U6962 ( .A1(n4629), .A2(n4628), .ZN(n2093) );
  NAND2_X2 U6963 ( .A1(n2702), .A2(n2938), .ZN(n4630) );
  NAND2_X2 U6964 ( .A1(n4631), .A2(n4630), .ZN(n2094) );
  NAND2_X2 U6965 ( .A1(n7372), .A2(n4667), .ZN(n4635) );
  AOI22_X2 U6966 ( .A1(net224957), .A2(n2930), .B1(n2702), .B2(n2936), .ZN(
        n4634) );
  NAND3_X2 U6967 ( .A1(n4635), .A2(n4652), .A3(n4634), .ZN(n2095) );
  NAND2_X2 U6968 ( .A1(n2926), .A2(n4667), .ZN(n4637) );
  AOI22_X2 U6969 ( .A1(net224957), .A2(n2773), .B1(n2702), .B2(n2935), .ZN(
        n4636) );
  NAND3_X2 U6970 ( .A1(n4637), .A2(n4652), .A3(n4636), .ZN(n2096) );
  NAND2_X2 U6971 ( .A1(n7371), .A2(n4667), .ZN(n4639) );
  AOI22_X2 U6972 ( .A1(net224957), .A2(n2763), .B1(n2702), .B2(n2934), .ZN(
        n4638) );
  NAND3_X2 U6973 ( .A1(n4639), .A2(n4652), .A3(n4638), .ZN(n2097) );
  NAND2_X2 U6974 ( .A1(n7370), .A2(n4667), .ZN(n4641) );
  AOI22_X2 U6975 ( .A1(net224957), .A2(n2764), .B1(n2702), .B2(n2933), .ZN(
        n4640) );
  NAND3_X2 U6976 ( .A1(n4641), .A2(n4652), .A3(n4640), .ZN(n2098) );
  NAND2_X2 U6977 ( .A1(n7378), .A2(n4658), .ZN(n4643) );
  AOI22_X2 U6978 ( .A1(n7369), .A2(n4667), .B1(net224957), .B2(n2906), .ZN(
        n4642) );
  NAND3_X2 U6979 ( .A1(n4643), .A2(n4652), .A3(n4642), .ZN(n2099) );
  NAND2_X2 U6980 ( .A1(n3074), .A2(n4667), .ZN(n4645) );
  AOI22_X2 U6981 ( .A1(net224957), .A2(n2901), .B1(n2702), .B2(n2870), .ZN(
        n4644) );
  NAND3_X2 U6982 ( .A1(n4645), .A2(n4652), .A3(n4644), .ZN(n2100) );
  NAND2_X2 U6983 ( .A1(n3073), .A2(n4667), .ZN(n4646) );
  NAND3_X2 U6984 ( .A1(n4646), .A2(n4652), .A3(net223721), .ZN(n2101) );
  NAND2_X2 U6985 ( .A1(n3072), .A2(n4667), .ZN(n4648) );
  AOI22_X2 U6986 ( .A1(net224957), .A2(n2931), .B1(n2702), .B2(n2765), .ZN(
        n4647) );
  NAND3_X2 U6987 ( .A1(n4648), .A2(n4652), .A3(n4647), .ZN(n2102) );
  NAND2_X2 U6988 ( .A1(n3071), .A2(n4667), .ZN(n4650) );
  AOI22_X2 U6989 ( .A1(net224957), .A2(n2917), .B1(n2702), .B2(n2720), .ZN(
        n4649) );
  NAND3_X2 U6990 ( .A1(n4650), .A2(n4652), .A3(n4649), .ZN(n2103) );
  NAND2_X2 U6991 ( .A1(n2702), .A2(n2766), .ZN(n4653) );
  AOI22_X2 U6992 ( .A1(n2835), .A2(n4667), .B1(net224957), .B2(n2932), .ZN(
        n4651) );
  NAND3_X2 U6993 ( .A1(n4653), .A2(n4652), .A3(n4651), .ZN(n2104) );
  NAND2_X2 U6994 ( .A1(net224957), .A2(n2859), .ZN(n4654) );
  NAND2_X2 U6995 ( .A1(n4655), .A2(n4654), .ZN(n2105) );
  OAI22_X2 U6996 ( .A1(n7726), .A2(net224943), .B1(n4658), .B2(n6330), .ZN(
        n2106) );
  OAI22_X2 U6997 ( .A1(n7722), .A2(net224943), .B1(n4658), .B2(n6329), .ZN(
        n2107) );
  OAI22_X2 U6998 ( .A1(n7725), .A2(net224943), .B1(n4658), .B2(n6328), .ZN(
        n2108) );
  NAND2_X2 U6999 ( .A1(net224937), .A2(n2958), .ZN(n6327) );
  OAI22_X2 U7000 ( .A1(n7724), .A2(net224943), .B1(n4658), .B2(n6327), .ZN(
        n2109) );
  NAND2_X2 U7001 ( .A1(net224937), .A2(n2938), .ZN(n6326) );
  OAI22_X2 U7002 ( .A1(net33193), .A2(net224943), .B1(n4658), .B2(n6326), .ZN(
        n7880) );
  NAND2_X2 U7003 ( .A1(net224937), .A2(n2936), .ZN(n6325) );
  OAI22_X2 U7004 ( .A1(n7743), .A2(net224943), .B1(n4658), .B2(n6325), .ZN(
        n7879) );
  NAND2_X2 U7005 ( .A1(net224937), .A2(n2935), .ZN(n6324) );
  OAI22_X2 U7006 ( .A1(n7744), .A2(net224943), .B1(n4658), .B2(n6324), .ZN(
        n7878) );
  NAND2_X2 U7007 ( .A1(net224937), .A2(n2934), .ZN(n6323) );
  OAI22_X2 U7008 ( .A1(n7745), .A2(net224943), .B1(n4658), .B2(n6323), .ZN(
        n7877) );
  NAND2_X2 U7009 ( .A1(net224937), .A2(n2933), .ZN(n6322) );
  OAI22_X2 U7010 ( .A1(n7746), .A2(net224943), .B1(n4658), .B2(n6322), .ZN(
        n7876) );
  NAND2_X2 U7011 ( .A1(net224937), .A2(n4657), .ZN(n4659) );
  OAI22_X2 U7012 ( .A1(n7721), .A2(net224943), .B1(n7556), .B2(n4659), .ZN(
        n2116) );
  NAND2_X2 U7013 ( .A1(net224937), .A2(n2761), .ZN(n6300) );
  OAI22_X2 U7014 ( .A1(n7748), .A2(net224943), .B1(n4658), .B2(n6300), .ZN(
        n7887) );
  OAI22_X2 U7015 ( .A1(n7720), .A2(net224943), .B1(n7555), .B2(n4659), .ZN(
        n2118) );
  NAND2_X2 U7016 ( .A1(net224939), .A2(n2720), .ZN(n6301) );
  OAI22_X2 U7017 ( .A1(n7749), .A2(net224943), .B1(n4658), .B2(n6301), .ZN(
        n7885) );
  OAI22_X2 U7018 ( .A1(n7733), .A2(net224943), .B1(n7554), .B2(n4659), .ZN(
        n2120) );
  INV_X4 U7019 ( .A(n4660), .ZN(n4675) );
  NAND2_X2 U7020 ( .A1(n2795), .A2(n2724), .ZN(n6332) );
  NAND2_X2 U7021 ( .A1(net224957), .A2(n2824), .ZN(n4661) );
  NAND2_X2 U7022 ( .A1(net224957), .A2(n2825), .ZN(n4662) );
  OAI221_X2 U7023 ( .B1(n4663), .B2(n6332), .C1(n2846), .C2(n4671), .A(n4662), 
        .ZN(n2126) );
  NAND2_X2 U7024 ( .A1(net224937), .A2(op0_1), .ZN(n6331) );
  NAND2_X2 U7025 ( .A1(op0_2), .A2(net224957), .ZN(n4664) );
  NAND2_X2 U7026 ( .A1(n6331), .A2(n4664), .ZN(n2127) );
  OAI22_X2 U7027 ( .A1(n7718), .A2(net224943), .B1(n7556), .B2(n4665), .ZN(
        n2129) );
  MUX2_X2 U7028 ( .A(n2867), .B(n6311), .S(net224943), .Z(n2130) );
  MUX2_X2 U7029 ( .A(n2971), .B(n4667), .S(net224943), .Z(n2131) );
  OAI22_X2 U7030 ( .A1(n7644), .A2(net224943), .B1(n4670), .B2(n4669), .ZN(
        n2133) );
  NAND2_X2 U7031 ( .A1(n4676), .A2(n4675), .ZN(n4677) );
  MUX2_X2 U7032 ( .A(net224747), .B(n3095), .S(net224943), .Z(n2136) );
  NAND2_X2 U7033 ( .A1(net224957), .A2(n2704), .ZN(n4685) );
  NAND4_X2 U7034 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n2137)
         );
  NAND2_X2 U7035 ( .A1(rd_2[0]), .A2(net224957), .ZN(n4689) );
  OAI221_X2 U7036 ( .B1(n6291), .B2(n4691), .C1(n4690), .C2(n6327), .A(n4689), 
        .ZN(n2138) );
  MUX2_X2 U7037 ( .A(instruction[1]), .B(n2720), .S(n3931), .Z(n2140) );
  MUX2_X2 U7038 ( .A(instruction[3]), .B(n2761), .S(n3931), .Z(n2142) );
  MUX2_X2 U7039 ( .A(instruction[5]), .B(n2847), .S(n3931), .Z(n2144) );
  MUX2_X2 U7040 ( .A(instruction[6]), .B(n2933), .S(n3931), .Z(n2145) );
  MUX2_X2 U7041 ( .A(instruction[7]), .B(n2934), .S(n3931), .Z(n2146) );
  MUX2_X2 U7042 ( .A(instruction[8]), .B(n2935), .S(n3931), .Z(n2147) );
  MUX2_X2 U7043 ( .A(instruction[9]), .B(n2936), .S(n3931), .Z(n2148) );
  MUX2_X2 U7044 ( .A(instruction[10]), .B(n2938), .S(n3931), .Z(n2149) );
  MUX2_X2 U7045 ( .A(instruction[11]), .B(n2958), .S(n3931), .Z(n2150) );
  MUX2_X2 U7046 ( .A(instruction[12]), .B(n2957), .S(n3930), .Z(n2151) );
  MUX2_X2 U7047 ( .A(instruction[13]), .B(n2956), .S(n3930), .Z(n2152) );
  MUX2_X2 U7048 ( .A(instruction[14]), .B(n2955), .S(n3930), .Z(n2153) );
  MUX2_X2 U7049 ( .A(instruction[15]), .B(n2939), .S(n3930), .Z(n2154) );
  MUX2_X2 U7050 ( .A(instruction[16]), .B(n2963), .S(n3930), .Z(n2155) );
  MUX2_X2 U7051 ( .A(instruction[17]), .B(n2952), .S(n3930), .Z(n2156) );
  MUX2_X2 U7052 ( .A(instruction[18]), .B(n2953), .S(n3930), .Z(n2157) );
  MUX2_X2 U7053 ( .A(instruction[19]), .B(n2954), .S(n3930), .Z(n2158) );
  MUX2_X2 U7054 ( .A(instruction[20]), .B(n2968), .S(n3930), .Z(n2159) );
  MUX2_X2 U7055 ( .A(instruction[21]), .B(rs1[0]), .S(n3930), .Z(n2160) );
  MUX2_X2 U7056 ( .A(instruction[22]), .B(rs1[1]), .S(n3930), .Z(n2161) );
  MUX2_X2 U7057 ( .A(instruction[23]), .B(rs1[2]), .S(n3930), .Z(n2162) );
  MUX2_X2 U7058 ( .A(instruction[24]), .B(rs1[3]), .S(n3930), .Z(n2163) );
  MUX2_X2 U7059 ( .A(instruction[25]), .B(rs1[4]), .S(n3929), .Z(n2164) );
  MUX2_X2 U7060 ( .A(instruction[26]), .B(op0_1), .S(n3929), .Z(n2165) );
  MUX2_X2 U7061 ( .A(instruction[27]), .B(n4692), .S(n3929), .Z(n2166) );
  MUX2_X2 U7062 ( .A(instruction[28]), .B(n2855), .S(n3929), .Z(n2167) );
  MUX2_X2 U7063 ( .A(instruction[29]), .B(n2868), .S(n3929), .Z(n2168) );
  MUX2_X2 U7064 ( .A(instruction[30]), .B(n2858), .S(n3929), .Z(n2169) );
  MUX2_X2 U7065 ( .A(instruction[31]), .B(n2849), .S(n3929), .Z(n2170) );
  MUX2_X2 U7066 ( .A(n2808), .B(n2987), .S(net224943), .Z(n2175) );
  MUX2_X2 U7067 ( .A(n2809), .B(n3018), .S(net224943), .Z(n2177) );
  MUX2_X2 U7068 ( .A(n2626), .B(n3018), .S(n3929), .Z(n2178) );
  MUX2_X2 U7069 ( .A(n2810), .B(n3019), .S(net224943), .Z(n2179) );
  MUX2_X2 U7070 ( .A(n4694), .B(n3019), .S(n3929), .Z(n2180) );
  MUX2_X2 U7071 ( .A(n2811), .B(n3020), .S(net224943), .Z(n2181) );
  MUX2_X2 U7072 ( .A(n4695), .B(n3020), .S(n3929), .Z(n2182) );
  MUX2_X2 U7073 ( .A(n2812), .B(n3021), .S(net224943), .Z(n2183) );
  MUX2_X2 U7074 ( .A(n4696), .B(n3021), .S(n3929), .Z(n2184) );
  MUX2_X2 U7075 ( .A(n2813), .B(n3022), .S(net224943), .Z(n2185) );
  MUX2_X2 U7076 ( .A(n2686), .B(n3022), .S(n3929), .Z(n2186) );
  MUX2_X2 U7077 ( .A(n2814), .B(n3023), .S(net224933), .Z(n2187) );
  MUX2_X2 U7078 ( .A(n4698), .B(n3023), .S(n3929), .Z(n2188) );
  MUX2_X2 U7079 ( .A(n3035), .B(n2829), .S(net224933), .Z(n2189) );
  MUX2_X2 U7080 ( .A(n4699), .B(n2829), .S(n3929), .Z(n2190) );
  MUX2_X2 U7081 ( .A(n2815), .B(n3024), .S(net224943), .Z(n2191) );
  MUX2_X2 U7082 ( .A(n4700), .B(n3024), .S(n3929), .Z(n2192) );
  MUX2_X2 U7083 ( .A(n2816), .B(n3025), .S(net224933), .Z(n2193) );
  MUX2_X2 U7084 ( .A(n2685), .B(n3025), .S(n3931), .Z(n2194) );
  MUX2_X2 U7085 ( .A(n2817), .B(n3026), .S(net224933), .Z(n2195) );
  MUX2_X2 U7086 ( .A(n4702), .B(n3026), .S(n3930), .Z(n2196) );
  MUX2_X2 U7087 ( .A(n2818), .B(n3027), .S(net224933), .Z(n2197) );
  MUX2_X2 U7088 ( .A(n4703), .B(n3027), .S(n3932), .Z(n2198) );
  MUX2_X2 U7089 ( .A(n3036), .B(n2830), .S(net224933), .Z(n2199) );
  MUX2_X2 U7090 ( .A(n4704), .B(n2830), .S(n3931), .Z(n2200) );
  MUX2_X2 U7091 ( .A(n3037), .B(n2831), .S(net224933), .Z(n2201) );
  MUX2_X2 U7092 ( .A(n4705), .B(n2831), .S(n3930), .Z(n2202) );
  MUX2_X2 U7093 ( .A(n2819), .B(n3028), .S(net224933), .Z(n2203) );
  MUX2_X2 U7094 ( .A(n4706), .B(n3028), .S(n3932), .Z(n2204) );
  MUX2_X2 U7095 ( .A(n3038), .B(n2832), .S(net224933), .Z(n2205) );
  MUX2_X2 U7096 ( .A(n4707), .B(n2832), .S(n3931), .Z(n2206) );
  MUX2_X2 U7097 ( .A(n2820), .B(n3029), .S(net224933), .Z(n2207) );
  MUX2_X2 U7098 ( .A(n4708), .B(n3029), .S(n3930), .Z(n2208) );
  MUX2_X2 U7099 ( .A(n2821), .B(n3030), .S(net224933), .Z(n2209) );
  MUX2_X2 U7100 ( .A(n4709), .B(n3030), .S(n3932), .Z(n2210) );
  MUX2_X2 U7101 ( .A(n3039), .B(n2833), .S(net224933), .Z(n2211) );
  MUX2_X2 U7102 ( .A(n4710), .B(n2833), .S(n3931), .Z(n2212) );
  MUX2_X2 U7103 ( .A(n2822), .B(n3031), .S(net224933), .Z(n2213) );
  MUX2_X2 U7104 ( .A(n4712), .B(n3031), .S(n3930), .Z(n2214) );
  NAND4_X2 U7105 ( .A1(n2697), .A2(n3175), .A3(\wb/dsize_reg/z2 [7]), .A4(
        net225251), .ZN(n5309) );
  NAND4_X2 U7106 ( .A1(n3118), .A2(net228697), .A3(net224787), .A4(net225251), 
        .ZN(n5088) );
  NAND4_X2 U7107 ( .A1(n3813), .A2(net225251), .A3(\wb/dsize_reg/z2 [31]), 
        .A4(n7921), .ZN(n5308) );
  INV_X4 U7108 ( .A(n7527), .ZN(n4719) );
  AOI211_X4 U7109 ( .C1(n4731), .C2(net225216), .A(n4729), .B(n4730), .ZN(
        n5145) );
  NAND3_X2 U7110 ( .A1(n4734), .A2(net224783), .A3(net224993), .ZN(n4739) );
  NOR3_X4 U7112 ( .A1(n3905), .A2(n3899), .A3(n7574), .ZN(n4743) );
  OAI21_X4 U7114 ( .B1(n4750), .B2(net223242), .A(n4749), .ZN(n5149) );
  OAI21_X4 U7115 ( .B1(n4753), .B2(net223242), .A(n4752), .ZN(n5150) );
  NAND3_X4 U7116 ( .A1(\wb/dsize_reg/z2 [31]), .A2(n4881), .A3(n3412), .ZN(
        n4762) );
  NOR2_X4 U7117 ( .A1(n4762), .A2(n3291), .ZN(n4764) );
  NOR3_X4 U7118 ( .A1(n4772), .A2(net228233), .A3(net229307), .ZN(n5244) );
  INV_X4 U7119 ( .A(n5003), .ZN(n4997) );
  INV_X4 U7120 ( .A(n5358), .ZN(n4776) );
  INV_X4 U7121 ( .A(n3864), .ZN(n4781) );
  NAND2_X2 U7122 ( .A1(reg31Val_0[2]), .A2(net224783), .ZN(n4978) );
  NOR2_X4 U7123 ( .A1(n7568), .A2(n3290), .ZN(n4782) );
  OAI21_X4 U7124 ( .B1(net224999), .B2(n4978), .A(n4783), .ZN(n5624) );
  INV_X4 U7125 ( .A(n5616), .ZN(n5626) );
  NAND2_X2 U7126 ( .A1(n4786), .A2(n5626), .ZN(regWrData[2]) );
  INV_X4 U7127 ( .A(regWrData[2]), .ZN(n5284) );
  INV_X4 U7128 ( .A(n4787), .ZN(n4788) );
  NAND2_X2 U7130 ( .A1(n4789), .A2(net225214), .ZN(n5586) );
  INV_X4 U7131 ( .A(n4792), .ZN(regWrData[1]) );
  INV_X4 U7132 ( .A(n4973), .ZN(n4794) );
  INV_X4 U7133 ( .A(n4974), .ZN(n4793) );
  OAI22_X2 U7134 ( .A1(n2784), .A2(n3855), .B1(n5009), .B2(n3291), .ZN(n5577)
         );
  NAND2_X2 U7135 ( .A1(n3771), .A2(net224995), .ZN(n5575) );
  OAI22_X2 U7136 ( .A1(n7566), .A2(net225015), .B1(n3935), .B2(n3087), .ZN(
        n4796) );
  INV_X4 U7137 ( .A(n4796), .ZN(n5580) );
  NAND2_X2 U7138 ( .A1(reg31Val_0[6]), .A2(net224783), .ZN(n4800) );
  INV_X4 U7139 ( .A(n4800), .ZN(n5095) );
  NAND2_X2 U7140 ( .A1(n5095), .A2(net224995), .ZN(n5436) );
  INV_X4 U7141 ( .A(n2581), .ZN(n4801) );
  NOR2_X4 U7142 ( .A1(net224783), .A2(n2732), .ZN(n4804) );
  NAND4_X2 U7143 ( .A1(n3813), .A2(net230143), .A3(\wb/dsize_reg/z2 [30]), 
        .A4(net224787), .ZN(n5441) );
  NAND2_X2 U7145 ( .A1(n4812), .A2(memAddr[11]), .ZN(n5035) );
  NOR2_X4 U7146 ( .A1(n3903), .A2(n2947), .ZN(n4813) );
  NAND2_X2 U7147 ( .A1(reg31Val_0[11]), .A2(net224783), .ZN(n4958) );
  INV_X4 U7148 ( .A(n4958), .ZN(n4815) );
  INV_X4 U7149 ( .A(n4818), .ZN(\ex_mem/N110 ) );
  OAI21_X4 U7150 ( .B1(net223242), .B2(n4826), .A(n4825), .ZN(n5341) );
  NAND2_X2 U7152 ( .A1(n4830), .A2(n3904), .ZN(n4831) );
  INV_X4 U7153 ( .A(n4831), .ZN(n5118) );
  NAND2_X2 U7155 ( .A1(net223245), .A2(n2746), .ZN(n5022) );
  NAND2_X2 U7156 ( .A1(reg31Val_0[12]), .A2(net224783), .ZN(n5271) );
  NOR2_X4 U7159 ( .A1(n3899), .A2(n2948), .ZN(n4836) );
  NAND3_X2 U7160 ( .A1(n4836), .A2(n4856), .A3(net225047), .ZN(n4837) );
  INV_X4 U7161 ( .A(n4840), .ZN(\ex_mem/N111 ) );
  NAND2_X2 U7162 ( .A1(\wb/dsize_reg/z2 [13]), .A2(n3898), .ZN(n5421) );
  NAND2_X2 U7163 ( .A1(reg31Val_0[13]), .A2(net225237), .ZN(n5417) );
  INV_X4 U7164 ( .A(n4841), .ZN(n5112) );
  NAND2_X2 U7165 ( .A1(n3086), .A2(n3898), .ZN(n5418) );
  NOR2_X4 U7166 ( .A1(n5379), .A2(n5377), .ZN(n5131) );
  INV_X4 U7167 ( .A(n4849), .ZN(n4950) );
  INV_X4 U7168 ( .A(n5382), .ZN(n4853) );
  NAND2_X2 U7169 ( .A1(\wb/dsize_reg/z2 [10]), .A2(n3898), .ZN(n5383) );
  INV_X4 U7170 ( .A(n5378), .ZN(n4852) );
  NAND2_X2 U7171 ( .A1(reg31Val_0[30]), .A2(net224783), .ZN(n4860) );
  INV_X4 U7172 ( .A(n4860), .ZN(n5667) );
  NAND2_X2 U7173 ( .A1(n4861), .A2(net225047), .ZN(n4862) );
  INV_X4 U7174 ( .A(regWrData[19]), .ZN(n4870) );
  OAI21_X4 U7176 ( .B1(n4870), .B2(n3940), .A(n4869), .ZN(net221491) );
  NAND3_X4 U7177 ( .A1(reg31Val_0[5]), .A2(net224781), .A3(net225045), .ZN(
        n5527) );
  NAND3_X4 U7178 ( .A1(\wb/dsize_reg/z2 [5]), .A2(n4856), .A3(net225045), .ZN(
        n5523) );
  NAND3_X4 U7179 ( .A1(n5527), .A2(n5058), .A3(n5523), .ZN(n5547) );
  INV_X4 U7180 ( .A(n5547), .ZN(n4872) );
  INV_X4 U7181 ( .A(n5548), .ZN(n4871) );
  NAND2_X2 U7182 ( .A1(n4872), .A2(n4871), .ZN(regWrData[5]) );
  INV_X4 U7183 ( .A(regWrData[5]), .ZN(n5691) );
  INV_X4 U7184 ( .A(n4873), .ZN(n4874) );
  INV_X4 U7185 ( .A(n5474), .ZN(n5043) );
  INV_X4 U7186 ( .A(n4966), .ZN(n4895) );
  NOR2_X4 U7187 ( .A1(n3933), .A2(n4896), .ZN(n5770) );
  OAI22_X2 U7188 ( .A1(n7412), .A2(n2623), .B1(n7683), .B2(net225243), .ZN(
        n5767) );
  NAND2_X2 U7189 ( .A1(n3906), .A2(reg31Val_0[18]), .ZN(n4898) );
  NAND3_X2 U7190 ( .A1(n4900), .A2(net224783), .A3(net224993), .ZN(n4906) );
  INV_X4 U7191 ( .A(n3875), .ZN(n4907) );
  NAND3_X2 U7192 ( .A1(n4908), .A2(net224783), .A3(net225251), .ZN(n4914) );
  NAND2_X2 U7193 ( .A1(n4909), .A2(net225251), .ZN(n4913) );
  AOI21_X4 U7194 ( .B1(n4911), .B2(net225251), .A(n4910), .ZN(n4912) );
  NOR3_X4 U7195 ( .A1(n3905), .A2(n3899), .A3(n7551), .ZN(n4926) );
  OAI21_X4 U7196 ( .B1(n4933), .B2(net223242), .A(n4932), .ZN(n6165) );
  OAI21_X4 U7197 ( .B1(n3291), .B2(n4937), .A(n4936), .ZN(n5652) );
  INV_X4 U7198 ( .A(n5652), .ZN(n4938) );
  NAND2_X2 U7199 ( .A1(n4938), .A2(n5650), .ZN(regWrData[17]) );
  INV_X4 U7200 ( .A(regWrData[17]), .ZN(n4939) );
  OAI21_X4 U7201 ( .B1(n4939), .B2(n3941), .A(n5655), .ZN(n6349) );
  INV_X4 U7203 ( .A(n4940), .ZN(n4945) );
  NAND2_X2 U7204 ( .A1(reg31Val_0[14]), .A2(n3937), .ZN(n4947) );
  OAI21_X4 U7205 ( .B1(n3933), .B2(n2964), .A(n4951), .ZN(n5798) );
  INV_X4 U7206 ( .A(n5499), .ZN(n4959) );
  INV_X4 U7207 ( .A(n5561), .ZN(n4961) );
  NAND2_X2 U7208 ( .A1(net225011), .A2(n2992), .ZN(n5558) );
  NAND3_X4 U7209 ( .A1(n4961), .A2(n5560), .A3(n5558), .ZN(regWrData[16]) );
  INV_X4 U7210 ( .A(n6053), .ZN(n4962) );
  NAND2_X2 U7211 ( .A1(net225011), .A2(n3077), .ZN(n6051) );
  INV_X4 U7212 ( .A(n4964), .ZN(n5404) );
  OAI22_X2 U7213 ( .A1(n2700), .A2(n2837), .B1(n7559), .B2(net225015), .ZN(
        n4965) );
  INV_X4 U7214 ( .A(n4965), .ZN(n5403) );
  MUX2_X2 U7216 ( .A(net224843), .B(n7151), .S(n5779), .Z(n4972) );
  NAND4_X2 U7217 ( .A1(n4973), .A2(n4974), .A3(n5588), .A4(n5585), .ZN(n5594)
         );
  NAND2_X2 U7218 ( .A1(net224737), .A2(n4974), .ZN(n4976) );
  NAND2_X2 U7219 ( .A1(n7749), .A2(net224747), .ZN(n4975) );
  OAI21_X4 U7220 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(n5593) );
  OAI21_X4 U7221 ( .B1(n5594), .B2(n5596), .A(n5595), .ZN(n6965) );
  INV_X4 U7222 ( .A(n6965), .ZN(n7230) );
  NAND2_X2 U7223 ( .A1(\wb/dsize_reg/z2 [2]), .A2(net224751), .ZN(n4982) );
  NOR2_X4 U7224 ( .A1(net225051), .A2(n2650), .ZN(n4983) );
  NAND3_X4 U7225 ( .A1(n4984), .A2(n4985), .A3(n2943), .ZN(n5568) );
  INV_X4 U7226 ( .A(n4993), .ZN(n4994) );
  NOR3_X4 U7228 ( .A1(n4999), .A2(n4998), .A3(n4997), .ZN(n5000) );
  NAND2_X2 U7229 ( .A1(n7721), .A2(net224747), .ZN(n5544) );
  NAND3_X4 U7230 ( .A1(n3611), .A2(n5544), .A3(n5545), .ZN(n6842) );
  NAND3_X2 U7231 ( .A1(n5010), .A2(n5015), .A3(net224993), .ZN(n5215) );
  NAND3_X2 U7232 ( .A1(n5219), .A2(n5215), .A3(n5216), .ZN(n5018) );
  NAND3_X2 U7233 ( .A1(n5218), .A2(n5220), .A3(net224737), .ZN(n5017) );
  NAND2_X2 U7234 ( .A1(n7748), .A2(net224747), .ZN(n5016) );
  OAI21_X4 U7235 ( .B1(n5018), .B2(n5017), .A(n5016), .ZN(n5631) );
  NAND2_X2 U7236 ( .A1(n3916), .A2(n3523), .ZN(n6461) );
  NAND3_X4 U7237 ( .A1(n5019), .A2(net224731), .A3(n5773), .ZN(n5020) );
  NAND2_X2 U7238 ( .A1(n7740), .A2(net224747), .ZN(n5771) );
  INV_X4 U7239 ( .A(n5022), .ZN(n5023) );
  INV_X4 U7241 ( .A(n3280), .ZN(n5037) );
  NAND2_X2 U7242 ( .A1(n7724), .A2(net224745), .ZN(n5492) );
  NAND2_X2 U7243 ( .A1(n7726), .A2(net224745), .ZN(n5469) );
  INV_X4 U7244 ( .A(n5053), .ZN(n6068) );
  NOR2_X4 U7245 ( .A1(n7548), .A2(n3905), .ZN(n5054) );
  OAI21_X4 U7246 ( .B1(n5061), .B2(n5062), .A(n5060), .ZN(n6015) );
  INV_X4 U7247 ( .A(n5064), .ZN(n5067) );
  NAND2_X2 U7248 ( .A1(n5228), .A2(n5229), .ZN(n5070) );
  MUX2_X2 U7249 ( .A(n2897), .B(n5071), .S(net224735), .Z(n6538) );
  NAND2_X2 U7250 ( .A1(n7743), .A2(net224747), .ZN(n6811) );
  NOR2_X4 U7251 ( .A1(n6538), .A2(n5078), .ZN(n5107) );
  MUX2_X2 U7252 ( .A(n2903), .B(n6579), .S(net224735), .Z(n5079) );
  INV_X4 U7253 ( .A(n5089), .ZN(n5090) );
  NAND2_X2 U7254 ( .A1(n7745), .A2(net224745), .ZN(n5325) );
  OAI21_X4 U7255 ( .B1(n5091), .B2(n5090), .A(n5325), .ZN(n6685) );
  NAND2_X2 U7256 ( .A1(n7746), .A2(net224745), .ZN(n5443) );
  NAND2_X2 U7257 ( .A1(n5095), .A2(net224995), .ZN(n5174) );
  NAND3_X2 U7258 ( .A1(n5097), .A2(n3638), .A3(net225238), .ZN(n5369) );
  NOR2_X4 U7259 ( .A1(n7565), .A2(n3290), .ZN(n5099) );
  INV_X4 U7261 ( .A(n5117), .ZN(n5197) );
  NAND2_X2 U7262 ( .A1(n7744), .A2(net224745), .ZN(n5330) );
  NAND3_X2 U7263 ( .A1(n5197), .A2(n5196), .A3(n5366), .ZN(n5123) );
  INV_X4 U7264 ( .A(n5303), .ZN(n5125) );
  INV_X4 U7265 ( .A(n5311), .ZN(n5124) );
  INV_X4 U7266 ( .A(n5324), .ZN(n5127) );
  NAND3_X4 U7267 ( .A1(n5127), .A2(net224731), .A3(n5126), .ZN(n5128) );
  NAND2_X2 U7268 ( .A1(net33193), .A2(net224745), .ZN(n5133) );
  NOR2_X4 U7269 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  NAND2_X2 U7270 ( .A1(n7738), .A2(net224745), .ZN(n5147) );
  MUX2_X2 U7271 ( .A(n7735), .B(n5151), .S(net224735), .Z(n5159) );
  NOR3_X4 U7273 ( .A1(n5165), .A2(n5164), .A3(n5166), .ZN(n5662) );
  INV_X4 U7274 ( .A(regWrData[31]), .ZN(n5169) );
  AOI22_X2 U7275 ( .A1(n5710), .A2(n2714), .B1(n5709), .B2(memAddr[31]), .ZN(
        n5168) );
  OAI21_X4 U7276 ( .B1(n5169), .B2(n3941), .A(n5168), .ZN(n6861) );
  INV_X4 U7277 ( .A(n5173), .ZN(n5175) );
  NAND2_X2 U7278 ( .A1(n5178), .A2(net229596), .ZN(n5180) );
  NAND3_X4 U7279 ( .A1(n7737), .A2(n7746), .A3(net224743), .ZN(n5179) );
  INV_X4 U7280 ( .A(n3854), .ZN(n5184) );
  NOR3_X4 U7281 ( .A1(n5188), .A2(n5186), .A3(n2579), .ZN(n5213) );
  NAND2_X2 U7282 ( .A1(n7730), .A2(net224747), .ZN(n6381) );
  NOR3_X4 U7283 ( .A1(n5201), .A2(n5200), .A3(n5202), .ZN(n5212) );
  NOR3_X4 U7284 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(n5211) );
  MUX2_X2 U7285 ( .A(n2918), .B(n5222), .S(net224733), .Z(n6932) );
  NOR2_X4 U7286 ( .A1(n3935), .A2(n2983), .ZN(n7351) );
  NAND2_X2 U7287 ( .A1(n5710), .A2(n2751), .ZN(n5225) );
  NAND2_X2 U7288 ( .A1(n5709), .A2(memAddr[25]), .ZN(n5224) );
  NAND2_X2 U7289 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  OAI21_X4 U7290 ( .B1(n7352), .B2(n3941), .A(n5227), .ZN(n6974) );
  NAND2_X2 U7291 ( .A1(n5709), .A2(memAddr[6]), .ZN(n6223) );
  NAND2_X2 U7292 ( .A1(n5710), .A2(n2753), .ZN(n6224) );
  NAND2_X2 U7293 ( .A1(n6223), .A2(n6224), .ZN(n5232) );
  NAND2_X2 U7295 ( .A1(n5233), .A2(net224995), .ZN(n5234) );
  OAI21_X4 U7296 ( .B1(n5238), .B2(n5237), .A(n5236), .ZN(n5373) );
  NAND2_X2 U7297 ( .A1(n6661), .A2(n5876), .ZN(n5295) );
  NAND2_X2 U7298 ( .A1(n5242), .A2(net225047), .ZN(n6215) );
  NAND2_X2 U7299 ( .A1(n5710), .A2(n2755), .ZN(n6221) );
  NAND2_X2 U7300 ( .A1(n5709), .A2(memAddr[0]), .ZN(n6220) );
  NAND2_X2 U7301 ( .A1(n6221), .A2(n6220), .ZN(n5243) );
  NAND3_X4 U7302 ( .A1(reg31Val_0[0]), .A2(net224781), .A3(net225045), .ZN(
        n6216) );
  NAND3_X4 U7303 ( .A1(\wb/dsize_reg/z2 [0]), .A2(n4856), .A3(net225045), .ZN(
        n6214) );
  OAI21_X4 U7304 ( .B1(n5247), .B2(n5248), .A(n5246), .ZN(n7179) );
  OAI21_X4 U7306 ( .B1(n5481), .B2(n3941), .A(n5477), .ZN(n6335) );
  NAND2_X2 U7307 ( .A1(n3197), .A2(n3916), .ZN(n5253) );
  INV_X4 U7308 ( .A(regWrData[16]), .ZN(n5250) );
  INV_X4 U7309 ( .A(n5563), .ZN(n5249) );
  OAI21_X4 U7310 ( .B1(n5250), .B2(n3941), .A(n5249), .ZN(n7134) );
  INV_X4 U7311 ( .A(regWrData[23]), .ZN(n5255) );
  OAI21_X4 U7313 ( .B1(n5255), .B2(n3941), .A(n5254), .ZN(n7046) );
  INV_X4 U7314 ( .A(n7048), .ZN(n7044) );
  NAND2_X2 U7315 ( .A1(net225017), .A2(n3096), .ZN(n6232) );
  NOR2_X4 U7316 ( .A1(n3933), .A2(n2949), .ZN(n6229) );
  NOR2_X4 U7317 ( .A1(n2700), .A2(n2959), .ZN(n6227) );
  INV_X4 U7319 ( .A(n2617), .ZN(n5259) );
  OAI21_X4 U7320 ( .B1(n3944), .B2(n6233), .A(n3133), .ZN(n5353) );
  INV_X4 U7321 ( .A(n5353), .ZN(n5258) );
  OAI21_X4 U7322 ( .B1(n5351), .B2(n5259), .A(n5258), .ZN(n5260) );
  NAND3_X2 U7323 ( .A1(n5988), .A2(n5987), .A3(n3947), .ZN(n5732) );
  NAND2_X2 U7325 ( .A1(n3955), .A2(n6616), .ZN(n5294) );
  NOR2_X4 U7326 ( .A1(n3935), .A2(n2916), .ZN(n6093) );
  NAND2_X2 U7327 ( .A1(n6093), .A2(n3945), .ZN(n5267) );
  OAI22_X2 U7328 ( .A1(n7695), .A2(n3909), .B1(n7422), .B2(n3911), .ZN(n6101)
         );
  NAND3_X4 U7329 ( .A1(n5267), .A2(n5266), .A3(n5265), .ZN(n6359) );
  NAND2_X2 U7330 ( .A1(n6359), .A2(net225029), .ZN(n6125) );
  INV_X4 U7331 ( .A(n6125), .ZN(n6394) );
  NAND3_X2 U7332 ( .A1(n6192), .A2(n6193), .A3(n3947), .ZN(n5873) );
  NAND2_X2 U7333 ( .A1(n5873), .A2(n5967), .ZN(n5278) );
  INV_X4 U7334 ( .A(n5268), .ZN(n5269) );
  AOI21_X4 U7335 ( .B1(n5270), .B2(net224993), .A(n5269), .ZN(n6245) );
  NOR2_X4 U7336 ( .A1(n7560), .A2(n3905), .ZN(n5273) );
  NAND3_X2 U7337 ( .A1(n5276), .A2(n6184), .A3(n3947), .ZN(n5872) );
  NAND2_X2 U7338 ( .A1(n5872), .A2(n6944), .ZN(n5277) );
  NAND3_X4 U7339 ( .A1(n5278), .A2(n5734), .A3(n5277), .ZN(n5762) );
  NAND2_X2 U7340 ( .A1(n7176), .A2(n5762), .ZN(n5293) );
  NOR2_X4 U7341 ( .A1(n3936), .A2(n2981), .ZN(n6250) );
  NAND2_X2 U7342 ( .A1(n5710), .A2(n2750), .ZN(n6254) );
  NOR2_X4 U7343 ( .A1(n6250), .A2(n5280), .ZN(n5279) );
  INV_X4 U7344 ( .A(n5279), .ZN(n5283) );
  INV_X4 U7345 ( .A(n5280), .ZN(n5281) );
  AOI21_X4 U7346 ( .B1(n5281), .B2(n3941), .A(net225083), .ZN(n5282) );
  OAI21_X4 U7347 ( .B1(n6249), .B2(n5283), .A(n5282), .ZN(n6634) );
  NAND2_X2 U7348 ( .A1(n6791), .A2(net225029), .ZN(n6793) );
  INV_X4 U7349 ( .A(n6793), .ZN(n6788) );
  NAND3_X2 U7350 ( .A1(n3699), .A2(n3947), .A3(n5977), .ZN(n5998) );
  NAND2_X2 U7351 ( .A1(n5967), .A2(n5998), .ZN(n5291) );
  INV_X4 U7352 ( .A(regWrData[21]), .ZN(n5286) );
  OAI21_X4 U7354 ( .B1(n5286), .B2(n3941), .A(n5285), .ZN(n6342) );
  NAND2_X2 U7355 ( .A1(n6342), .A2(net225029), .ZN(n5940) );
  INV_X4 U7356 ( .A(n5940), .ZN(n7108) );
  INV_X4 U7358 ( .A(n5398), .ZN(n5799) );
  OAI21_X4 U7359 ( .B1(n8010), .B2(n3941), .A(n5799), .ZN(n6485) );
  INV_X4 U7360 ( .A(n6502), .ZN(n6504) );
  NAND2_X2 U7361 ( .A1(n6944), .A2(n7168), .ZN(n5290) );
  NAND3_X4 U7362 ( .A1(n5291), .A2(n5290), .A3(n5734), .ZN(n5864) );
  INV_X4 U7363 ( .A(n5658), .ZN(n5302) );
  OAI22_X2 U7364 ( .A1(n7542), .A2(n3901), .B1(net225243), .B2(n7685), .ZN(
        n6298) );
  NAND2_X2 U7365 ( .A1(n5600), .A2(n5605), .ZN(n5300) );
  NAND2_X2 U7366 ( .A1(n5599), .A2(n5605), .ZN(n5299) );
  NAND2_X2 U7367 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  AOI21_X4 U7368 ( .B1(n5306), .B2(n5305), .A(n5304), .ZN(n5307) );
  OAI21_X4 U7369 ( .B1(n5316), .B2(n5315), .A(n5314), .ZN(n6688) );
  AOI21_X4 U7370 ( .B1(n5321), .B2(n4718), .A(n5320), .ZN(n5322) );
  NAND2_X2 U7371 ( .A1(n5325), .A2(net224747), .ZN(n5326) );
  OAI21_X4 U7372 ( .B1(n5327), .B2(n5328), .A(n5326), .ZN(n5329) );
  AOI21_X4 U7373 ( .B1(n5336), .B2(n5335), .A(n5342), .ZN(n5456) );
  NAND3_X4 U7374 ( .A1(n5456), .A2(n5457), .A3(n6583), .ZN(n6824) );
  NAND3_X4 U7375 ( .A1(n5350), .A2(n5349), .A3(n5348), .ZN(n5453) );
  INV_X4 U7376 ( .A(n5351), .ZN(n5354) );
  OAI22_X2 U7377 ( .A1(n7533), .A2(n3911), .B1(n7686), .B2(n3909), .ZN(n5355)
         );
  NAND2_X2 U7378 ( .A1(n5356), .A2(\wb/dsize_reg/z2 [25]), .ZN(n6238) );
  INV_X4 U7379 ( .A(n6238), .ZN(n5357) );
  NAND2_X2 U7380 ( .A1(n5357), .A2(net225047), .ZN(n5362) );
  XNOR2_X2 U7382 ( .A(n5367), .B(n5366), .ZN(n5458) );
  XNOR2_X2 U7383 ( .A(n5373), .B(net224861), .ZN(n5793) );
  XNOR2_X2 U7384 ( .A(n5374), .B(n5793), .ZN(n5375) );
  INV_X4 U7385 ( .A(n5383), .ZN(n5384) );
  INV_X4 U7386 ( .A(n5387), .ZN(n5388) );
  AOI221_X2 U7387 ( .B1(n5398), .B2(net225029), .C1(n5397), .C2(n2672), .A(
        n5896), .ZN(n5434) );
  NAND3_X2 U7388 ( .A1(regWrData[11]), .A2(n3133), .A3(n3945), .ZN(n5399) );
  NAND2_X2 U7389 ( .A1(n5713), .A2(net225029), .ZN(n5500) );
  INV_X4 U7390 ( .A(n5402), .ZN(n5699) );
  AOI21_X4 U7391 ( .B1(n5699), .B2(n3941), .A(net225083), .ZN(n5406) );
  NAND3_X4 U7392 ( .A1(n5404), .A2(n5403), .A3(n5699), .ZN(n5405) );
  NOR3_X4 U7393 ( .A1(n7973), .A2(n3920), .A3(net225015), .ZN(n5419) );
  XNOR2_X2 U7394 ( .A(net224869), .B(n7722), .ZN(n5423) );
  INV_X4 U7395 ( .A(n5443), .ZN(n5444) );
  AOI21_X4 U7396 ( .B1(n5445), .B2(net224731), .A(n5444), .ZN(n5446) );
  XNOR2_X2 U7397 ( .A(n5448), .B(net224861), .ZN(n5449) );
  NOR2_X4 U7398 ( .A1(n6588), .A2(n5450), .ZN(n5466) );
  OAI21_X4 U7399 ( .B1(n5465), .B2(n5466), .A(n5464), .ZN(n6155) );
  INV_X4 U7400 ( .A(net222515), .ZN(net221442) );
  XNOR2_X2 U7401 ( .A(net227791), .B(n5469), .ZN(n5471) );
  NOR2_X4 U7402 ( .A1(net225083), .A2(net224871), .ZN(n5634) );
  NAND2_X2 U7403 ( .A1(n5477), .A2(net224859), .ZN(n5478) );
  NAND2_X2 U7404 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  XNOR2_X2 U7405 ( .A(n5486), .B(net224865), .ZN(n5489) );
  NAND2_X2 U7406 ( .A1(n5492), .A2(n7946), .ZN(n5496) );
  XNOR2_X2 U7407 ( .A(n5497), .B(net228323), .ZN(n5504) );
  NAND2_X2 U7408 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NOR2_X4 U7409 ( .A1(n2989), .A2(n5502), .ZN(n5503) );
  OAI21_X4 U7410 ( .B1(n2591), .B2(n6714), .A(n6548), .ZN(n6524) );
  NAND3_X4 U7411 ( .A1(n6524), .A2(n3698), .A3(n3629), .ZN(n6152) );
  XNOR2_X2 U7412 ( .A(n3360), .B(n5506), .ZN(n6530) );
  OAI21_X4 U7413 ( .B1(n5510), .B2(n5902), .A(n5911), .ZN(n5808) );
  NAND3_X4 U7414 ( .A1(n7144), .A2(n6152), .A3(n5813), .ZN(n7054) );
  NOR2_X4 U7415 ( .A1(n5548), .A2(n5547), .ZN(n5516) );
  INV_X4 U7416 ( .A(n5514), .ZN(n5690) );
  AOI21_X4 U7417 ( .B1(n5516), .B2(n5690), .A(n5515), .ZN(n5540) );
  NAND3_X2 U7418 ( .A1(n5518), .A2(n5523), .A3(n5527), .ZN(n5520) );
  INV_X4 U7419 ( .A(n5523), .ZN(n5524) );
  INV_X4 U7420 ( .A(n5527), .ZN(n5528) );
  NAND3_X2 U7421 ( .A1(n5534), .A2(n3200), .A3(n6400), .ZN(n5535) );
  NOR3_X4 U7422 ( .A1(n5542), .A2(n6702), .A3(n3769), .ZN(n5557) );
  NAND3_X4 U7423 ( .A1(n5543), .A2(n5544), .A3(n5545), .ZN(n5642) );
  XNOR2_X2 U7424 ( .A(n5642), .B(net224859), .ZN(n5546) );
  AOI22_X2 U7425 ( .A1(n3945), .A2(n5548), .B1(n3945), .B2(n5547), .ZN(n5549)
         );
  AOI21_X4 U7426 ( .B1(n5549), .B2(n5690), .A(net225084), .ZN(n5550) );
  NOR2_X4 U7427 ( .A1(n6594), .A2(n5462), .ZN(n5552) );
  NAND3_X2 U7428 ( .A1(n5556), .A2(n5557), .A3(n2621), .ZN(n5809) );
  INV_X4 U7429 ( .A(n5558), .ZN(n5559) );
  INV_X4 U7430 ( .A(n5560), .ZN(n5562) );
  NAND2_X2 U7431 ( .A1(n3652), .A2(n7136), .ZN(n5647) );
  INV_X4 U7432 ( .A(n5567), .ZN(n5569) );
  NOR2_X4 U7433 ( .A1(n5568), .A2(n5569), .ZN(n5570) );
  NAND2_X2 U7434 ( .A1(net225029), .A2(n5571), .ZN(n5618) );
  INV_X4 U7435 ( .A(n5578), .ZN(n6206) );
  NAND2_X2 U7436 ( .A1(n6206), .A2(n5575), .ZN(n5576) );
  AOI21_X4 U7437 ( .B1(n5581), .B2(n5580), .A(n5579), .ZN(n6758) );
  NAND2_X2 U7438 ( .A1(n5710), .A2(n2754), .ZN(n6210) );
  NAND2_X2 U7439 ( .A1(n5588), .A2(n5587), .ZN(n5591) );
  AOI21_X4 U7440 ( .B1(n5589), .B2(n3941), .A(net225083), .ZN(n5590) );
  OAI21_X4 U7441 ( .B1(n5592), .B2(n5591), .A(n5590), .ZN(n6770) );
  AOI22_X2 U7442 ( .A1(n5596), .A2(n5595), .B1(n5595), .B2(n5594), .ZN(n5597)
         );
  XNOR2_X2 U7443 ( .A(n5597), .B(net224859), .ZN(n5598) );
  NAND3_X2 U7444 ( .A1(n6750), .A2(n6678), .A3(n6748), .ZN(n5811) );
  NAND2_X2 U7446 ( .A1(n7733), .A2(net224747), .ZN(n5602) );
  NAND2_X2 U7447 ( .A1(n5602), .A2(net224861), .ZN(n5603) );
  NOR2_X4 U7448 ( .A1(n5604), .A2(n5603), .ZN(n5610) );
  XNOR2_X2 U7449 ( .A(n6770), .B(net224861), .ZN(n5611) );
  INV_X4 U7450 ( .A(n5624), .ZN(n5614) );
  NAND2_X2 U7451 ( .A1(n5614), .A2(n5613), .ZN(n5617) );
  NAND2_X2 U7452 ( .A1(n5618), .A2(net224871), .ZN(n5619) );
  INV_X4 U7453 ( .A(n5619), .ZN(n5623) );
  AOI211_X4 U7454 ( .C1(n5620), .C2(n3940), .A(net225084), .B(net224871), .ZN(
        n5622) );
  OAI21_X4 U7455 ( .B1(n5623), .B2(n5622), .A(n5621), .ZN(n5628) );
  NOR3_X4 U7456 ( .A1(n5627), .A2(n5628), .A3(n5629), .ZN(n5630) );
  AOI21_X4 U7458 ( .B1(n6751), .B2(n6750), .A(n5633), .ZN(n6011) );
  XNOR2_X2 U7459 ( .A(n5643), .B(n5642), .ZN(n6837) );
  OAI21_X4 U7460 ( .B1(n6011), .B2(n5644), .A(n3241), .ZN(n5645) );
  INV_X4 U7461 ( .A(n7156), .ZN(n7150) );
  INV_X4 U7462 ( .A(n5650), .ZN(n5651) );
  NOR2_X4 U7463 ( .A1(n5652), .A2(n5651), .ZN(n5656) );
  AOI21_X4 U7464 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5657) );
  XNOR2_X2 U7465 ( .A(n5657), .B(net224865), .ZN(net222370) );
  NAND2_X2 U7466 ( .A1(n6683), .A2(n6462), .ZN(n6954) );
  INV_X4 U7468 ( .A(n5661), .ZN(n5660) );
  NOR2_X4 U7469 ( .A1(n2700), .A2(n2982), .ZN(n5659) );
  INV_X4 U7470 ( .A(n5659), .ZN(n7348) );
  NAND2_X2 U7471 ( .A1(n5660), .A2(n3942), .ZN(n6046) );
  NAND3_X2 U7472 ( .A1(n6954), .A2(n6955), .A3(n3947), .ZN(n5946) );
  NAND3_X2 U7474 ( .A1(n6951), .A2(n6950), .A3(n3947), .ZN(n5948) );
  INV_X4 U7475 ( .A(n6514), .ZN(n5722) );
  INV_X4 U7476 ( .A(n5666), .ZN(n6260) );
  NAND2_X2 U7477 ( .A1(n6260), .A2(n6258), .ZN(n5673) );
  OAI21_X4 U7478 ( .B1(n5673), .B2(n6257), .A(n5672), .ZN(n6423) );
  NAND3_X2 U7479 ( .A1(n5679), .A2(n5678), .A3(n2649), .ZN(n5929) );
  AOI22_X2 U7480 ( .A1(n5710), .A2(n2716), .B1(n5709), .B2(memAddr[22]), .ZN(
        n5680) );
  OAI21_X4 U7481 ( .B1(n5681), .B2(n3940), .A(n5680), .ZN(n7074) );
  NAND2_X2 U7482 ( .A1(n5989), .A2(net220656), .ZN(n5931) );
  NAND2_X2 U7483 ( .A1(n6810), .A2(n6462), .ZN(n5930) );
  NAND3_X2 U7484 ( .A1(n5930), .A2(n5931), .A3(n3947), .ZN(n5725) );
  NAND2_X2 U7485 ( .A1(n5967), .A2(n5725), .ZN(n5682) );
  NAND3_X4 U7486 ( .A1(n5683), .A2(n5969), .A3(n5682), .ZN(n6620) );
  INV_X4 U7487 ( .A(n6031), .ZN(n5684) );
  NAND2_X2 U7488 ( .A1(n5684), .A2(n3945), .ZN(n5689) );
  NOR2_X4 U7489 ( .A1(n3936), .A2(n2960), .ZN(n6028) );
  NAND2_X2 U7490 ( .A1(n6028), .A2(n3945), .ZN(n5688) );
  NAND2_X2 U7491 ( .A1(n3934), .A2(\wb/dsize_reg/z2 [26]), .ZN(n6029) );
  INV_X4 U7492 ( .A(n6029), .ZN(n5686) );
  NAND2_X2 U7493 ( .A1(n6341), .A2(net225029), .ZN(n6017) );
  INV_X4 U7494 ( .A(n6017), .ZN(n6013) );
  NAND2_X2 U7495 ( .A1(n6462), .A2(n6013), .ZN(n6458) );
  OAI22_X2 U7496 ( .A1(n7544), .A2(net225015), .B1(n2734), .B2(n2699), .ZN(
        n5694) );
  INV_X4 U7497 ( .A(n5694), .ZN(n7346) );
  NOR2_X4 U7498 ( .A1(n3935), .A2(n2974), .ZN(n7345) );
  NAND2_X2 U7499 ( .A1(n5710), .A2(n2752), .ZN(n5696) );
  NAND2_X2 U7500 ( .A1(n5709), .A2(memAddr[18]), .ZN(n5695) );
  NAND2_X2 U7501 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  AOI21_X4 U7502 ( .B1(n3944), .B2(n7345), .A(n5697), .ZN(n5698) );
  OAI21_X4 U7503 ( .B1(n7346), .B2(n3940), .A(n5698), .ZN(n6343) );
  INV_X4 U7504 ( .A(n5776), .ZN(n5841) );
  INV_X4 U7506 ( .A(regWrData[13]), .ZN(n5700) );
  NAND2_X2 U7507 ( .A1(n6533), .A2(net225029), .ZN(n6535) );
  INV_X4 U7508 ( .A(n6535), .ZN(n6522) );
  NAND2_X2 U7510 ( .A1(n6944), .A2(n6457), .ZN(n5703) );
  INV_X4 U7512 ( .A(n6188), .ZN(n6406) );
  NAND3_X2 U7513 ( .A1(n5854), .A2(n5855), .A3(n3947), .ZN(n6004) );
  AOI22_X2 U7515 ( .A1(n5710), .A2(n2717), .B1(n5709), .B2(memAddr[20]), .ZN(
        n5711) );
  OAI21_X4 U7516 ( .B1(n5712), .B2(n3940), .A(n5711), .ZN(n6357) );
  AOI22_X2 U7518 ( .A1(n5860), .A2(n7176), .B1(n5835), .B2(n7239), .ZN(n5720)
         );
  INV_X4 U7519 ( .A(n5730), .ZN(n5723) );
  NAND2_X2 U7520 ( .A1(n6003), .A2(n5967), .ZN(n5727) );
  NAND2_X2 U7521 ( .A1(n3955), .A2(n5876), .ZN(n5739) );
  NAND2_X2 U7522 ( .A1(n5967), .A2(n5731), .ZN(n5735) );
  NAND2_X2 U7523 ( .A1(n5732), .A2(n6944), .ZN(n5733) );
  NAND3_X4 U7524 ( .A1(n5735), .A2(n5734), .A3(n5733), .ZN(n6600) );
  NAND2_X2 U7525 ( .A1(n7239), .A2(n6600), .ZN(n5738) );
  NAND2_X2 U7526 ( .A1(n6661), .A2(n5762), .ZN(n5737) );
  NAND2_X2 U7527 ( .A1(n7176), .A2(n5864), .ZN(n5736) );
  MUX2_X2 U7528 ( .A(net224851), .B(n3913), .S(n5841), .Z(n5745) );
  NAND2_X2 U7529 ( .A1(n5745), .A2(n2838), .ZN(n5757) );
  NAND2_X2 U7530 ( .A1(n7176), .A2(n6600), .ZN(n5750) );
  INV_X4 U7531 ( .A(n7941), .ZN(n6005) );
  OAI21_X4 U7532 ( .B1(n6005), .B2(n5960), .A(n3922), .ZN(n6668) );
  INV_X4 U7533 ( .A(n6668), .ZN(n5746) );
  NAND2_X2 U7534 ( .A1(n5746), .A2(n7239), .ZN(n5749) );
  NOR2_X4 U7535 ( .A1(n6546), .A2(n3954), .ZN(n5755) );
  AOI211_X4 U7536 ( .C1(n5757), .C2(n5756), .A(n5754), .B(n5755), .ZN(n5786)
         );
  NAND2_X2 U7537 ( .A1(n6661), .A2(n6616), .ZN(n5765) );
  NAND2_X2 U7538 ( .A1(n3916), .A2(n5972), .ZN(n5950) );
  AOI22_X2 U7539 ( .A1(n7169), .A2(n5998), .B1(n7168), .B2(n5967), .ZN(n5760)
         );
  NAND2_X2 U7541 ( .A1(n7127), .A2(n7918), .ZN(n5784) );
  INV_X4 U7542 ( .A(n5766), .ZN(n5782) );
  INV_X4 U7543 ( .A(n5767), .ZN(n5768) );
  INV_X4 U7544 ( .A(n5771), .ZN(n5772) );
  AOI21_X4 U7545 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  XNOR2_X2 U7546 ( .A(n5775), .B(net227884), .ZN(n5840) );
  XNOR2_X2 U7547 ( .A(n5840), .B(n5776), .ZN(n6909) );
  NAND4_X2 U7548 ( .A1(n5784), .A2(n5786), .A3(n5783), .A4(n5785), .ZN(
        \ex_mem/N214 ) );
  AOI22_X2 U7549 ( .A1(n7127), .A2(n7133), .B1(n3924), .B2(n2690), .ZN(n5828)
         );
  NAND2_X2 U7550 ( .A1(n3954), .A2(n2701), .ZN(n5825) );
  NAND2_X2 U7551 ( .A1(n6661), .A2(n5860), .ZN(n5791) );
  INV_X4 U7552 ( .A(n5890), .ZN(n5792) );
  INV_X4 U7553 ( .A(n6698), .ZN(n6550) );
  INV_X4 U7554 ( .A(n6156), .ZN(n5806) );
  NAND2_X2 U7555 ( .A1(n3945), .A2(n5798), .ZN(n5800) );
  OAI211_X2 U7556 ( .C1(n5801), .C2(n3942), .A(n5800), .B(n5799), .ZN(n5802)
         );
  NAND2_X2 U7557 ( .A1(n5802), .A2(net225029), .ZN(n5804) );
  XNOR2_X2 U7558 ( .A(n5804), .B(n5803), .ZN(n6552) );
  INV_X4 U7559 ( .A(n6552), .ZN(n5805) );
  OAI21_X4 U7560 ( .B1(n6550), .B2(n5806), .A(n5805), .ZN(n5807) );
  OAI21_X4 U7561 ( .B1(n5646), .B2(n7984), .A(n5810), .ZN(n6558) );
  XNOR2_X2 U7562 ( .A(n5815), .B(n7142), .ZN(n7308) );
  MUX2_X2 U7563 ( .A(net224843), .B(n7151), .S(n3197), .Z(n5817) );
  NAND3_X2 U7564 ( .A1(n5826), .A2(n5828), .A3(n5827), .ZN(\ex_mem/N211 ) );
  INV_X4 U7565 ( .A(n6357), .ZN(n5829) );
  MUX2_X2 U7566 ( .A(net224843), .B(n7151), .S(n6040), .Z(n5832) );
  OAI21_X4 U7567 ( .B1(n3763), .B2(n6005), .A(n3922), .ZN(n6610) );
  NAND2_X2 U7571 ( .A1(net222151), .A2(n7020), .ZN(n5845) );
  NAND2_X2 U7572 ( .A1(net222151), .A2(n7004), .ZN(n5844) );
  XNOR2_X2 U7573 ( .A(n5847), .B(n5871), .ZN(net221922) );
  XNOR2_X2 U7574 ( .A(n5848), .B(net228341), .ZN(n7324) );
  NAND3_X2 U7575 ( .A1(n3916), .A2(n5972), .A3(net221494), .ZN(n5851) );
  INV_X4 U7576 ( .A(n5854), .ZN(n5857) );
  INV_X4 U7577 ( .A(n5855), .ZN(n5856) );
  OAI21_X4 U7578 ( .B1(n5857), .B2(n5856), .A(n7242), .ZN(n7226) );
  AOI22_X2 U7579 ( .A1(n7239), .A2(n5860), .B1(n3955), .B2(n2696), .ZN(n5862)
         );
  NAND2_X2 U7580 ( .A1(n5746), .A2(n7176), .ZN(n5868) );
  NAND2_X2 U7581 ( .A1(n7239), .A2(n6602), .ZN(n5867) );
  NAND2_X2 U7582 ( .A1(n6661), .A2(n6600), .ZN(n5866) );
  NAND2_X2 U7583 ( .A1(n3955), .A2(n5864), .ZN(n5865) );
  AOI22_X2 U7584 ( .A1(n7169), .A2(n5873), .B1(n5967), .B2(n5872), .ZN(n5874)
         );
  NAND2_X2 U7585 ( .A1(n7239), .A2(n5876), .ZN(n5878) );
  NAND2_X2 U7586 ( .A1(n7176), .A2(n6616), .ZN(n5877) );
  MUX2_X2 U7587 ( .A(net224853), .B(n7182), .S(n5886), .Z(n5887) );
  NAND2_X2 U7588 ( .A1(n5887), .A2(n2838), .ZN(n5919) );
  INV_X4 U7589 ( .A(n6489), .ZN(n5894) );
  AOI211_X4 U7590 ( .C1(n5901), .C2(n5900), .A(n5898), .B(n5899), .ZN(n6525)
         );
  NAND2_X2 U7591 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  NAND2_X2 U7592 ( .A1(n6699), .A2(n6705), .ZN(n6557) );
  INV_X4 U7593 ( .A(n6557), .ZN(n5906) );
  XNOR2_X2 U7594 ( .A(n3544), .B(n5910), .ZN(n7284) );
  NAND4_X2 U7596 ( .A1(n5921), .A2(n5923), .A3(n5920), .A4(n5922), .ZN(
        \ex_mem/N210 ) );
  INV_X4 U7597 ( .A(n6342), .ZN(n7124) );
  INV_X4 U7598 ( .A(n7046), .ZN(n5926) );
  INV_X4 U7599 ( .A(n6974), .ZN(n6351) );
  INV_X4 U7600 ( .A(n6341), .ZN(n5928) );
  NAND3_X2 U7601 ( .A1(n5931), .A2(n3947), .A3(n5930), .ZN(n5932) );
  NAND2_X2 U7602 ( .A1(n7169), .A2(n5932), .ZN(n6443) );
  NAND2_X2 U7603 ( .A1(n5938), .A2(n5937), .ZN(n6469) );
  OAI21_X4 U7604 ( .B1(n5939), .B2(n3916), .A(n6469), .ZN(n5943) );
  OAI21_X4 U7605 ( .B1(n5943), .B2(n5942), .A(n7201), .ZN(n5945) );
  NAND2_X2 U7606 ( .A1(n5967), .A2(n6457), .ZN(n5944) );
  INV_X4 U7607 ( .A(n5951), .ZN(n5952) );
  INV_X4 U7608 ( .A(n6427), .ZN(n5964) );
  NAND2_X2 U7609 ( .A1(n5962), .A2(n5989), .ZN(n6426) );
  INV_X4 U7610 ( .A(n6426), .ZN(n5963) );
  NOR2_X4 U7611 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  NAND3_X4 U7612 ( .A1(n5970), .A2(n5968), .A3(n7935), .ZN(n6660) );
  INV_X4 U7613 ( .A(n3878), .ZN(n6618) );
  INV_X4 U7614 ( .A(n6080), .ZN(n6114) );
  INV_X4 U7616 ( .A(n5977), .ZN(n5978) );
  INV_X4 U7617 ( .A(n7175), .ZN(n5982) );
  INV_X4 U7618 ( .A(n3850), .ZN(n5994) );
  NAND2_X2 U7619 ( .A1(n7027), .A2(n6944), .ZN(n5990) );
  NOR2_X4 U7620 ( .A1(n3521), .A2(n5991), .ZN(n5992) );
  AOI22_X2 U7621 ( .A1(n3955), .A2(n2681), .B1(n3747), .B2(n6661), .ZN(n5995)
         );
  NAND2_X2 U7622 ( .A1(n7176), .A2(n6669), .ZN(n6002) );
  OAI21_X4 U7623 ( .B1(n6005), .B2(n5998), .A(n3922), .ZN(n6671) );
  INV_X4 U7624 ( .A(n6671), .ZN(n6169) );
  NAND2_X2 U7625 ( .A1(n6169), .A2(n6661), .ZN(n6001) );
  NAND2_X2 U7626 ( .A1(n7239), .A2(n7255), .ZN(n6006) );
  INV_X4 U7627 ( .A(n6006), .ZN(n5999) );
  NAND3_X4 U7628 ( .A1(n6002), .A2(n6001), .A3(n6000), .ZN(n6851) );
  OAI21_X4 U7629 ( .B1(n6005), .B2(n6003), .A(n3922), .ZN(n6606) );
  OAI21_X4 U7630 ( .B1(n6004), .B2(n6005), .A(n3922), .ZN(n6607) );
  NOR3_X4 U7631 ( .A1(n6007), .A2(n6008), .A3(n6009), .ZN(n6980) );
  MUX2_X2 U7632 ( .A(net224851), .B(n3913), .S(n6013), .Z(n6014) );
  NAND2_X2 U7633 ( .A1(n7358), .A2(n6341), .ZN(n6016) );
  OAI221_X2 U7634 ( .B1(n3274), .B2(n3954), .C1(n6086), .C2(n3923), .A(n6026), 
        .ZN(\ex_mem/N200 ) );
  INV_X4 U7635 ( .A(n6340), .ZN(n6027) );
  INV_X4 U7636 ( .A(n6028), .ZN(n6030) );
  NAND3_X4 U7637 ( .A1(n6031), .A2(n6030), .A3(n6029), .ZN(regWrData[26]) );
  NOR2_X4 U7638 ( .A1(n6033), .A2(n6034), .ZN(n6036) );
  OAI21_X4 U7639 ( .B1(n6037), .B2(n6036), .A(n6035), .ZN(net221806) );
  NAND3_X4 U7640 ( .A1(net221481), .A2(n3411), .A3(n6373), .ZN(net220767) );
  INV_X4 U7641 ( .A(n6049), .ZN(n6050) );
  INV_X4 U7642 ( .A(n6051), .ZN(n6052) );
  NOR2_X4 U7643 ( .A1(n6053), .A2(n6052), .ZN(n6056) );
  AOI21_X4 U7644 ( .B1(n6057), .B2(n6056), .A(n6055), .ZN(net221905) );
  XNOR2_X2 U7646 ( .A(n6063), .B(net224865), .ZN(n6064) );
  XNOR2_X2 U7647 ( .A(n6065), .B(n6066), .ZN(net220720) );
  INV_X4 U7649 ( .A(regWrData[26]), .ZN(n6076) );
  INV_X4 U7650 ( .A(n6070), .ZN(n6071) );
  MUX2_X2 U7651 ( .A(net224853), .B(n7182), .S(n6114), .Z(net221862) );
  NAND2_X2 U7652 ( .A1(n7358), .A2(n6340), .ZN(n6079) );
  OAI221_X2 U7653 ( .B1(n3274), .B2(n3918), .C1(n6086), .C2(n2701), .A(n6085), 
        .ZN(\ex_mem/N222 ) );
  INV_X4 U7654 ( .A(n6359), .ZN(n6094) );
  NAND2_X2 U7655 ( .A1(n6088), .A2(net224995), .ZN(n6092) );
  NOR2_X4 U7656 ( .A1(n6093), .A2(n6104), .ZN(n6106) );
  MUX2_X2 U7657 ( .A(net224843), .B(n7151), .S(n6394), .Z(n6097) );
  INV_X4 U7658 ( .A(n6607), .ZN(n6098) );
  NAND2_X2 U7659 ( .A1(n7255), .A2(n3649), .ZN(n6170) );
  OAI22_X2 U7660 ( .A1(n6836), .A2(n3954), .B1(n6100), .B2(n3923), .ZN(n6123)
         );
  OAI211_X2 U7661 ( .C1(n3945), .C2(n3508), .A(net225029), .B(net224865), .ZN(
        n6103) );
  INV_X4 U7662 ( .A(n6101), .ZN(n6107) );
  OAI21_X4 U7663 ( .B1(n6107), .B2(net225083), .A(net224861), .ZN(n6102) );
  NAND2_X2 U7665 ( .A1(n6105), .A2(n6104), .ZN(n6109) );
  INV_X4 U7667 ( .A(n6115), .ZN(n6116) );
  OAI21_X4 U7668 ( .B1(n6991), .B2(n6116), .A(n6117), .ZN(net221802) );
  NAND2_X2 U7669 ( .A1(n6663), .A2(n6478), .ZN(n6132) );
  NAND2_X2 U7670 ( .A1(n7176), .A2(n6622), .ZN(n6131) );
  NAND2_X2 U7671 ( .A1(n6661), .A2(n6129), .ZN(n6130) );
  NAND4_X2 U7672 ( .A1(n6134), .A2(n6136), .A3(n6135), .A4(n6137), .ZN(
        \ex_mem/N223 ) );
  INV_X4 U7674 ( .A(net221763), .ZN(net221762) );
  NOR2_X4 U7675 ( .A1(net221762), .A2(net227982), .ZN(n6144) );
  NAND2_X2 U7676 ( .A1(n6145), .A2(net220644), .ZN(n6146) );
  NOR2_X4 U7677 ( .A1(n3416), .A2(n3042), .ZN(n6646) );
  NAND2_X2 U7679 ( .A1(n6661), .A2(n6669), .ZN(n6172) );
  NAND2_X2 U7680 ( .A1(n6169), .A2(n6663), .ZN(n6171) );
  INV_X4 U7681 ( .A(n6801), .ZN(n6766) );
  NOR2_X4 U7682 ( .A1(n6766), .A2(n3954), .ZN(n6182) );
  MUX2_X2 U7683 ( .A(net224853), .B(n3913), .S(n6406), .Z(n6173) );
  OAI21_X4 U7684 ( .B1(n6836), .B2(n3923), .A(n6180), .ZN(n6181) );
  INV_X4 U7686 ( .A(n6193), .ZN(n6194) );
  OAI21_X4 U7687 ( .B1(n6195), .B2(n6194), .A(n6956), .ZN(n6196) );
  INV_X4 U7688 ( .A(regWrData[3]), .ZN(n6207) );
  INV_X4 U7689 ( .A(n6356), .ZN(n6757) );
  INV_X4 U7690 ( .A(n6791), .ZN(n6208) );
  INV_X4 U7691 ( .A(n6783), .ZN(n6211) );
  INV_X4 U7692 ( .A(n6219), .ZN(regWrData[0]) );
  OAI211_X2 U7693 ( .C1(n6219), .C2(n3942), .A(n6221), .B(n6220), .ZN(n7190)
         );
  INV_X4 U7694 ( .A(n7190), .ZN(n6222) );
  INV_X4 U7695 ( .A(regWrData[6]), .ZN(n6225) );
  INV_X4 U7696 ( .A(n6350), .ZN(n6736) );
  INV_X4 U7697 ( .A(n6686), .ZN(n6226) );
  INV_X4 U7698 ( .A(n6227), .ZN(n6231) );
  INV_X4 U7699 ( .A(regWrData[8]), .ZN(n6235) );
  INV_X4 U7700 ( .A(n3644), .ZN(n6234) );
  INV_X4 U7701 ( .A(n6334), .ZN(n6580) );
  INV_X4 U7702 ( .A(n6237), .ZN(n6240) );
  INV_X4 U7703 ( .A(regWrData[9]), .ZN(n6243) );
  INV_X4 U7704 ( .A(n6815), .ZN(n6244) );
  INV_X4 U7705 ( .A(n6358), .ZN(n6717) );
  INV_X4 U7706 ( .A(regWrData[12]), .ZN(n6247) );
  INV_X4 U7707 ( .A(n6355), .ZN(n6565) );
  INV_X4 U7708 ( .A(n6533), .ZN(n6248) );
  INV_X4 U7709 ( .A(n6250), .ZN(n6251) );
  NAND2_X2 U7710 ( .A1(n6252), .A2(n6251), .ZN(regWrData[29]) );
  INV_X4 U7711 ( .A(regWrData[29]), .ZN(n6255) );
  OAI211_X2 U7712 ( .C1(n6255), .C2(n3942), .A(n6254), .B(n6253), .ZN(n6632)
         );
  INV_X4 U7713 ( .A(n6632), .ZN(n6256) );
  NAND2_X2 U7714 ( .A1(n6259), .A2(n6258), .ZN(regWrData[30]) );
  INV_X4 U7715 ( .A(regWrData[30]), .ZN(n6262) );
  INV_X4 U7716 ( .A(n6422), .ZN(n6263) );
  NAND3_X2 U7717 ( .A1(n2738), .A2(n2836), .A3(n3085), .ZN(n6265) );
  NOR4_X2 U7718 ( .A1(n6265), .A2(n7622), .A3(n7623), .A4(n7619), .ZN(n6276)
         );
  NOR4_X2 U7719 ( .A1(n3117), .A2(instr_2[27]), .A3(instr_2[26]), .A4(
        instr_2[17]), .ZN(n6275) );
  NAND2_X2 U7720 ( .A1(valid_3), .A2(n6268), .ZN(n6294) );
  INV_X4 U7721 ( .A(n6294), .ZN(n6287) );
  XNOR2_X2 U7722 ( .A(rd_3[1]), .B(rd_2[1]), .ZN(n6270) );
  NAND4_X2 U7723 ( .A1(n7618), .A2(n6287), .A3(n6270), .A4(n6269), .ZN(n6273)
         );
  NAND3_X2 U7724 ( .A1(n6276), .A2(n6275), .A3(n6274), .ZN(n6297) );
  INV_X4 U7725 ( .A(n6297), .ZN(n6277) );
  NOR2_X4 U7726 ( .A1(rs1[3]), .A2(net224955), .ZN(n6278) );
  MUX2_X2 U7727 ( .A(n6278), .B(n2926), .S(rd_3[3]), .Z(n6286) );
  XOR2_X2 U7728 ( .A(rs1[2]), .B(rd_3[2]), .Z(n6279) );
  XOR2_X2 U7729 ( .A(rd_3[4]), .B(rs1[4]), .Z(n6283) );
  XOR2_X2 U7730 ( .A(rd_3[1]), .B(rs1[1]), .Z(n6282) );
  XOR2_X2 U7731 ( .A(rs1[0]), .B(rd_3[0]), .Z(n6281) );
  XNOR2_X2 U7732 ( .A(rd_3[3]), .B(\hazard_detect/eq_83/A[3] ), .ZN(n6290) );
  XNOR2_X2 U7733 ( .A(rd_3[2]), .B(\hazard_detect/eq_83/A[2] ), .ZN(n6289) );
  XNOR2_X2 U7734 ( .A(rd_3[4]), .B(\hazard_detect/eq_83/A[4] ), .ZN(n6288) );
  XNOR2_X2 U7735 ( .A(rd_3[1]), .B(\hazard_detect/eq_83/A[1] ), .ZN(n6293) );
  XNOR2_X2 U7736 ( .A(n6291), .B(n2856), .ZN(n6292) );
  NAND2_X2 U7737 ( .A1(n6293), .A2(n6292), .ZN(n6295) );
  INV_X4 U7738 ( .A(n6300), .ZN(n7362) );
  INV_X4 U7739 ( .A(n6301), .ZN(n7361) );
  NOR2_X4 U7740 ( .A1(n7362), .A2(n7361), .ZN(n6305) );
  NOR2_X4 U7741 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  NAND2_X2 U7742 ( .A1(n6305), .A2(n6304), .ZN(n6307) );
  INV_X4 U7743 ( .A(n7884), .ZN(n6306) );
  AOI211_X2 U7744 ( .C1(n7711), .C2(n6307), .A(n6306), .B(n3119), .ZN(n6320)
         );
  INV_X4 U7745 ( .A(n7628), .ZN(n6308) );
  INV_X4 U7746 ( .A(n6309), .ZN(n6310) );
  INV_X4 U7747 ( .A(n6315), .ZN(n6316) );
  OAI211_X2 U7748 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n6317), .ZN(
        \id_ex/N37 ) );
  INV_X4 U7749 ( .A(n6322), .ZN(n7363) );
  INV_X4 U7750 ( .A(n6323), .ZN(n7364) );
  INV_X4 U7751 ( .A(n6324), .ZN(n7365) );
  INV_X4 U7752 ( .A(n6325), .ZN(n7366) );
  INV_X4 U7753 ( .A(n6326), .ZN(n7367) );
  INV_X4 U7754 ( .A(n6327), .ZN(n7368) );
  INV_X4 U7755 ( .A(n6328), .ZN(n7373) );
  INV_X4 U7756 ( .A(n6329), .ZN(n7374) );
  INV_X4 U7757 ( .A(n6330), .ZN(n7375) );
  INV_X4 U7758 ( .A(n6331), .ZN(n7359) );
  INV_X4 U7759 ( .A(n6332), .ZN(n7360) );
  NAND4_X2 U7760 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(n6367)
         );
  NAND4_X2 U7761 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6366)
         );
  NAND4_X2 U7762 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6365)
         );
  NAND4_X2 U7763 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n6364)
         );
  NOR4_X2 U7764 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .ZN(
        \ex_mem/N232 ) );
  MUX2_X2 U7765 ( .A(net224853), .B(n7182), .S(net221494), .Z(n6368) );
  NAND2_X2 U7766 ( .A1(n6368), .A2(n2838), .ZN(n6371) );
  INV_X4 U7767 ( .A(net221492), .ZN(net221489) );
  INV_X4 U7768 ( .A(n6384), .ZN(n6389) );
  MUX2_X2 U7769 ( .A(net224853), .B(n3913), .S(n6867), .Z(n6383) );
  NAND2_X2 U7770 ( .A1(n6383), .A2(n2838), .ZN(n6388) );
  NAND2_X2 U7771 ( .A1(n6384), .A2(net224843), .ZN(n6385) );
  NAND2_X2 U7772 ( .A1(n6394), .A2(n6393), .ZN(n6410) );
  INV_X4 U7773 ( .A(n6880), .ZN(n6407) );
  NOR2_X4 U7774 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  OAI21_X4 U7775 ( .B1(n3868), .B2(n6410), .A(n6409), .ZN(n6412) );
  INV_X4 U7776 ( .A(net220890), .ZN(net220865) );
  INV_X4 U7777 ( .A(n6416), .ZN(n6420) );
  INV_X4 U7778 ( .A(n6417), .ZN(n6418) );
  NAND4_X2 U7779 ( .A1(n3271), .A2(net230730), .A3(net221416), .A4(n6418), 
        .ZN(n6419) );
  AOI22_X2 U7780 ( .A1(n7358), .A2(n6422), .B1(n3953), .B2(n6859), .ZN(n6482)
         );
  NAND3_X2 U7781 ( .A1(n6427), .A2(n7936), .A3(n6426), .ZN(n6428) );
  INV_X4 U7782 ( .A(n6429), .ZN(n7210) );
  NAND3_X2 U7783 ( .A1(n3587), .A2(n7198), .A3(n7210), .ZN(n6435) );
  NAND2_X2 U7784 ( .A1(n6444), .A2(n6443), .ZN(n6456) );
  NAND3_X2 U7785 ( .A1(n6445), .A2(n3947), .A3(n3649), .ZN(n6446) );
  NOR2_X4 U7786 ( .A1(n6447), .A2(n6446), .ZN(n6454) );
  NOR2_X4 U7787 ( .A1(n6449), .A2(n6448), .ZN(n6453) );
  OAI21_X4 U7788 ( .B1(n6451), .B2(n3877), .A(n7242), .ZN(n6452) );
  NAND4_X2 U7789 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n7244), .ZN(n6455)
         );
  INV_X4 U7790 ( .A(n7222), .ZN(n6477) );
  INV_X4 U7792 ( .A(n6469), .ZN(n6472) );
  NAND2_X2 U7793 ( .A1(n6470), .A2(n3948), .ZN(n6471) );
  NAND2_X2 U7794 ( .A1(n6661), .A2(n6478), .ZN(n6480) );
  AOI22_X2 U7795 ( .A1(n7944), .A2(n3921), .B1(n7127), .B2(n6804), .ZN(n6481)
         );
  NAND4_X2 U7796 ( .A1(n6481), .A2(n6484), .A3(n6482), .A4(n6483), .ZN(
        \ex_mem/N226 ) );
  INV_X4 U7797 ( .A(n6512), .ZN(n7357) );
  NOR2_X4 U7798 ( .A1(n6696), .A2(n2701), .ZN(n6511) );
  INV_X4 U7799 ( .A(n6680), .ZN(n6593) );
  INV_X4 U7800 ( .A(n6826), .ZN(n6490) );
  NAND2_X2 U7801 ( .A1(n6710), .A2(n6677), .ZN(n6492) );
  AOI21_X4 U7802 ( .B1(n6493), .B2(n6492), .A(n6491), .ZN(n6494) );
  XNOR2_X2 U7803 ( .A(n6494), .B(n6552), .ZN(n7306) );
  INV_X4 U7804 ( .A(n6495), .ZN(n6496) );
  NOR2_X4 U7805 ( .A1(n6496), .A2(n7205), .ZN(n6499) );
  NOR2_X4 U7806 ( .A1(n6609), .A2(n3914), .ZN(n6498) );
  MUX2_X2 U7808 ( .A(n2902), .B(n6500), .S(net224733), .Z(n6501) );
  INV_X4 U7809 ( .A(n6501), .ZN(n6505) );
  MUX2_X2 U7810 ( .A(net224853), .B(n7182), .S(n6504), .Z(n6506) );
  NAND3_X2 U7811 ( .A1(n6520), .A2(n6519), .A3(n6518), .ZN(\ex_mem/N206 ) );
  NAND2_X2 U7812 ( .A1(n7127), .A2(n6521), .ZN(n6544) );
  MUX2_X2 U7813 ( .A(net224853), .B(n3913), .S(n6522), .Z(n6523) );
  AOI21_X4 U7814 ( .B1(n6529), .B2(n6528), .A(n6527), .ZN(n6531) );
  NAND2_X2 U7815 ( .A1(n7358), .A2(n6533), .ZN(n6534) );
  NAND2_X2 U7816 ( .A1(n7918), .A2(n3953), .ZN(n6542) );
  AOI22_X2 U7817 ( .A1(n7123), .A2(n6545), .B1(n3921), .B2(n6540), .ZN(n6541)
         );
  NAND4_X2 U7818 ( .A1(n6542), .A2(n6541), .A3(n6543), .A4(n6544), .ZN(
        \ex_mem/N209 ) );
  INV_X4 U7819 ( .A(n6545), .ZN(n6547) );
  OAI22_X2 U7820 ( .A1(n6547), .A2(n3954), .B1(n6546), .B2(n2701), .ZN(n6576)
         );
  NOR2_X4 U7821 ( .A1(n6550), .A2(n6701), .ZN(n6555) );
  INV_X4 U7822 ( .A(n6699), .ZN(n6551) );
  AOI211_X4 U7823 ( .C1(n6555), .C2(n6554), .A(n6553), .B(n2912), .ZN(n6561)
         );
  XNOR2_X2 U7824 ( .A(n6563), .B(n6562), .ZN(n7282) );
  MUX2_X2 U7825 ( .A(net224843), .B(n7151), .S(n6568), .Z(n6564) );
  NOR2_X2 U7826 ( .A1(n6576), .A2(n6575), .ZN(n6578) );
  MUX2_X2 U7827 ( .A(n2903), .B(n3160), .S(net224733), .Z(n6584) );
  MUX2_X2 U7828 ( .A(net224843), .B(n7151), .S(n6583), .Z(n6585) );
  INV_X4 U7829 ( .A(n6705), .ZN(n6587) );
  NAND3_X2 U7830 ( .A1(n6590), .A2(n7296), .A3(n6589), .ZN(n6597) );
  INV_X4 U7831 ( .A(n6600), .ZN(n6601) );
  NOR2_X4 U7832 ( .A1(n6601), .A2(n7205), .ZN(n6605) );
  NOR2_X4 U7833 ( .A1(n3914), .A2(n6668), .ZN(n6604) );
  NOR3_X4 U7834 ( .A1(n6605), .A2(n6603), .A3(n6604), .ZN(n7098) );
  OAI22_X2 U7835 ( .A1(n6607), .A2(n6672), .B1(n2703), .B2(n6606), .ZN(n6613)
         );
  NOR2_X4 U7836 ( .A1(n6609), .A2(n7205), .ZN(n6612) );
  MUX2_X2 U7837 ( .A(net224853), .B(n7182), .S(n3209), .Z(n6630) );
  NAND2_X2 U7838 ( .A1(n6630), .A2(n2838), .ZN(n6638) );
  NAND2_X2 U7839 ( .A1(n7358), .A2(n6632), .ZN(n6633) );
  INV_X4 U7840 ( .A(n6641), .ZN(n6642) );
  INV_X4 U7841 ( .A(n7205), .ZN(n6663) );
  AOI22_X2 U7842 ( .A1(n6663), .A2(n6662), .B1(n6660), .B2(n6661), .ZN(n6664)
         );
  INV_X4 U7843 ( .A(n7040), .ZN(n7000) );
  NOR3_X4 U7844 ( .A1(n6675), .A2(n6674), .A3(n6673), .ZN(n7026) );
  NAND2_X2 U7845 ( .A1(n6677), .A2(n3745), .ZN(n6731) );
  NAND3_X2 U7846 ( .A1(n6679), .A2(n2599), .A3(n6677), .ZN(n6732) );
  INV_X4 U7847 ( .A(n6682), .ZN(n7305) );
  MUX2_X2 U7848 ( .A(net224853), .B(n3913), .S(n6683), .Z(n6684) );
  NAND2_X2 U7849 ( .A1(n7358), .A2(n6686), .ZN(n6687) );
  OAI221_X2 U7850 ( .B1(n7071), .B2(n3954), .C1(n7000), .C2(n3923), .A(n6695), 
        .ZN(\ex_mem/N203 ) );
  AOI21_X4 U7851 ( .B1(n6711), .B2(n6703), .A(n2912), .ZN(n6713) );
  NAND3_X2 U7852 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6712) );
  MUX2_X2 U7853 ( .A(net224843), .B(n7151), .S(n2759), .Z(n6716) );
  NOR2_X2 U7854 ( .A1(n6727), .A2(n6726), .ZN(n6730) );
  MUX2_X2 U7855 ( .A(net224843), .B(n7151), .S(n6739), .Z(n6734) );
  OAI221_X2 U7856 ( .B1(n3274), .B2(n3923), .C1(n7000), .C2(n3954), .A(n6747), 
        .ZN(\ex_mem/N202 ) );
  INV_X4 U7857 ( .A(n6799), .ZN(n6752) );
  MUX2_X2 U7858 ( .A(net224853), .B(n7182), .S(n3773), .Z(n6759) );
  OAI21_X2 U7859 ( .B1(n6766), .B2(n3918), .A(n6765), .ZN(n6767) );
  NAND2_X2 U7860 ( .A1(n6769), .A2(n6768), .ZN(\ex_mem/N198 ) );
  MUX2_X2 U7861 ( .A(net224853), .B(n3913), .S(n7230), .Z(n6771) );
  INV_X4 U7862 ( .A(n6773), .ZN(n6774) );
  AOI22_X2 U7863 ( .A1(n7358), .A2(n6783), .B1(n7127), .B2(n6859), .ZN(n6785)
         );
  AOI22_X2 U7864 ( .A1(n7944), .A2(n7123), .B1(n3953), .B2(n6804), .ZN(n6784)
         );
  NAND4_X2 U7865 ( .A1(n6784), .A2(n6786), .A3(n6785), .A4(n6787), .ZN(
        \ex_mem/N196 ) );
  MUX2_X2 U7866 ( .A(net224853), .B(n7182), .S(n6788), .Z(n6789) );
  NAND2_X2 U7867 ( .A1(n6789), .A2(n2838), .ZN(n6797) );
  NAND2_X2 U7868 ( .A1(n7358), .A2(n6791), .ZN(n6792) );
  NAND2_X2 U7869 ( .A1(n3951), .A2(n2794), .ZN(n6807) );
  AOI22_X2 U7870 ( .A1(n7127), .A2(n6802), .B1(n3921), .B2(n6801), .ZN(n6806)
         );
  NAND4_X2 U7871 ( .A1(n6805), .A2(n6807), .A3(n6806), .A4(n6808), .ZN(
        \ex_mem/N197 ) );
  MUX2_X2 U7872 ( .A(net224853), .B(n3913), .S(n6810), .Z(n6813) );
  NAND2_X2 U7873 ( .A1(n7358), .A2(n6815), .ZN(n6816) );
  INV_X4 U7874 ( .A(n6822), .ZN(n6828) );
  XNOR2_X2 U7875 ( .A(n6830), .B(n3683), .ZN(n7302) );
  OAI221_X2 U7876 ( .B1(n7104), .B2(n3954), .C1(n7103), .C2(n3923), .A(n6834), 
        .ZN(\ex_mem/N205 ) );
  NOR2_X4 U7877 ( .A1(n6836), .A2(n3918), .ZN(n6850) );
  MUX2_X2 U7878 ( .A(net224853), .B(n7182), .S(n6840), .Z(n6841) );
  NOR4_X2 U7879 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6857)
         );
  NAND2_X2 U7880 ( .A1(n3921), .A2(n6851), .ZN(n6856) );
  NAND4_X2 U7881 ( .A1(n6855), .A2(n6854), .A3(n6856), .A4(n6857), .ZN(
        \ex_mem/N199 ) );
  AOI22_X2 U7882 ( .A1(net224855), .A2(n3255), .B1(n7127), .B2(n6858), .ZN(
        n6972) );
  NAND2_X2 U7883 ( .A1(n3924), .A2(n6859), .ZN(n6860) );
  INV_X4 U7884 ( .A(n6860), .ZN(n6864) );
  OAI22_X2 U7885 ( .A1(n6264), .A2(n2840), .B1(n7193), .B2(n3954), .ZN(n6863)
         );
  XNOR2_X2 U7887 ( .A(n6865), .B(net224859), .ZN(n6866) );
  INV_X4 U7889 ( .A(net220888), .ZN(net220838) );
  XNOR2_X2 U7890 ( .A(net220305), .B(net224861), .ZN(n6921) );
  INV_X4 U7891 ( .A(n6921), .ZN(n6910) );
  NAND2_X2 U7893 ( .A1(n6887), .A2(n6926), .ZN(n6908) );
  AOI21_X4 U7894 ( .B1(n3496), .B2(n6902), .A(n6889), .ZN(n6894) );
  NAND3_X2 U7895 ( .A1(n6891), .A2(n6892), .A3(n6902), .ZN(n6893) );
  OAI21_X4 U7896 ( .B1(n6894), .B2(n6900), .A(n6893), .ZN(n6898) );
  NAND3_X2 U7897 ( .A1(n6901), .A2(n3639), .A3(n3622), .ZN(n6903) );
  NAND3_X2 U7898 ( .A1(n6917), .A2(n6914), .A3(n3254), .ZN(n6907) );
  NOR3_X4 U7899 ( .A1(n6919), .A2(n6920), .A3(net220838), .ZN(n6922) );
  OAI21_X4 U7900 ( .B1(n6925), .B2(n6924), .A(n6923), .ZN(n7339) );
  NOR3_X4 U7901 ( .A1(n6929), .A2(n6928), .A3(n6927), .ZN(n6930) );
  NAND2_X2 U7902 ( .A1(n7176), .A2(n3862), .ZN(n7225) );
  NOR2_X4 U7903 ( .A1(n6934), .A2(n7244), .ZN(n6938) );
  OAI21_X4 U7904 ( .B1(n6938), .B2(n6937), .A(n7176), .ZN(n7228) );
  NOR2_X4 U7905 ( .A1(n6942), .A2(n7201), .ZN(n6963) );
  NAND2_X2 U7906 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  OAI21_X4 U7907 ( .B1(n6962), .B2(n6963), .A(n3955), .ZN(n7232) );
  AOI22_X2 U7908 ( .A1(n3921), .A2(n6968), .B1(n7151), .B2(n6967), .ZN(n6969)
         );
  NAND4_X2 U7909 ( .A1(n6972), .A2(n6969), .A3(n6970), .A4(n6971), .ZN(
        \ex_mem/N227 ) );
  MUX2_X2 U7910 ( .A(net224853), .B(n3913), .S(net220780), .Z(n6973) );
  NAND2_X2 U7911 ( .A1(n7358), .A2(n6974), .ZN(n6975) );
  NOR2_X4 U7912 ( .A1(n7026), .A2(n3923), .ZN(n6997) );
  NOR2_X4 U7913 ( .A1(n7057), .A2(n3482), .ZN(n7139) );
  NAND3_X2 U7914 ( .A1(n6982), .A2(n6981), .A3(n7055), .ZN(n6995) );
  OAI221_X2 U7915 ( .B1(n3274), .B2(n2701), .C1(n7000), .C2(n3918), .A(n6999), 
        .ZN(\ex_mem/N221 ) );
  NAND2_X2 U7916 ( .A1(net220882), .A2(n7002), .ZN(n7003) );
  INV_X4 U7917 ( .A(n7004), .ZN(n7005) );
  INV_X4 U7918 ( .A(n7008), .ZN(n7085) );
  NAND2_X2 U7919 ( .A1(n7085), .A2(n7009), .ZN(n7011) );
  NAND2_X2 U7920 ( .A1(n7011), .A2(n7010), .ZN(n7012) );
  INV_X4 U7921 ( .A(n7018), .ZN(n7333) );
  INV_X4 U7922 ( .A(n7024), .ZN(n7332) );
  INV_X4 U7924 ( .A(n7025), .ZN(n7279) );
  OAI22_X2 U7925 ( .A1(n7279), .A2(n3950), .B1(n7026), .B2(n3954), .ZN(n7038)
         );
  MUX2_X2 U7926 ( .A(net224853), .B(n7182), .S(n7027), .Z(n7028) );
  NAND2_X2 U7927 ( .A1(n3921), .A2(n7040), .ZN(n7041) );
  NAND3_X2 U7928 ( .A1(n7043), .A2(n7042), .A3(n7041), .ZN(\ex_mem/N220 ) );
  MUX2_X2 U7929 ( .A(net224853), .B(n3913), .S(n7044), .Z(n7045) );
  NAND2_X2 U7930 ( .A1(n7358), .A2(n7046), .ZN(n7047) );
  OAI221_X2 U7931 ( .B1(n7071), .B2(n2701), .C1(n7103), .C2(n3918), .A(n7070), 
        .ZN(\ex_mem/N219 ) );
  MUX2_X2 U7932 ( .A(net224853), .B(n7182), .S(net220656), .Z(n7072) );
  NAND3_X2 U7933 ( .A1(n7090), .A2(n7087), .A3(n7088), .ZN(n7093) );
  NAND2_X2 U7934 ( .A1(n7090), .A2(n7091), .ZN(n7092) );
  OAI21_X4 U7935 ( .B1(n7096), .B2(n7095), .A(n7094), .ZN(n7097) );
  OAI221_X2 U7936 ( .B1(n7104), .B2(n3918), .C1(n7103), .C2(n2701), .A(n7102), 
        .ZN(\ex_mem/N218 ) );
  MUX2_X2 U7937 ( .A(net224843), .B(n7151), .S(n7108), .Z(n7105) );
  NAND2_X2 U7938 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  NAND4_X2 U7939 ( .A1(n7130), .A2(n7131), .A3(n7132), .A4(n7129), .ZN(
        \ex_mem/N217 ) );
  NAND2_X2 U7941 ( .A1(n3923), .A2(n3918), .ZN(n7161) );
  INV_X4 U7942 ( .A(n7136), .ZN(n7137) );
  NAND2_X2 U7943 ( .A1(n7147), .A2(n7146), .ZN(n7304) );
  MUX2_X2 U7944 ( .A(net224843), .B(n7151), .S(n7150), .Z(n7152) );
  AOI211_X4 U7945 ( .C1(n7160), .C2(n7161), .A(n7158), .B(n7159), .ZN(n7162)
         );
  NAND3_X2 U7946 ( .A1(n7164), .A2(n7162), .A3(n7163), .ZN(\ex_mem/N212 ) );
  NAND2_X2 U7947 ( .A1(setInv_2), .A2(net220307), .ZN(n7165) );
  XNOR2_X2 U7948 ( .A(setInv_2), .B(net220310), .ZN(n7166) );
  INV_X4 U7949 ( .A(net220537), .ZN(net220535) );
  INV_X4 U7950 ( .A(n7170), .ZN(n7174) );
  NAND2_X2 U7951 ( .A1(n7176), .A2(n3953), .ZN(n7267) );
  INV_X4 U7952 ( .A(n7290), .ZN(n7189) );
  INV_X4 U7953 ( .A(n7178), .ZN(n7180) );
  MUX2_X2 U7954 ( .A(net224851), .B(n3913), .S(n7181), .Z(n7185) );
  OAI21_X4 U7955 ( .B1(n7189), .B2(n2706), .A(n7188), .ZN(n7260) );
  NAND2_X2 U7956 ( .A1(n7358), .A2(n7190), .ZN(n7191) );
  OAI21_X4 U7957 ( .B1(n7193), .B2(n3918), .A(n7191), .ZN(n7259) );
  INV_X4 U7958 ( .A(n7199), .ZN(n7208) );
  NOR2_X4 U7959 ( .A1(n7200), .A2(n7208), .ZN(n7211) );
  AND2_X2 U7960 ( .A1(n7202), .A2(n7201), .ZN(n7204) );
  NAND2_X2 U7961 ( .A1(n7204), .A2(n7203), .ZN(n7207) );
  OAI21_X4 U7962 ( .B1(n7208), .B2(n7207), .A(n7206), .ZN(n7209) );
  AOI21_X4 U7963 ( .B1(n7211), .B2(n7210), .A(n7209), .ZN(n7215) );
  NOR2_X4 U7964 ( .A1(n7252), .A2(n3088), .ZN(n7214) );
  NOR3_X4 U7965 ( .A1(n7216), .A2(n7215), .A3(n7214), .ZN(n7238) );
  INV_X4 U7966 ( .A(n7221), .ZN(n7223) );
  NOR2_X4 U7967 ( .A1(n7223), .A2(n7222), .ZN(n7236) );
  INV_X4 U7968 ( .A(n7228), .ZN(n7229) );
  NOR3_X4 U7969 ( .A1(n7229), .A2(n7231), .A3(n7230), .ZN(n7233) );
  OAI21_X4 U7970 ( .B1(n7235), .B2(n7236), .A(n7234), .ZN(n7271) );
  NAND3_X2 U7971 ( .A1(n7258), .A2(n7257), .A3(n7196), .ZN(n7265) );
  INV_X4 U7972 ( .A(n7259), .ZN(n7263) );
  NAND2_X2 U7973 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  OAI21_X4 U7974 ( .B1(n7268), .B2(n7267), .A(n7266), .ZN(n7269) );
  AOI21_X4 U7975 ( .B1(n7270), .B2(n3953), .A(n7269), .ZN(n7272) );
  NAND2_X2 U7976 ( .A1(n3567), .A2(n8012), .ZN(n7278) );
  NAND3_X2 U7977 ( .A1(n7279), .A2(n3250), .A3(n7324), .ZN(n7281) );
  NOR3_X4 U7978 ( .A1(n7281), .A2(n7280), .A3(n7318), .ZN(n7315) );
  NOR3_X4 U7979 ( .A1(n7286), .A2(n7284), .A3(n7285), .ZN(n7314) );
  NAND3_X2 U7980 ( .A1(n7294), .A2(n7293), .A3(n7292), .ZN(n7299) );
  NOR3_X4 U7981 ( .A1(n7309), .A2(n7308), .A3(n7307), .ZN(n7313) );
  AOI21_X4 U7982 ( .B1(n7316), .B2(n7315), .A(n7317), .ZN(n7322) );
  NOR2_X4 U7983 ( .A1(n7320), .A2(n7319), .ZN(n7321) );
  NOR3_X4 U7984 ( .A1(n3721), .A2(n7322), .A3(n7321), .ZN(net220285) );
  NAND3_X2 U7985 ( .A1(n7325), .A2(n7323), .A3(n7324), .ZN(n7329) );
  NOR2_X4 U7986 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  NOR2_X4 U7987 ( .A1(n7330), .A2(n7336), .ZN(net220294) );
  NOR2_X4 U7988 ( .A1(n7337), .A2(n7336), .ZN(net220295) );
  INV_X4 U7989 ( .A(n7338), .ZN(n7340) );
  NOR2_X4 U7990 ( .A1(n7340), .A2(n7339), .ZN(n7344) );
  INV_X4 U7991 ( .A(n7345), .ZN(n7347) );
  NAND2_X2 U7992 ( .A1(n7347), .A2(n7346), .ZN(regWrData[18]) );
  INV_X4 U7993 ( .A(n7351), .ZN(n7353) );
  NAND2_X2 U7994 ( .A1(n7353), .A2(n7352), .ZN(regWrData[25]) );
  OAI222_X2 U7995 ( .A1(n7381), .A2(net224765), .B1(net224755), .B2(n2737), 
        .C1(net36084), .C2(n7541), .ZN(memWrData[16]) );
  OAI222_X2 U7996 ( .A1(n7405), .A2(net224767), .B1(net224755), .B2(n2726), 
        .C1(net36084), .C2(n7411), .ZN(memWrData[17]) );
  OAI222_X2 U7997 ( .A1(n7406), .A2(net224765), .B1(net224755), .B2(n2734), 
        .C1(net36084), .C2(n7412), .ZN(memWrData[18]) );
  OAI222_X2 U7998 ( .A1(n7407), .A2(net224767), .B1(net224755), .B2(n2728), 
        .C1(net36084), .C2(n7415), .ZN(memWrData[20]) );
  OAI222_X2 U7999 ( .A1(n7383), .A2(net224767), .B1(net224755), .B2(n2732), 
        .C1(net36084), .C2(n7539), .ZN(memWrData[22]) );
  OAI222_X2 U8000 ( .A1(n7384), .A2(net224767), .B1(net224755), .B2(n2729), 
        .C1(net36084), .C2(n7538), .ZN(memWrData[23]) );
  OAI222_X2 U8001 ( .A1(n7385), .A2(net224767), .B1(net224755), .B2(n2730), 
        .C1(net36084), .C2(n7537), .ZN(memWrData[24]) );
  OAI222_X2 U8002 ( .A1(n7386), .A2(net224767), .B1(net224755), .B2(n2733), 
        .C1(net224773), .C2(n7536), .ZN(memWrData[25]) );
  OAI222_X2 U8004 ( .A1(n7409), .A2(net224765), .B1(net224759), .B2(n2784), 
        .C1(net224773), .C2(n7422), .ZN(memWrData[27]) );
  OAI222_X2 U8005 ( .A1(n7410), .A2(net224765), .B1(net224755), .B2(n2787), 
        .C1(net224773), .C2(n7424), .ZN(memWrData[28]) );
  OAI222_X2 U8006 ( .A1(n7395), .A2(net224765), .B1(net224759), .B2(n2791), 
        .C1(net224773), .C2(n7526), .ZN(memWrData[29]) );
  OAI222_X2 U8007 ( .A1(n7401), .A2(net224765), .B1(net224755), .B2(n2781), 
        .C1(net224773), .C2(n7500), .ZN(memWrData[30]) );
  OAI222_X2 U8008 ( .A1(n7387), .A2(net224765), .B1(net224759), .B2(n2731), 
        .C1(net224773), .C2(n7535), .ZN(memWrData[31]) );
  MUX2_X1 U8009 ( .A(rd_3[4]), .B(rd[4]), .S(net224717), .Z(n7752) );
  MUX2_X1 U8010 ( .A(rd_3[3]), .B(rd[3]), .S(net224717), .Z(n7753) );
  MUX2_X1 U8011 ( .A(rd_3[2]), .B(rd[2]), .S(net224717), .Z(n7754) );
  MUX2_X1 U8012 ( .A(rd_3[1]), .B(rd[1]), .S(net224717), .Z(n7755) );
  MUX2_X1 U8013 ( .A(rd_3[0]), .B(rd[0]), .S(net224717), .Z(n7756) );
  INV_X1 U8014 ( .A(n7580), .ZN(n7758) );
  MUX2_X1 U8015 ( .A(n7533), .B(n7569), .S(net224719), .Z(n7580) );
  INV_X1 U8016 ( .A(n7581), .ZN(n7759) );
  MUX2_X1 U8017 ( .A(n7525), .B(n7561), .S(net224719), .Z(n7581) );
  INV_X1 U8018 ( .A(n7582), .ZN(n7760) );
  MUX2_X1 U8019 ( .A(n7535), .B(n7571), .S(net224719), .Z(n7582) );
  INV_X1 U8020 ( .A(n7583), .ZN(n7761) );
  MUX2_X1 U8021 ( .A(n7500), .B(n7557), .S(net224719), .Z(n7583) );
  INV_X1 U8022 ( .A(n7584), .ZN(n7762) );
  MUX2_X1 U8023 ( .A(n7526), .B(n7562), .S(net224719), .Z(n7584) );
  INV_X1 U8024 ( .A(n7585), .ZN(n7763) );
  MUX2_X1 U8025 ( .A(n7424), .B(n7551), .S(net224719), .Z(n7585) );
  INV_X1 U8026 ( .A(n7586), .ZN(n7764) );
  MUX2_X1 U8027 ( .A(n7422), .B(n7550), .S(net224719), .Z(n7586) );
  INV_X1 U8028 ( .A(n7587), .ZN(n7765) );
  MUX2_X1 U8029 ( .A(n7421), .B(n7549), .S(net224719), .Z(n7587) );
  INV_X1 U8030 ( .A(n7588), .ZN(n7766) );
  MUX2_X1 U8031 ( .A(n7536), .B(n7572), .S(net224719), .Z(n7588) );
  INV_X1 U8032 ( .A(n7589), .ZN(n7767) );
  MUX2_X1 U8033 ( .A(n7537), .B(n7573), .S(net224719), .Z(n7589) );
  INV_X1 U8034 ( .A(n7590), .ZN(n7768) );
  MUX2_X1 U8035 ( .A(n7538), .B(n7574), .S(net224719), .Z(n7590) );
  INV_X1 U8036 ( .A(n7591), .ZN(n7769) );
  MUX2_X1 U8037 ( .A(n7539), .B(n7575), .S(net224719), .Z(n7591) );
  INV_X1 U8038 ( .A(n7592), .ZN(n7770) );
  MUX2_X1 U8039 ( .A(n7540), .B(n7576), .S(net224719), .Z(n7592) );
  INV_X1 U8040 ( .A(n7593), .ZN(n7771) );
  MUX2_X1 U8041 ( .A(n7415), .B(n7546), .S(net224719), .Z(n7593) );
  INV_X1 U8042 ( .A(net35483), .ZN(net33021) );
  INV_X1 U8043 ( .A(n7594), .ZN(n7772) );
  MUX2_X1 U8044 ( .A(n7412), .B(n7544), .S(net224719), .Z(n7594) );
  INV_X1 U8045 ( .A(n7595), .ZN(n7773) );
  MUX2_X1 U8046 ( .A(n7411), .B(n7543), .S(net224719), .Z(n7595) );
  INV_X1 U8047 ( .A(n7596), .ZN(n7774) );
  MUX2_X1 U8048 ( .A(n7541), .B(n7577), .S(net224719), .Z(n7596) );
  INV_X1 U8049 ( .A(n7597), .ZN(n7775) );
  MUX2_X1 U8050 ( .A(n7414), .B(n7545), .S(net224721), .Z(n7597) );
  INV_X1 U8051 ( .A(n7598), .ZN(n7776) );
  MUX2_X1 U8052 ( .A(n7417), .B(n7547), .S(net224721), .Z(n7598) );
  INV_X1 U8053 ( .A(n7599), .ZN(n7777) );
  MUX2_X1 U8054 ( .A(n7523), .B(n7559), .S(net224721), .Z(n7599) );
  INV_X1 U8055 ( .A(n7600), .ZN(n7778) );
  MUX2_X1 U8056 ( .A(n7524), .B(n7560), .S(net224721), .Z(n7600) );
  INV_X1 U8057 ( .A(n7601), .ZN(n7779) );
  MUX2_X1 U8058 ( .A(n7528), .B(n7564), .S(net224721), .Z(n7601) );
  INV_X1 U8059 ( .A(n7602), .ZN(n7780) );
  MUX2_X1 U8060 ( .A(n7522), .B(n7558), .S(net224721), .Z(n7602) );
  MUX2_X1 U8063 ( .A(memRdData[0]), .B(\wb/dsize_reg/z2 [0]), .S(net224721), 
        .Z(n2267) );
  MUX2_X1 U8064 ( .A(memRdData[1]), .B(\wb/dsize_reg/z2 [1]), .S(net224721), 
        .Z(n2266) );
  MUX2_X1 U8065 ( .A(memRdData[2]), .B(\wb/dsize_reg/z2 [2]), .S(net224721), 
        .Z(n2265) );
  MUX2_X1 U8066 ( .A(memRdData[3]), .B(\wb/dsize_reg/z2 [3]), .S(net224721), 
        .Z(n2264) );
  MUX2_X1 U8067 ( .A(memRdData[4]), .B(\wb/dsize_reg/z2 [4]), .S(net224721), 
        .Z(n2263) );
  MUX2_X1 U8068 ( .A(memRdData[5]), .B(\wb/dsize_reg/z2 [5]), .S(net224721), 
        .Z(n2262) );
  MUX2_X1 U8069 ( .A(memRdData[6]), .B(\wb/dsize_reg/z2 [6]), .S(net224721), 
        .Z(n2261) );
  MUX2_X1 U8070 ( .A(memRdData[7]), .B(\wb/dsize_reg/z2 [7]), .S(net224721), 
        .Z(n2260) );
  MUX2_X1 U8071 ( .A(memRdData[8]), .B(\wb/dsize_reg/z2 [8]), .S(net224721), 
        .Z(n2259) );
  MUX2_X1 U8072 ( .A(memRdData[9]), .B(\wb/dsize_reg/z2 [9]), .S(net224721), 
        .Z(n2258) );
  MUX2_X1 U8073 ( .A(memRdData[10]), .B(\wb/dsize_reg/z2 [10]), .S(net224721), 
        .Z(n2257) );
  MUX2_X1 U8074 ( .A(memRdData[11]), .B(\wb/dsize_reg/z2 [11]), .S(net224721), 
        .Z(n2256) );
  MUX2_X1 U8075 ( .A(memRdData[12]), .B(\wb/dsize_reg/z2 [12]), .S(net224723), 
        .Z(n2255) );
  MUX2_X1 U8076 ( .A(memRdData[13]), .B(\wb/dsize_reg/z2 [13]), .S(net224723), 
        .Z(n2254) );
  MUX2_X1 U8077 ( .A(memRdData[14]), .B(\wb/dsize_reg/z2 [14]), .S(net224723), 
        .Z(n2253) );
  MUX2_X1 U8078 ( .A(memRdData[15]), .B(\wb/dsize_reg/z2 [15]), .S(net224723), 
        .Z(n2252) );
  MUX2_X1 U8079 ( .A(memRdData[16]), .B(\wb/dsize_reg/z2 [16]), .S(net224723), 
        .Z(n2251) );
  MUX2_X1 U8080 ( .A(memRdData[17]), .B(\wb/dsize_reg/z2 [17]), .S(net224723), 
        .Z(n2250) );
  MUX2_X1 U8081 ( .A(memRdData[18]), .B(\wb/dsize_reg/z2 [18]), .S(net224723), 
        .Z(n2249) );
  MUX2_X1 U8082 ( .A(memRdData[19]), .B(\wb/dsize_reg/z2 [19]), .S(net224723), 
        .Z(n2248) );
  MUX2_X1 U8083 ( .A(memRdData[20]), .B(\wb/dsize_reg/z2 [20]), .S(net224723), 
        .Z(n2247) );
  MUX2_X1 U8084 ( .A(memRdData[21]), .B(\wb/dsize_reg/z2 [21]), .S(net224723), 
        .Z(n2246) );
  MUX2_X1 U8085 ( .A(memRdData[22]), .B(\wb/dsize_reg/z2 [22]), .S(net224723), 
        .Z(n2245) );
  MUX2_X1 U8086 ( .A(memRdData[23]), .B(\wb/dsize_reg/z2 [23]), .S(net224723), 
        .Z(n2244) );
  MUX2_X1 U8087 ( .A(memRdData[24]), .B(\wb/dsize_reg/z2 [24]), .S(net224723), 
        .Z(n2243) );
  MUX2_X1 U8088 ( .A(memRdData[25]), .B(\wb/dsize_reg/z2 [25]), .S(net224723), 
        .Z(n2242) );
  MUX2_X1 U8089 ( .A(memRdData[27]), .B(\wb/dsize_reg/z2 [27]), .S(net224723), 
        .Z(n2240) );
  MUX2_X1 U8090 ( .A(memRdData[28]), .B(\wb/dsize_reg/z2 [28]), .S(net224723), 
        .Z(n2239) );
  MUX2_X1 U8091 ( .A(memRdData[29]), .B(\wb/dsize_reg/z2 [29]), .S(net224725), 
        .Z(n2238) );
  MUX2_X1 U8092 ( .A(memRdData[30]), .B(\wb/dsize_reg/z2 [30]), .S(net224725), 
        .Z(n2237) );
  MUX2_X1 U8093 ( .A(memRdData[31]), .B(\wb/dsize_reg/z2 [31]), .S(net224725), 
        .Z(n2236) );
  INV_X1 U8094 ( .A(n7608), .ZN(n2235) );
  MUX2_X1 U8095 ( .A(n7542), .B(n7578), .S(net224725), .Z(n7608) );
  INV_X1 U8096 ( .A(n7609), .ZN(n2227) );
  MUX2_X1 U8097 ( .A(n7534), .B(n7570), .S(net224725), .Z(n7609) );
  INV_X1 U8098 ( .A(n7610), .ZN(n2225) );
  MUX2_X1 U8099 ( .A(n7532), .B(n7568), .S(net224725), .Z(n7610) );
  INV_X1 U8100 ( .A(n7611), .ZN(n2224) );
  MUX2_X1 U8101 ( .A(n7531), .B(n7567), .S(net224725), .Z(n7611) );
  INV_X1 U8102 ( .A(n7612), .ZN(n2223) );
  MUX2_X1 U8103 ( .A(n7530), .B(n7566), .S(net224725), .Z(n7612) );
  INV_X1 U8104 ( .A(n7613), .ZN(n2222) );
  MUX2_X1 U8105 ( .A(n7529), .B(n7565), .S(net224725), .Z(n7613) );
  INV_X1 U8106 ( .A(n7614), .ZN(n2220) );
  MUX2_X1 U8107 ( .A(n7527), .B(n7563), .S(net224725), .Z(n7614) );
  INV_X1 U8108 ( .A(n7616), .ZN(n1948) );
  MUX2_X1 U8109 ( .A(n7420), .B(n7548), .S(net224725), .Z(n7616) );
  OR2_X1 U8110 ( .A1(net224685), .A2(initPC[30]), .ZN(n1914) );
  NAND2_X1 U8111 ( .A1(initPC[30]), .A2(net224725), .ZN(n1913) );
  OR2_X1 U8112 ( .A1(net224685), .A2(initPC[29]), .ZN(n1912) );
  NAND2_X1 U8113 ( .A1(initPC[29]), .A2(net224725), .ZN(n1911) );
  OR2_X1 U8114 ( .A1(net224685), .A2(initPC[28]), .ZN(n1910) );
  NAND2_X1 U8115 ( .A1(initPC[28]), .A2(net224725), .ZN(n1909) );
  OR2_X1 U8116 ( .A1(net224685), .A2(initPC[27]), .ZN(n1908) );
  NAND2_X1 U8117 ( .A1(initPC[27]), .A2(net224725), .ZN(n1907) );
  OR2_X1 U8118 ( .A1(net224685), .A2(initPC[26]), .ZN(n1906) );
  NAND2_X1 U8119 ( .A1(initPC[26]), .A2(net224725), .ZN(n1905) );
  OR2_X1 U8120 ( .A1(net224645), .A2(initPC[25]), .ZN(n1904) );
  NAND2_X1 U8121 ( .A1(initPC[25]), .A2(net224725), .ZN(n1903) );
  OR2_X1 U8122 ( .A1(net224625), .A2(initPC[24]), .ZN(n1902) );
  NAND2_X1 U8123 ( .A1(initPC[24]), .A2(net224725), .ZN(n1901) );
  OR2_X1 U8124 ( .A1(net224663), .A2(initPC[23]), .ZN(n1900) );
  NAND2_X1 U8125 ( .A1(initPC[23]), .A2(net224725), .ZN(n1899) );
  OR2_X1 U8126 ( .A1(net224661), .A2(initPC[22]), .ZN(n1898) );
  NAND2_X1 U8127 ( .A1(initPC[22]), .A2(net224725), .ZN(n1897) );
  OR2_X1 U8128 ( .A1(net224673), .A2(initPC[21]), .ZN(n1896) );
  NAND2_X1 U8129 ( .A1(initPC[21]), .A2(net224727), .ZN(n1895) );
  OR2_X1 U8130 ( .A1(net224637), .A2(initPC[20]), .ZN(n1894) );
  NAND2_X1 U8131 ( .A1(initPC[20]), .A2(net224727), .ZN(n1893) );
  OR2_X1 U8132 ( .A1(net224621), .A2(initPC[19]), .ZN(n1892) );
  NAND2_X1 U8133 ( .A1(initPC[19]), .A2(net224727), .ZN(n1891) );
  OR2_X1 U8134 ( .A1(net224627), .A2(initPC[18]), .ZN(n1890) );
  NAND2_X1 U8135 ( .A1(initPC[18]), .A2(net224727), .ZN(n1889) );
  OR2_X1 U8136 ( .A1(net224629), .A2(initPC[17]), .ZN(n1888) );
  NAND2_X1 U8137 ( .A1(initPC[17]), .A2(net224727), .ZN(n1887) );
  OR2_X1 U8138 ( .A1(net224657), .A2(initPC[16]), .ZN(n1886) );
  NAND2_X1 U8139 ( .A1(initPC[16]), .A2(net224727), .ZN(n1885) );
  OR2_X1 U8140 ( .A1(net224623), .A2(initPC[15]), .ZN(n1884) );
  NAND2_X1 U8141 ( .A1(initPC[15]), .A2(net224727), .ZN(n1883) );
  OR2_X1 U8142 ( .A1(net224633), .A2(initPC[14]), .ZN(n1882) );
  NAND2_X1 U8143 ( .A1(initPC[14]), .A2(net224727), .ZN(n1881) );
  OR2_X1 U8144 ( .A1(net224669), .A2(initPC[13]), .ZN(n1880) );
  NAND2_X1 U8145 ( .A1(initPC[13]), .A2(net224727), .ZN(n1879) );
  OR2_X1 U8146 ( .A1(net224675), .A2(initPC[11]), .ZN(n1878) );
  NAND2_X1 U8147 ( .A1(initPC[11]), .A2(net224727), .ZN(n1877) );
  OR2_X1 U8148 ( .A1(net224631), .A2(initPC[10]), .ZN(n1876) );
  NAND2_X1 U8149 ( .A1(initPC[10]), .A2(net224727), .ZN(n1875) );
  OR2_X1 U8150 ( .A1(net224659), .A2(initPC[0]), .ZN(n1874) );
  NAND2_X1 U8151 ( .A1(initPC[0]), .A2(net224727), .ZN(n1873) );
  OR2_X1 U8152 ( .A1(net224653), .A2(initPC[1]), .ZN(n1872) );
  NAND2_X1 U8153 ( .A1(initPC[1]), .A2(net224727), .ZN(n1871) );
  OR2_X1 U8154 ( .A1(net224635), .A2(initPC[2]), .ZN(n1870) );
  NAND2_X1 U8155 ( .A1(initPC[2]), .A2(net224727), .ZN(n1869) );
  OR2_X1 U8156 ( .A1(net224631), .A2(initPC[3]), .ZN(n1868) );
  NAND2_X1 U8157 ( .A1(initPC[3]), .A2(net224727), .ZN(n1867) );
  OR2_X1 U8158 ( .A1(net224655), .A2(initPC[4]), .ZN(n1866) );
  NAND2_X1 U8159 ( .A1(initPC[4]), .A2(net224727), .ZN(n1865) );
  OR2_X1 U8160 ( .A1(net224613), .A2(initPC[6]), .ZN(n1864) );
  NAND2_X1 U8161 ( .A1(initPC[6]), .A2(net224727), .ZN(n1863) );
  OR2_X1 U8162 ( .A1(net224611), .A2(initPC[7]), .ZN(n1862) );
  NAND2_X1 U8163 ( .A1(initPC[7]), .A2(net224727), .ZN(n1861) );
  OR2_X1 U8164 ( .A1(net224613), .A2(initPC[8]), .ZN(n1860) );
  NAND2_X1 U8165 ( .A1(initPC[8]), .A2(net224727), .ZN(n1859) );
  OR2_X1 U8166 ( .A1(net224679), .A2(initPC[9]), .ZN(n1858) );
  NAND2_X1 U8167 ( .A1(initPC[9]), .A2(net224727), .ZN(n1857) );
  OR2_X1 U8168 ( .A1(net224611), .A2(initPC[12]), .ZN(n1856) );
  NAND2_X1 U8169 ( .A1(initPC[12]), .A2(net224727), .ZN(n1855) );
  OR2_X1 U8170 ( .A1(net224679), .A2(initPC[5]), .ZN(n1854) );
  NAND2_X1 U8171 ( .A1(initPC[5]), .A2(net224727), .ZN(n1853) );
  OR2_X1 U8172 ( .A1(net224679), .A2(initPC[31]), .ZN(n1852) );
  NAND2_X1 U8173 ( .A1(initPC[31]), .A2(net224727), .ZN(n1851) );
  OAI222_X1 U8174 ( .A1(n7533), .A2(net224773), .B1(n7389), .B2(net224767), 
        .C1(n2927), .C2(net224759), .ZN(memWrData[9]) );
  OAI222_X1 U8175 ( .A1(n7525), .A2(net224773), .B1(n7396), .B2(net224767), 
        .C1(n2949), .C2(net224759), .ZN(memWrData[8]) );
  OAI222_X1 U8176 ( .A1(n7527), .A2(net224773), .B1(n7380), .B2(net224767), 
        .C1(n2783), .C2(net224759), .ZN(memWrData[7]) );
  OAI222_X1 U8177 ( .A1(n7529), .A2(net224773), .B1(n7393), .B2(net224767), 
        .C1(n3010), .C2(net224759), .ZN(memWrData[6]) );
  OAI222_X1 U8178 ( .A1(n7420), .A2(net224773), .B1(n7402), .B2(net224767), 
        .C1(n2779), .C2(net224759), .ZN(memWrData[5]) );
  OAI222_X1 U8179 ( .A1(n7534), .A2(net224773), .B1(n7388), .B2(net224767), 
        .C1(n2777), .C2(net224759), .ZN(memWrData[4]) );
  OAI222_X1 U8180 ( .A1(n7530), .A2(net224773), .B1(n7392), .B2(net224765), 
        .C1(n3772), .C2(net224759), .ZN(memWrData[3]) );
  OAI222_X1 U8181 ( .A1(n7532), .A2(net224773), .B1(n7390), .B2(net224765), 
        .C1(n2780), .C2(net224759), .ZN(memWrData[2]) );
  OAI222_X1 U8182 ( .A1(n7531), .A2(net224773), .B1(n7391), .B2(net224765), 
        .C1(n2785), .C2(net224759), .ZN(memWrData[1]) );
  OAI222_X1 U8183 ( .A1(n7414), .A2(net224773), .B1(n7404), .B2(net224765), 
        .C1(n2967), .C2(net224759), .ZN(memWrData[15]) );
  OAI222_X1 U8184 ( .A1(n7417), .A2(net224773), .B1(n7403), .B2(net224765), 
        .C1(n2782), .C2(net224759), .ZN(memWrData[14]) );
  OAI222_X1 U8185 ( .A1(n7523), .A2(net224773), .B1(n7398), .B2(net224765), 
        .C1(n3078), .C2(net224759), .ZN(memWrData[13]) );
  OAI222_X1 U8186 ( .A1(n7524), .A2(net224773), .B1(n7397), .B2(net224765), 
        .C1(n2948), .C2(net224759), .ZN(memWrData[12]) );
  OAI222_X1 U8187 ( .A1(n7528), .A2(net224773), .B1(n7394), .B2(net224765), 
        .C1(n2947), .C2(net224759), .ZN(memWrData[11]) );
  OAI222_X1 U8188 ( .A1(n7522), .A2(net224773), .B1(n7399), .B2(net224765), 
        .C1(n2964), .C2(net224759), .ZN(memWrData[10]) );
  OAI222_X1 U8189 ( .A1(n7542), .A2(net36084), .B1(n7478), .B2(net224767), 
        .C1(n2727), .C2(net224755), .ZN(memWrData[0]) );
  NAND2_X1 U8190 ( .A1(n7469), .A2(n2723), .ZN(net36084) );
  NAND3_X1 U8191 ( .A1(instr_2[2]), .A2(instr_2[4]), .A3(instr_2[0]), .ZN(
        n7617) );
  NOR2_X1 U8192 ( .A1(instr_2[6]), .A2(instr_2[7]), .ZN(n7618) );
  NAND3_X1 U8193 ( .A1(n7484), .A2(n7483), .A3(n7485), .ZN(n7620) );
  NAND4_X1 U8194 ( .A1(n7482), .A2(n7481), .A3(n7621), .A4(n7480), .ZN(n7619)
         );
  NOR2_X1 U8195 ( .A1(instr_2[8]), .A2(instr_2[9]), .ZN(n7621) );
  NAND3_X1 U8196 ( .A1(n7490), .A2(n7489), .A3(n7491), .ZN(n7623) );
  NAND4_X1 U8197 ( .A1(n7488), .A2(n7487), .A3(n7624), .A4(n7486), .ZN(n7622)
         );
  NOR2_X1 U8198 ( .A1(instr_2[18]), .A2(instr_2[19]), .ZN(n7624) );
  XOR2_X1 U8199 ( .A(n2871), .B(rd_2[2]), .Z(n7627) );
  XOR2_X1 U8200 ( .A(n2899), .B(rd_2[3]), .Z(n7626) );
  XNOR2_X1 U8201 ( .A(rd_3[4]), .B(rd_2[4]), .ZN(n7625) );
  NOR2_X1 U8202 ( .A1(n7713), .A2(n2855), .ZN(n7628) );
  DFFR_X1 \if_id/instr_q_reg[20]  ( .D(n2159), .CK(clk), .RN(net224637), .Q(
        n2968), .QN(n7649) );
  DFFR_X1 \if_id/instr_q_reg[19]  ( .D(n2158), .CK(clk), .RN(net224673), .Q(
        n2954), .QN(n7648) );
  DFFR_X1 \if_id/instr_q_reg[18]  ( .D(n2157), .CK(clk), .RN(net224625), .Q(
        n2953), .QN(n7647) );
  DFFR_X1 \if_id/instr_q_reg[17]  ( .D(n2156), .CK(clk), .RN(net224663), .Q(
        n2952), .QN(n7646) );
  DFFR_X1 \if_id/instr_q_reg[16]  ( .D(n2155), .CK(clk), .RN(net224625), .Q(
        n2963), .QN(n7645) );
  DFFR_X1 \if_id/instr_q_reg[30]  ( .D(n2169), .CK(clk), .RN(net224625), .Q(
        n2858), .QN(n7713) );
  DFFR_X1 \if_id/instr_q_reg[5]  ( .D(n2144), .CK(clk), .RN(net224623), .Q(
        n2847), .QN(n7711) );
  DFFR_X1 \if_id/instr_q_reg[3]  ( .D(n2142), .CK(clk), .RN(net224623), .Q(
        n2761), .QN(net33230) );
  DFFR_X1 \if_id/instr_q_reg[1]  ( .D(n2140), .CK(clk), .RN(net224625), .Q(
        n2720), .QN(n7712) );
  DFFR_X1 \if_id/instr_q_reg[25]  ( .D(n2164), .CK(clk), .RN(net224625), .Q(
        rs1[4]), .QN(n2904) );
  DFFR_X1 \if_id/instr_q_reg[22]  ( .D(n2161), .CK(clk), .RN(net224621), .Q(
        rs1[1]), .QN(n2907) );
  DFFR_X1 \if_id/instr_q_reg[23]  ( .D(n2162), .CK(clk), .RN(net224625), .Q(
        rs1[2]), .QN(n2908) );
  DFFR_X1 \if_id/instr_q_reg[21]  ( .D(n2160), .CK(clk), .RN(net224625), .Q(
        rs1[0]), .QN(n2909) );
  DFFR_X1 \id_ex/busB_q_reg[31]  ( .D(n7813), .CK(clk), .RN(net224661), .Q(
        n2890), .QN(n7676) );
  DFFR_X1 \id_ex/busB_q_reg[27]  ( .D(n7817), .CK(clk), .RN(net224671), .Q(
        n2873), .QN(n7677) );
  DFFR_X1 \id_ex/busB_q_reg[26]  ( .D(n7818), .CK(clk), .RN(net224663), .Q(
        n2874), .QN(n7678) );
  DFFR_X1 \id_ex/busB_q_reg[25]  ( .D(n7819), .CK(clk), .RN(net224673), .Q(
        n2891), .QN(n7679) );
  DFFR_X1 \id_ex/busB_q_reg[22]  ( .D(n7822), .CK(clk), .RN(net224663), .Q(
        n2875), .QN(n7680) );
  DFFR_X1 \id_ex/busB_q_reg[21]  ( .D(n7823), .CK(clk), .RN(net224673), .Q(
        n2888), .QN(n7681) );
  DFFR_X1 \id_ex/busB_q_reg[20]  ( .D(n7824), .CK(clk), .RN(net224663), .Q(
        n2876), .QN(n7682) );
  DFFR_X1 \id_ex/busB_q_reg[19]  ( .D(n7825), .CK(clk), .RN(net224663), .Q(
        n2862), .QN(net33280) );
  DFFR_X1 \id_ex/busB_q_reg[18]  ( .D(n7826), .CK(clk), .RN(net224673), .Q(
        n2877), .QN(n7683) );
  DFFR_X1 \id_ex/busB_q_reg[16]  ( .D(n7828), .CK(clk), .RN(net224673), .Q(
        n2889), .QN(n7684) );
  DFFR_X1 \id_ex/busB_q_reg[0]  ( .D(n7844), .CK(clk), .RN(net224663), .Q(
        n2878), .QN(n7685) );
  DFFR_X1 \id_ex/busA_q_reg[30]  ( .D(n7782), .CK(clk), .RN(net224675), .Q(
        n2864), .QN(n7692) );
  DFFR_X1 \id_ex/busA_q_reg[28]  ( .D(n7784), .CK(clk), .RN(net224679), .Q(
        n2860), .QN(n7694) );
  DFFR_X1 \id_ex/busA_q_reg[27]  ( .D(n7785), .CK(clk), .RN(net224675), .Q(
        n2872), .QN(n7695) );
  DFFR_X1 \id_ex/busA_q_reg[26]  ( .D(n7786), .CK(clk), .RN(net224679), .Q(
        n2866), .QN(n7696) );
  DFFR_X1 \id_ex/busA_q_reg[24]  ( .D(n7788), .CK(clk), .RN(net224679), .Q(
        n2879), .QN(n7697) );
  DFFR_X1 \id_ex/busA_q_reg[17]  ( .D(n7795), .CK(clk), .RN(net224669), .Q(
        n2880), .QN(n7699) );
  DFFR_X1 \id_ex/busA_q_reg[16]  ( .D(n7796), .CK(clk), .RN(net224675), .Q(
        n2892), .QN(n7700) );
  DFFR_X1 \id_ex/busA_q_reg[15]  ( .D(n7797), .CK(clk), .RN(net224613), .Q(
        n2881), .QN(n7701) );
  DFFR_X1 \id_ex/busA_q_reg[14]  ( .D(n7798), .CK(clk), .RN(net224675), .Q(
        n2861), .QN(n7702) );
  DFFR_X1 \id_ex/busA_q_reg[13]  ( .D(n7799), .CK(clk), .RN(net224611), .Q(
        n2893), .QN(n7703) );
  DFFR_X1 \id_ex/busA_q_reg[12]  ( .D(n7800), .CK(clk), .RN(net224675), .Q(
        n3744) );
  DFFR_X1 \id_ex/busA_q_reg[11]  ( .D(n7801), .CK(clk), .RN(net224679), .Q(
        n2895), .QN(n7705) );
  DFFR_X1 \ex_mem/op0_q_reg  ( .D(\ex_mem/N237 ), .CK(clk), .RN(net224645), 
        .QN(n3281) );
  DFFR_X1 \ex_mem/imm32_q_reg[2]  ( .D(\ex_mem/N133 ), .CK(clk), .RN(net224641), .QN(n7438) );
  DFFR_X1 \ex_mem/busB_q_reg[11]  ( .D(\ex_mem/N110 ), .CK(clk), .RN(net224631), .QN(n7394) );
  DFFR_X1 \ex_mem/imm32_q_reg[5]  ( .D(\ex_mem/N136 ), .CK(clk), .RN(net224641), .Q(n3989), .QN(n7441) );
  DFFR_X1 \ex_mem/imm32_q_reg[0]  ( .D(\ex_mem/N131 ), .CK(clk), .RN(net224641), .Q(n4462) );
  DFFR_X1 \ex_mem/incPC_q_reg[30]  ( .D(\ex_mem/N65 ), .CK(clk), .RN(net224617), .Q(n2669), .QN(n7501) );
  DFFR_X1 \ex_mem/busB_q_reg[17]  ( .D(\ex_mem/N116 ), .CK(clk), .RN(net224633), .QN(n7405) );
  DFFR_X1 \ex_mem/branch_q_reg  ( .D(\ex_mem/N234 ), .CK(clk), .RN(net224641), 
        .QN(n7473) );
  DFFR_X1 \ex_mem/busB_q_reg[18]  ( .D(\ex_mem/N117 ), .CK(clk), .RN(net224633), .QN(n7406) );
  DFFR_X1 \ex_mem/imm32_q_reg[15]  ( .D(\ex_mem/N146 ), .CK(clk), .RN(
        net224643), .Q(n4010), .QN(n7451) );
  DFFR_X1 \ex_mem/busB_q_reg[23]  ( .D(\ex_mem/N122 ), .CK(clk), .RN(net224629), .QN(n7384) );
  DFFR_X1 \ex_mem/jump_q_reg  ( .D(\ex_mem/N233 ), .CK(clk), .RN(net224617), 
        .QN(n7472) );
  DFFR_X1 \ex_mem/incPC_q_reg[31]  ( .D(\ex_mem/N66 ), .CK(clk), .RN(net224631), .QN(n7400) );
  DFFR_X1 \ex_mem/busB_q_reg[13]  ( .D(\ex_mem/N112 ), .CK(clk), .RN(net224631), .QN(n7398) );
  DFFR_X1 \ex_mem/imm32_q_reg[30]  ( .D(\ex_mem/N161 ), .CK(clk), .RN(
        net224645), .QN(n7466) );
  DFFR_X1 \ex_mem/imm32_q_reg[29]  ( .D(\ex_mem/N160 ), .CK(clk), .RN(
        net224645), .QN(n7465) );
  DFFR_X1 \ex_mem/imm32_q_reg[23]  ( .D(\ex_mem/N154 ), .CK(clk), .RN(
        net224645), .QN(n7459) );
  DFFR_X1 \ex_mem/imm32_q_reg[22]  ( .D(\ex_mem/N153 ), .CK(clk), .RN(
        net224645), .QN(n7458) );
  DFFR_X1 \ex_mem/imm32_q_reg[21]  ( .D(\ex_mem/N152 ), .CK(clk), .RN(
        net224645), .QN(n7457) );
  DFFR_X1 \ex_mem/busB_q_reg[7]  ( .D(\ex_mem/N106 ), .CK(clk), .RN(net224629), 
        .QN(n7380) );
  DFFR_X1 \ex_mem/busB_q_reg[0]  ( .D(\ex_mem/N99 ), .CK(clk), .RN(net224623), 
        .QN(n7478) );
  DFFR_X1 \ex_mem/busB_q_reg[12]  ( .D(\ex_mem/N111 ), .CK(clk), .RN(net224631), .QN(n7397) );
  DFFR_X1 \ex_mem/busA_q_reg[4]  ( .D(n2557), .CK(clk), .RN(net224639), .QN(
        n7430) );
  DFFR_X1 \ex_mem/busB_q_reg[22]  ( .D(\ex_mem/N121 ), .CK(clk), .RN(net224629), .QN(n7383) );
  DFFR_X1 \ex_mem/busB_q_reg[5]  ( .D(\ex_mem/N104 ), .CK(clk), .RN(net224633), 
        .QN(n7402) );
  DFFR_X1 \ex_mem/busA_q_reg[10]  ( .D(n7357), .CK(clk), .RN(net224619), .QN(
        n7521) );
  DFFR_X1 \ex_mem/busB_q_reg[24]  ( .D(\ex_mem/N123 ), .CK(clk), .RN(net224629), .QN(n7385) );
  DFFR_X1 \ex_mem/busB_q_reg[10]  ( .D(\ex_mem/N109 ), .CK(clk), .RN(net224631), .QN(n7399) );
  DFFR_X1 \ex_mem/busB_q_reg[4]  ( .D(\ex_mem/N103 ), .CK(clk), .RN(net224629), 
        .QN(n7388) );
  DFFR_X1 \ex_mem/busB_q_reg[1]  ( .D(\ex_mem/N100 ), .CK(clk), .RN(net224631), 
        .QN(n7391) );
  DFFR_X1 \ex_mem/busA_q_reg[21]  ( .D(n2528), .CK(clk), .RN(net224635), .QN(
        n7418) );
  DFFR_X1 \ex_mem/busA_q_reg[15]  ( .D(n2547), .CK(clk), .RN(net224635), .QN(
        n7413) );
  DFFR_X1 \ex_mem/busA_q_reg[0]  ( .D(n7845), .CK(clk), .RN(net224641), .QN(
        n7435) );
  DFFR_X1 \ex_mem/busA_q_reg[31]  ( .D(n2530), .CK(clk), .RN(net224631), .QN(
        n7468) );
  DFFR_X1 \ex_mem/busA_q_reg[28]  ( .D(n2559), .CK(clk), .RN(net224637), .QN(
        n7423) );
  DFFR_X1 \ex_mem/busB_q_reg[2]  ( .D(\ex_mem/N101 ), .CK(clk), .RN(net224631), 
        .QN(n7390) );
  DFFR_X1 \ex_mem/busB_q_reg[30]  ( .D(\ex_mem/N129 ), .CK(clk), .RN(net224633), .QN(n7401) );
  DFFR_X1 \ex_mem/busA_q_reg[1]  ( .D(n7846), .CK(clk), .RN(net224641), .QN(
        n7434) );
  DFFR_X1 \ex_mem/busB_q_reg[15]  ( .D(\ex_mem/N114 ), .CK(clk), .RN(net224633), .QN(n7404) );
  DFFR_X1 \ex_mem/busB_q_reg[25]  ( .D(\ex_mem/N124 ), .CK(clk), .RN(net224629), .QN(n7386) );
  DFFR_X1 \ex_mem/busB_q_reg[3]  ( .D(\ex_mem/N102 ), .CK(clk), .RN(net224631), 
        .QN(n7392) );
  DFFR_X1 \ex_mem/busB_q_reg[26]  ( .D(\ex_mem/N125 ), .CK(clk), .RN(net224633), .QN(n7408) );
  DFFR_X1 \ex_mem/busB_q_reg[21]  ( .D(\ex_mem/N120 ), .CK(clk), .RN(net224639), .QN(n7382) );
  DFFR_X1 \ex_mem/busB_q_reg[27]  ( .D(\ex_mem/N126 ), .CK(clk), .RN(net224633), .QN(n7409) );
  DFFR_X1 \ex_mem/busB_q_reg[9]  ( .D(\ex_mem/N108 ), .CK(clk), .RN(net224631), 
        .QN(n7389) );
  DFFR_X1 \ex_mem/busB_q_reg[20]  ( .D(\ex_mem/N119 ), .CK(clk), .RN(net224633), .QN(n7407) );
  DFFR_X1 \ex_mem/busB_q_reg[29]  ( .D(\ex_mem/N128 ), .CK(clk), .RN(net224631), .QN(n7395) );
  DFFR_X1 \ex_mem/busA_q_reg[7]  ( .D(n2551), .CK(clk), .RN(net224655), .QN(
        n7467) );
  DFFR_X1 \ex_mem/busB_q_reg[31]  ( .D(\ex_mem/N130 ), .CK(clk), .RN(net224629), .QN(n7387) );
  DFFR_X1 \ex_mem/busB_q_reg[19]  ( .D(\ex_mem/N118 ), .CK(clk), .RN(net224633), .QN(net34613) );
  DFFR_X1 \ex_mem/busB_q_reg[28]  ( .D(\ex_mem/N127 ), .CK(clk), .RN(net224633), .QN(n7410) );
  DFFR_X1 \ex_mem/busB_q_reg[16]  ( .D(\ex_mem/N115 ), .CK(clk), .RN(net224631), .QN(n7381) );
  DFFR_X1 \ex_mem/busB_q_reg[8]  ( .D(\ex_mem/N107 ), .CK(clk), .RN(net224631), 
        .QN(n7396) );
  DFFR_X1 \ex_mem/busB_q_reg[6]  ( .D(\ex_mem/N105 ), .CK(clk), .RN(net224631), 
        .QN(n7393) );
  DFFR_X1 \ex_mem/busB_q_reg[14]  ( .D(\ex_mem/N113 ), .CK(clk), .RN(net224633), .QN(n7403) );
  DFFR_X1 \ex_mem/busA_q_reg[14]  ( .D(n2538), .CK(clk), .RN(net224635), .QN(
        n7416) );
  DFFR_X1 \id_ex/instr_q_reg[30]  ( .D(n7379), .CK(clk), .RN(net224615), .QN(
        n7494) );
  DFFR_X1 \id_ex/instr_q_reg[24]  ( .D(n2926), .CK(clk), .RN(net224613), .QN(
        n7490) );
  DFFR_X1 \id_ex/instr_q_reg[15]  ( .D(n7376), .CK(clk), .RN(net224611), .QN(
        n7485) );
  DFFR_X1 \id_ex/instr_q_reg[1]  ( .D(n7361), .CK(clk), .RN(net224615), .QN(
        n7497) );
  DFFR_X1 \id_ex/memWrData_sel_q_reg[0]  ( .D(\id_ex/N42 ), .CK(clk), .RN(
        net224635), .QN(n7477) );
  DFFR_X1 \id_ex/instr_q_reg[10]  ( .D(n7367), .CK(clk), .RN(net224611), .QN(
        n7480) );
  DFFR_X1 \id_ex/instr_q_reg[29]  ( .D(\id_ex/N33 ), .CK(clk), .RN(net224613), 
        .QN(n7493) );
  DFFR_X1 \id_ex/instr_q_reg[28]  ( .D(n7377), .CK(clk), .RN(net224613), .QN(
        n7492) );
  DFFR_X1 \id_ex/memWr_q_reg  ( .D(n7360), .CK(clk), .RN(net224615), .QN(n7495) );
  DFFR_X1 \id_ex/instr_q_reg[25]  ( .D(n7372), .CK(clk), .RN(net224613), .QN(
        n7491) );
  DFFR_X1 \ex_mem/rd_q_reg[3]  ( .D(\ex_mem/N246 ), .CK(clk), .RN(net224653), 
        .Q(rd_3[3]), .QN(n2899) );
  DFFR_X1 \ex_mem/rd_q_reg[2]  ( .D(\ex_mem/N245 ), .CK(clk), .RN(net224615), 
        .Q(rd_3[2]), .QN(n2871) );
  DFFR_X1 \ex_mem/rd_q_reg[0]  ( .D(\ex_mem/N243 ), .CK(clk), .RN(net224675), 
        .Q(rd_3[0]), .QN(n2856) );
  DFFR_X1 \ex_mem/imm32_q_reg[7]  ( .D(\ex_mem/N138 ), .CK(clk), .RN(net224643), .Q(n2998), .QN(n7443) );
  DFFR_X1 \ex_mem/imm32_q_reg[4]  ( .D(\ex_mem/N135 ), .CK(clk), .RN(net224641), .Q(n2999), .QN(n7440) );
  DFFR_X1 \ex_mem/memWrData_sel_q_reg[0]  ( .D(\ex_mem/N239 ), .CK(clk), .RN(
        net224615), .Q(n2723), .QN(n7475) );
  DFFR_X1 \ex_mem/jr_q_reg  ( .D(\ex_mem/N235 ), .CK(clk), .RN(net224639), .Q(
        n2941), .QN(n7474) );
  DFFR_X1 \ex_mem/incPC_q_reg[29]  ( .D(\ex_mem/N64 ), .CK(clk), .RN(net224617), .Q(n2887), .QN(n7502) );
  DFFR_X1 \ex_mem/incPC_q_reg[28]  ( .D(\ex_mem/N63 ), .CK(clk), .RN(net224617), .Q(n2769), .QN(n7503) );
  DFFR_X1 \ex_mem/incPC_q_reg[27]  ( .D(\ex_mem/N62 ), .CK(clk), .RN(net224617), .Q(n2774), .QN(n7504) );
  DFFR_X1 \ex_mem/incPC_q_reg[26]  ( .D(\ex_mem/N61 ), .CK(clk), .RN(net224617), .Q(n2771), .QN(n7505) );
  DFFR_X1 \ex_mem/incPC_q_reg[25]  ( .D(\ex_mem/N60 ), .CK(clk), .RN(net224617), .Q(n2776), .QN(n7506) );
  DFFR_X1 \ex_mem/incPC_q_reg[24]  ( .D(\ex_mem/N59 ), .CK(clk), .RN(net224617), .Q(n2770), .QN(n7507) );
  DFFR_X1 \ex_mem/imm32_q_reg[12]  ( .D(\ex_mem/N143 ), .CK(clk), .RN(
        net224643), .Q(n2997), .QN(n7448) );
  DFFR_X1 \ex_mem/imm32_q_reg[14]  ( .D(\ex_mem/N145 ), .CK(clk), .RN(
        net224643), .Q(n3001), .QN(n7450) );
  DFFR_X1 \ex_mem/imm32_q_reg[8]  ( .D(\ex_mem/N139 ), .CK(clk), .RN(net224643), .Q(n2996), .QN(n7444) );
  DFFR_X1 \ex_mem/imm32_q_reg[13]  ( .D(\ex_mem/N144 ), .CK(clk), .RN(
        net224643), .Q(n3000), .QN(n7449) );
  DFFR_X1 \ex_mem/memWrData_sel_q_reg[1]  ( .D(\ex_mem/N240 ), .CK(clk), .RN(
        net224621), .Q(n2758), .QN(n7469) );
  DFFR_X1 \ex_mem/memRd_q_reg  ( .D(\ex_mem/N229 ), .CK(clk), .RN(net224671), 
        .Q(n2969), .QN(n7471) );
  DFFR_X1 \ex_mem/incPC_q_reg[21]  ( .D(\ex_mem/N56 ), .CK(clk), .RN(net224617), .Q(n2857), .QN(n7510) );
  DFFR_X1 \ex_mem/incPC_q_reg[13]  ( .D(\ex_mem/N48 ), .CK(clk), .RN(net224619), .Q(n2775), .QN(n7518) );
  DFFR_X1 \ex_mem/incPC_q_reg[14]  ( .D(\ex_mem/N49 ), .CK(clk), .RN(net224619), .Q(n2768), .QN(n7517) );
  DFFR_X1 \ex_mem/imm32_q_reg[28]  ( .D(\ex_mem/N159 ), .CK(clk), .RN(
        net224645), .Q(n3003), .QN(n7464) );
  DFFR_X1 \ex_mem/imm32_q_reg[27]  ( .D(\ex_mem/N158 ), .CK(clk), .RN(
        net224645), .Q(n3004), .QN(n7463) );
  DFFR_X1 \ex_mem/imm32_q_reg[26]  ( .D(\ex_mem/N157 ), .CK(clk), .RN(
        net224645), .Q(n3007), .QN(n7462) );
  DFFR_X1 \ex_mem/imm32_q_reg[25]  ( .D(\ex_mem/N156 ), .CK(clk), .RN(
        net224645), .Q(n3005), .QN(n7461) );
  DFFR_X1 \ex_mem/imm32_q_reg[24]  ( .D(\ex_mem/N155 ), .CK(clk), .RN(
        net224645), .Q(n3006), .QN(n7460) );
  DFFR_X1 \id_ex/imm32_q_reg[5]  ( .D(n7883), .CK(clk), .RN(net224659), .Q(
        n2973), .QN(n7747) );
  DFFR_X1 \id_ex/valid_q_reg  ( .D(net224967), .CK(clk), .RN(net224659), .Q(
        valid_2), .QN(n2946) );
  DFFR_X1 \id_ex/fp_q_reg  ( .D(n2129), .CK(clk), .RN(net224661), .Q(n2767), 
        .QN(n7718) );
  DFFR_X1 \id_ex/incPC_q_reg[24]  ( .D(n2187), .CK(clk), .RN(net224621), .Q(
        n2814), .QN(n7656) );
  DFFR_X1 \id_ex/incPC_q_reg[23]  ( .D(n2189), .CK(clk), .RN(net224657), .Q(
        n3035), .QN(n7657) );
  DFFR_X1 \id_ex/incPC_q_reg[21]  ( .D(n2193), .CK(clk), .RN(net224657), .Q(
        n2816), .QN(n7659) );
  DFFR_X1 \id_ex/incPC_q_reg[20]  ( .D(n2195), .CK(clk), .RN(net224637), .Q(
        n2817), .QN(n7660) );
  DFFR_X1 \id_ex/incPC_q_reg[19]  ( .D(n2197), .CK(clk), .RN(net224675), .Q(
        n2818), .QN(n7661) );
  DFFR_X1 \id_ex/incPC_q_reg[18]  ( .D(n2199), .CK(clk), .RN(net224657), .Q(
        n3036), .QN(n7662) );
  DFFR_X1 \id_ex/incPC_q_reg[17]  ( .D(n2201), .CK(clk), .RN(net224669), .Q(
        n3037), .QN(n7663) );
  DFFR_X1 \id_ex/incPC_q_reg[16]  ( .D(n2203), .CK(clk), .RN(net224657), .Q(
        n2819), .QN(n7664) );
  DFFR_X1 \id_ex/incPC_q_reg[15]  ( .D(n2205), .CK(clk), .RN(net224617), .Q(
        n3038), .QN(n7665) );
  DFFR_X1 \id_ex/incPC_q_reg[14]  ( .D(n2207), .CK(clk), .RN(net224657), .Q(
        n2820), .QN(n7666) );
  DFFR_X1 \id_ex/incPC_q_reg[13]  ( .D(n2209), .CK(clk), .RN(net224625), .Q(
        n2821), .QN(n7667) );
  DFFR_X1 \id_ex/incPC_q_reg[11]  ( .D(n2211), .CK(clk), .RN(net224645), .Q(
        n3039), .QN(n7668) );
  DFFR_X1 \id_ex/incPC_q_reg[10]  ( .D(n2213), .CK(clk), .RN(net224659), .Q(
        n2822), .QN(n7669) );
  DFFR_X1 \id_ex/link_q_reg  ( .D(n2130), .CK(clk), .RN(net224613), .Q(n2867), 
        .QN(n7642) );
  DFFR_X1 \id_ex/incPC_q_reg[29]  ( .D(n2177), .CK(clk), .RN(net224657), .Q(
        n2809), .QN(n7651) );
  DFFR_X1 \id_ex/incPC_q_reg[28]  ( .D(n2179), .CK(clk), .RN(net224673), .Q(
        n2810), .QN(n7652) );
  DFFR_X1 \id_ex/incPC_q_reg[27]  ( .D(n2181), .CK(clk), .RN(net224657), .Q(
        n2811), .QN(n7653) );
  DFFR_X1 \id_ex/incPC_q_reg[26]  ( .D(n2183), .CK(clk), .RN(net224637), .Q(
        n2812), .QN(n7654) );
  DFFR_X1 \id_ex/incPC_q_reg[25]  ( .D(n2185), .CK(clk), .RN(net224657), .Q(
        n2813), .QN(n7655) );
  DFFR_X1 \id_ex/incPC_q_reg[22]  ( .D(n2191), .CK(clk), .RN(net224623), .Q(
        n2815), .QN(n7658) );
  DFFR_X1 \id_ex/incPC_q_reg[12]  ( .D(n1956), .CK(clk), .RN(net224657), .Q(
        n2802), .QN(n7632) );
  DFFR_X1 \id_ex/incPC_q_reg[8]  ( .D(n1962), .CK(clk), .RN(net224615), .Q(
        n2803), .QN(n7634) );
  DFFR_X1 \id_ex/incPC_q_reg[7]  ( .D(n1965), .CK(clk), .RN(net224655), .Q(
        n2804), .QN(n7635) );
  DFFR_X1 \id_ex/incPC_q_reg[5]  ( .D(n1945), .CK(clk), .RN(net224655), .Q(
        n2801), .QN(n7631) );
  DFFR_X1 \id_ex/incPC_q_reg[30]  ( .D(n2175), .CK(clk), .RN(net224657), .Q(
        n2808), .QN(n7650) );
  DFFR_X1 \id_ex/busA_q_reg[10]  ( .D(n7802), .CK(clk), .RN(net224679), .Q(
        n2894), .QN(n7706) );
  DFFR_X1 \id_ex/busA_q_reg[9]  ( .D(n7803), .CK(clk), .RN(net224673), .Q(
        n2882), .QN(n7686) );
  DFFR_X1 \id_ex/busA_q_reg[8]  ( .D(n7804), .CK(clk), .RN(net224663), .Q(
        n2865), .QN(n7687) );
  DFFR_X1 \id_ex/busA_q_reg[5]  ( .D(n7807), .CK(clk), .RN(net224673), .Q(
        n2883), .QN(n7689) );
  DFFR_X1 \id_ex/busA_q_reg[4]  ( .D(n7808), .CK(clk), .RN(net224679), .Q(
        n2884), .QN(n7690) );
  DFFR_X1 \id_ex/busA_q_reg[3]  ( .D(n7809), .CK(clk), .RN(net224675), .Q(
        n2885), .QN(n7691) );
  DFFR_X1 \id_ex/busA_q_reg[2]  ( .D(n7810), .CK(clk), .RN(net224679), .Q(
        n2886), .QN(n7693) );
  DFFR_X1 \id_ex/jump_q_reg  ( .D(n2131), .CK(clk), .RN(net224655), .Q(n2971), 
        .QN(n7643) );
  DFFR_X1 \id_ex/imm32_q_reg[8]  ( .D(n7878), .CK(clk), .RN(net224663), .Q(
        n2903), .QN(n7744) );
  DFFRS_X1 \ifetch/dffa/q_reg[4]  ( .D(n1974), .CK(clk), .RN(n1866), .SN(n1865), .Q(n3060) );
  DFFRS_X1 \ifetch/dffa/q_reg[2]  ( .D(n7866), .CK(clk), .RN(n1870), .SN(n1869), .Q(n3062) );
  DFFRS_X1 \ifetch/dffa/q_reg[10]  ( .D(n1996), .CK(clk), .RN(n1876), .SN(
        n1875), .Q(n3063) );
  DFFRS_X1 \ifetch/dffa/q_reg[3]  ( .D(n1978), .CK(clk), .RN(n1868), .SN(n1867), .Q(n3061) );
  DFFRS_X1 \ifetch/dffa/q_reg[11]  ( .D(n1997), .CK(clk), .RN(n1878), .SN(
        n1877), .Q(n3064) );
  DFFRS_X1 \ifetch/dffa/q_reg[7]  ( .D(n1967), .CK(clk), .RN(n1862), .SN(n1861), .Q(n3058) );
  DFFRS_X1 \ifetch/dffa/q_reg[12]  ( .D(n1958), .CK(clk), .RN(n1856), .SN(
        n1855), .Q(n3056) );
  DFFRS_X1 \ifetch/dffa/q_reg[6]  ( .D(n1970), .CK(clk), .RN(n1864), .SN(n1863), .Q(n3059) );
  DFFRS_X1 \ifetch/dffa/q_reg[5]  ( .D(n1947), .CK(clk), .RN(n1854), .SN(n1853), .Q(n3055) );
  DFFRS_X1 \ifetch/dffa/q_reg[9]  ( .D(n1961), .CK(clk), .RN(n1858), .SN(n1857), .Q(n3057) );
  DFFRS_X1 \ifetch/dffa/q_reg[13]  ( .D(n1998), .CK(clk), .RN(n1880), .SN(
        n1879), .Q(n3065) );
  DFFRS_X1 \ifetch/dffa/q_reg[18]  ( .D(n2003), .CK(clk), .RN(n1890), .SN(
        n1889), .Q(n3067) );
  DFFRS_X1 \ifetch/dffa/q_reg[17]  ( .D(n2002), .CK(clk), .RN(n1888), .SN(
        n1887), .Q(n3066) );
  DFFRS_X1 \ifetch/dffa/q_reg[21]  ( .D(n2006), .CK(clk), .RN(n1896), .SN(
        n1895), .Q(n3084) );
  DFFRS_X1 \ifetch/dffa/q_reg[24]  ( .D(n2009), .CK(clk), .RN(n1902), .SN(
        n1901), .Q(n3054) );
  DFFRS_X1 \ifetch/dffa/q_reg[26]  ( .D(n2011), .CK(clk), .RN(n1906), .SN(
        n1905), .Q(n3068) );
  DFFR_X2 \ex_mem/incPC_q_reg[5]  ( .D(\ex_mem/N40 ), .CK(clk), .RN(
        \mem_wb/N41 ), .Q(n4415), .QN(n7419) );
  DFFR_X2 \ex_mem/incPC_q_reg[12]  ( .D(\ex_mem/N47 ), .CK(clk), .RN(
        \mem_wb/N41 ), .Q(n4382), .QN(n7425) );
  DFFR_X1 \ex_mem/aluRes_q_reg[27]  ( .D(\ex_mem/N223 ), .CK(clk), .RN(
        net224637), .Q(memAddr[27]), .QN(n7422) );
  DFFR_X2 \ex_mem/imm32_q_reg[3]  ( .D(\ex_mem/N134 ), .CK(clk), .RN(
        \mem_wb/N41 ), .Q(n7912), .QN(n7439) );
  DFFR_X2 \ex_mem/incPC_q_reg[7]  ( .D(\ex_mem/N42 ), .CK(clk), .RN(net224639), 
        .Q(n4417), .QN(n7428) );
  DFFR_X2 \ex_mem/incPC_q_reg[15]  ( .D(\ex_mem/N50 ), .CK(clk), .RN(net224619), .Q(n4011), .QN(n7516) );
  AND3_X4 U2581 ( .A1(n6430), .A2(n7201), .A3(n7202), .ZN(n2972) );
  NAND2_X2 U2590 ( .A1(n6463), .A2(n3816), .ZN(n6464) );
  AOI21_X2 U2592 ( .B1(n5758), .B2(n5841), .A(n3751), .ZN(n5759) );
  NAND2_X2 U2594 ( .A1(net229691), .A2(net221905), .ZN(n7954) );
  NAND2_X2 U2595 ( .A1(n5505), .A2(n3301), .ZN(n3819) );
  INV_X8 U2599 ( .A(regWrData[28]), .ZN(n5705) );
  OAI222_X4 U2611 ( .A1(n3935), .A2(n3081), .B1(n2787), .B2(n2699), .C1(n7551), 
        .C2(net230145), .ZN(regWrData[28]) );
  NAND2_X1 U2614 ( .A1(n6462), .A2(n6522), .ZN(n5701) );
  NAND2_X2 U2620 ( .A1(n6462), .A2(n6944), .ZN(n6189) );
  NAND2_X1 U2622 ( .A1(n5172), .A2(n5369), .ZN(n5100) );
  INV_X4 U2625 ( .A(n5369), .ZN(n5445) );
  INV_X8 U2636 ( .A(n4834), .ZN(n5026) );
  BUF_X8 U2650 ( .A(n6817), .Z(n7909) );
  OAI21_X2 U2655 ( .B1(n6958), .B2(n6957), .A(n6956), .ZN(n6959) );
  NAND3_X2 U2672 ( .A1(n4950), .A2(n3898), .A3(net225216), .ZN(n4850) );
  NOR2_X4 U2688 ( .A1(regWrData[15]), .A2(n5475), .ZN(n5483) );
  BUF_X8 U2692 ( .A(net225601), .Z(n7910) );
  INV_X8 U2694 ( .A(net225600), .ZN(net225601) );
  INV_X4 U2709 ( .A(n6298), .ZN(n5298) );
  INV_X2 U2725 ( .A(n6349), .ZN(n4969) );
  INV_X8 U2733 ( .A(n5675), .ZN(n5779) );
  NAND2_X4 U2738 ( .A1(net227884), .A2(n3309), .ZN(n3236) );
  NAND2_X2 U2753 ( .A1(n3817), .A2(n3818), .ZN(n3820) );
  NAND2_X4 U2754 ( .A1(n3489), .A2(n3490), .ZN(n5505) );
  OAI21_X4 U2757 ( .B1(n5481), .B2(n2595), .A(n5480), .ZN(n5482) );
  AOI21_X4 U2759 ( .B1(n7227), .B2(n7226), .A(n7225), .ZN(n7231) );
  NAND3_X2 U2760 ( .A1(n4988), .A2(n4986), .A3(n4987), .ZN(n4989) );
  INV_X8 U2771 ( .A(n5463), .ZN(n3769) );
  INV_X1 U2776 ( .A(n7308), .ZN(n5819) );
  NAND2_X2 U2781 ( .A1(n3740), .A2(n4289), .ZN(n4296) );
  NAND2_X4 U2784 ( .A1(n4009), .A2(n4355), .ZN(n4019) );
  NAND2_X4 U2791 ( .A1(n4037), .A2(n4165), .ZN(n4009) );
  XNOR2_X1 U2804 ( .A(n4513), .B(iAddr[25]), .ZN(n4697) );
  INV_X8 U2820 ( .A(n4540), .ZN(n2624) );
  INV_X1 U2822 ( .A(n4276), .ZN(n4288) );
  XNOR2_X1 U2831 ( .A(n2624), .B(n4541), .ZN(n7911) );
  INV_X4 U2843 ( .A(n7912), .ZN(n7913) );
  INV_X2 U2844 ( .A(n4189), .ZN(n4182) );
  XNOR2_X2 U2845 ( .A(n2624), .B(n4541), .ZN(n2626) );
  BUF_X32 U2853 ( .A(n4470), .Z(n7914) );
  AOI21_X1 U2857 ( .B1(n4471), .B2(n7914), .A(n4469), .ZN(n4712) );
  BUF_X32 U2867 ( .A(n4480), .Z(n7915) );
  INV_X4 U2870 ( .A(iAddr[15]), .ZN(n4480) );
  OAI21_X4 U2873 ( .B1(n4233), .B2(n4202), .A(n4524), .ZN(n4205) );
  INV_X8 U2883 ( .A(n4201), .ZN(n4202) );
  NAND3_X1 U2892 ( .A1(n4153), .A2(n4152), .A3(n4083), .ZN(n7916) );
  INV_X2 U2906 ( .A(n6954), .ZN(n6958) );
  INV_X4 U2907 ( .A(n5946), .ZN(n5724) );
  INV_X1 U2931 ( .A(n4154), .ZN(n7917) );
  INV_X2 U2937 ( .A(n4142), .ZN(n4154) );
  NAND3_X2 U2943 ( .A1(n4351), .A2(n4349), .A3(n7931), .ZN(n4352) );
  OR2_X2 U2965 ( .A1(n7283), .A2(n3950), .ZN(n3155) );
  AOI21_X4 U2984 ( .B1(n5235), .B2(n3942), .A(net225083), .ZN(n5236) );
  INV_X8 U2991 ( .A(n5232), .ZN(n5235) );
  OAI221_X4 U2996 ( .B1(n5722), .B2(n3914), .C1(n5721), .C2(n7205), .A(n5720), 
        .ZN(n7918) );
  OAI221_X2 U2998 ( .B1(n5722), .B2(n3914), .C1(n5721), .C2(n7205), .A(n5720), 
        .ZN(n6539) );
  NAND3_X1 U3009 ( .A1(n4051), .A2(n4052), .A3(n4053), .ZN(n4054) );
  NAND2_X1 U3014 ( .A1(n3921), .A2(n6545), .ZN(n5785) );
  AOI22_X2 U3015 ( .A1(n7176), .A2(n3454), .B1(n7239), .B2(n6616), .ZN(n6617)
         );
  AOI22_X1 U3021 ( .A1(n3921), .A2(n7133), .B1(n2690), .B2(n3953), .ZN(n5920)
         );
  AOI22_X1 U3022 ( .A1(n3953), .A2(n7133), .B1(n2690), .B2(n3921), .ZN(n7164)
         );
  AOI22_X1 U3031 ( .A1(n2690), .A2(n7127), .B1(n7285), .B2(n3951), .ZN(n5741)
         );
  NOR2_X2 U3042 ( .A1(n6449), .A2(n5677), .ZN(n5678) );
  NAND2_X4 U3048 ( .A1(n5929), .A2(n7201), .ZN(n5683) );
  NOR3_X2 U3050 ( .A1(n3903), .A2(n6087), .A3(n7545), .ZN(n4889) );
  INV_X1 U3053 ( .A(n3907), .ZN(n7919) );
  NOR3_X4 U3059 ( .A1(n3275), .A2(n3753), .A3(n3276), .ZN(n3274) );
  INV_X2 U3083 ( .A(n5929), .ZN(n7920) );
  AND2_X2 U3089 ( .A1(n6622), .A2(n6661), .ZN(n3276) );
  INV_X8 U3101 ( .A(net224781), .ZN(n7921) );
  NAND2_X2 U3124 ( .A1(n5069), .A2(n3628), .ZN(net220778) );
  INV_X1 U3135 ( .A(n7073), .ZN(n7922) );
  NAND2_X4 U3144 ( .A1(n3230), .A2(n3231), .ZN(n5141) );
  INV_X8 U3152 ( .A(n5852), .ZN(n5949) );
  NAND2_X4 U3197 ( .A1(n5869), .A2(n3916), .ZN(n5852) );
  OAI211_X4 U3208 ( .C1(n6939), .C2(n7201), .A(n6128), .B(n6127), .ZN(n6478)
         );
  NOR2_X2 U3213 ( .A1(net225230), .A2(n7566), .ZN(n5008) );
  INV_X1 U3235 ( .A(n5047), .ZN(n7923) );
  INV_X4 U3243 ( .A(n7923), .ZN(n7924) );
  AND2_X4 U3250 ( .A1(n3843), .A2(n2640), .ZN(n2590) );
  NAND2_X4 U3257 ( .A1(n3577), .A2(n4904), .ZN(n3732) );
  INV_X4 U3261 ( .A(n5846), .ZN(n5142) );
  NAND3_X2 U3299 ( .A1(n7379), .A2(n7708), .A3(n2868), .ZN(n7925) );
  NAND3_X1 U3522 ( .A1(n7379), .A2(n7708), .A3(n2868), .ZN(n4674) );
  MUX2_X2 U3547 ( .A(n4696), .B(n3068), .S(n3927), .Z(n2011) );
  NAND2_X4 U3548 ( .A1(n4543), .A2(n2665), .ZN(n4540) );
  OAI21_X2 U3551 ( .B1(n4536), .B2(n4537), .A(n4535), .ZN(n4538) );
  INV_X4 U3555 ( .A(n4503), .ZN(n7926) );
  CLKBUF_X3 U3556 ( .A(n4061), .Z(n2684) );
  NOR2_X2 U3558 ( .A1(n4491), .A2(n4503), .ZN(n4493) );
  OAI21_X4 U3560 ( .B1(n4493), .B2(iAddr[20]), .A(n7928), .ZN(n4494) );
  INV_X1 U3569 ( .A(n4487), .ZN(n7927) );
  NAND2_X4 U3592 ( .A1(n4492), .A2(n3138), .ZN(n7928) );
  INV_X4 U3596 ( .A(n2666), .ZN(n3138) );
  AOI21_X1 U3597 ( .B1(n7927), .B2(n4489), .A(n7926), .ZN(n4704) );
  NAND2_X4 U3603 ( .A1(n4011), .A2(n4010), .ZN(n4036) );
  INV_X1 U3608 ( .A(n4469), .ZN(n7929) );
  XNOR2_X2 U3618 ( .A(n4518), .B(n3790), .ZN(n4695) );
  NOR3_X2 U3637 ( .A1(n7431), .A2(n3247), .A3(n3531), .ZN(n4423) );
  INV_X4 U3645 ( .A(n7419), .ZN(n7930) );
  NAND2_X4 U3647 ( .A1(n4068), .A2(n4070), .ZN(n4044) );
  NAND2_X4 U3797 ( .A1(n4050), .A2(n4060), .ZN(n7931) );
  NAND2_X2 U3816 ( .A1(n4050), .A2(n4060), .ZN(n4350) );
  INV_X8 U3845 ( .A(n4239), .ZN(n3139) );
  NAND2_X4 U3893 ( .A1(n6944), .A2(n5725), .ZN(n5726) );
  INV_X1 U3897 ( .A(n7439), .ZN(n7932) );
  INV_X2 U3902 ( .A(n6192), .ZN(n6195) );
  INV_X4 U3920 ( .A(n6735), .ZN(n7933) );
  OAI22_X4 U3926 ( .A1(n6697), .A2(n3923), .B1(n6696), .B2(n3918), .ZN(n6727)
         );
  NAND2_X4 U3930 ( .A1(n6659), .A2(n6661), .ZN(n5880) );
  INV_X4 U3963 ( .A(n5975), .ZN(n3774) );
  INV_X4 U3985 ( .A(n5070), .ZN(n5975) );
  INV_X4 U3997 ( .A(n3598), .ZN(n7942) );
  NAND2_X4 U4018 ( .A1(n4105), .A2(n4043), .ZN(n4068) );
  AOI21_X4 U4023 ( .B1(n5946), .B2(n3922), .A(n6005), .ZN(n3270) );
  INV_X8 U4025 ( .A(n4345), .ZN(n4508) );
  INV_X8 U4054 ( .A(n5833), .ZN(n5939) );
  OAI221_X1 U4065 ( .B1(n7521), .B2(n4465), .C1(n4087), .C2(n3895), .A(n4086), 
        .ZN(iAddr[10]) );
  INV_X4 U4074 ( .A(n3907), .ZN(n7994) );
  OAI22_X2 U4076 ( .A1(n7026), .A2(n3918), .B1(n2695), .B2(n2701), .ZN(n6694)
         );
  AOI222_X2 U4094 ( .A1(n3921), .A2(n6539), .B1(n6540), .B2(n3953), .C1(n7123), 
        .C2(n7133), .ZN(n5740) );
  INV_X2 U4102 ( .A(n5954), .ZN(n7935) );
  NOR3_X2 U4105 ( .A1(n6998), .A2(n6997), .A3(n6996), .ZN(n6999) );
  NAND2_X4 U4107 ( .A1(n6129), .A2(n6663), .ZN(n5959) );
  INV_X4 U4129 ( .A(n6450), .ZN(n6451) );
  NAND2_X4 U4130 ( .A1(n5989), .A2(n6867), .ZN(n6450) );
  OAI211_X2 U4133 ( .C1(n3712), .C2(n5871), .A(n5716), .B(n3856), .ZN(n3293)
         );
  INV_X4 U4163 ( .A(n2648), .ZN(n7936) );
  INV_X4 U4165 ( .A(n3947), .ZN(n2648) );
  INV_X4 U4171 ( .A(n5421), .ZN(n7937) );
  INV_X8 U4184 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U4191 ( .A1(n7169), .A2(n6457), .ZN(n6476) );
  NAND2_X2 U4214 ( .A1(n3601), .A2(n3602), .ZN(n5816) );
  NAND2_X2 U4232 ( .A1(n6809), .A2(n3953), .ZN(n3808) );
  AND2_X2 U4236 ( .A1(n3808), .A2(n3809), .ZN(n6626) );
  OAI222_X1 U4237 ( .A1(n7408), .A2(net224767), .B1(net224755), .B2(n2719), 
        .C1(net224773), .C2(n7421), .ZN(memWrData[26]) );
  INV_X16 U4238 ( .A(n6944), .ZN(n7939) );
  INV_X2 U4263 ( .A(n7217), .ZN(n7940) );
  INV_X4 U4279 ( .A(n7940), .ZN(n7941) );
  NAND2_X1 U4281 ( .A1(n7255), .A2(n6461), .ZN(n7217) );
  NAND2_X4 U4282 ( .A1(n3664), .A2(n3132), .ZN(n5188) );
  AND2_X4 U4292 ( .A1(n3601), .A2(n3403), .ZN(n3132) );
  NAND2_X4 U4293 ( .A1(n2696), .A2(n7176), .ZN(n6624) );
  NAND2_X4 U4299 ( .A1(n5204), .A2(net229606), .ZN(n3598) );
  OAI21_X2 U4323 ( .B1(net223242), .B2(n4826), .A(n4825), .ZN(n7943) );
  BUF_X4 U4338 ( .A(n6631), .Z(n3784) );
  NAND4_X2 U4341 ( .A1(n6437), .A2(n6438), .A3(n6439), .A4(n6436), .ZN(n7944)
         );
  NAND4_X2 U4350 ( .A1(n6437), .A2(n6438), .A3(n6439), .A4(n6436), .ZN(n6858)
         );
  NAND2_X4 U4355 ( .A1(n6435), .A2(n3848), .ZN(n6438) );
  NAND2_X4 U4360 ( .A1(n7239), .A2(n6662), .ZN(n6436) );
  NOR3_X2 U4370 ( .A1(n6864), .A2(n6863), .A3(n6862), .ZN(n6971) );
  NAND2_X2 U4378 ( .A1(n7239), .A2(n6620), .ZN(n6625) );
  AOI22_X2 U4389 ( .A1(n7123), .A2(n3166), .B1(n6803), .B2(n3953), .ZN(n6805)
         );
  AOI22_X4 U4391 ( .A1(n5834), .A2(n7239), .B1(n7176), .B2(n6608), .ZN(n5837)
         );
  NOR2_X2 U4395 ( .A1(n6725), .A2(n3954), .ZN(n6369) );
  NAND2_X1 U4418 ( .A1(n5989), .A2(n5841), .ZN(n5702) );
  INV_X8 U4434 ( .A(n5969), .ZN(n5954) );
  NAND2_X2 U4455 ( .A1(n3041), .A2(n5740), .ZN(\ex_mem/N213 ) );
  OAI211_X4 U4457 ( .C1(n6964), .C2(n7230), .A(n6480), .B(n6479), .ZN(n6804)
         );
  NAND3_X1 U4462 ( .A1(n6623), .A2(n6624), .A3(n6625), .ZN(n7968) );
  NAND2_X4 U4478 ( .A1(n6622), .A2(n7239), .ZN(n6479) );
  NAND2_X2 U4494 ( .A1(n3331), .A2(net228029), .ZN(net223343) );
  NAND2_X2 U4512 ( .A1(net223347), .A2(net225251), .ZN(net223339) );
  AOI21_X1 U4533 ( .B1(n2759), .B2(n6719), .A(n6718), .ZN(n6720) );
  BUF_X32 U4539 ( .A(n6245), .Z(n7945) );
  INV_X4 U4542 ( .A(n6779), .ZN(n3391) );
  INV_X8 U4564 ( .A(n6910), .ZN(n3254) );
  AOI22_X1 U4567 ( .A1(n5710), .A2(n2715), .B1(n5709), .B2(memAddr[23]), .ZN(
        n5254) );
  NAND2_X1 U4610 ( .A1(n5709), .A2(memAddr[14]), .ZN(n5109) );
  AOI22_X1 U4622 ( .A1(n5710), .A2(n2718), .B1(n5709), .B2(memAddr[19]), .ZN(
        n4869) );
  NAND2_X1 U4627 ( .A1(n5709), .A2(memAddr[28]), .ZN(n5704) );
  INV_X1 U4680 ( .A(n5713), .ZN(n5714) );
  NOR2_X2 U4682 ( .A1(n6228), .A2(n6233), .ZN(n5257) );
  INV_X2 U4716 ( .A(n5476), .ZN(n5477) );
  INV_X1 U4744 ( .A(n6054), .ZN(n5285) );
  OAI22_X2 U4754 ( .A1(n7500), .A2(n3911), .B1(n7692), .B2(n3909), .ZN(n5666)
         );
  NAND3_X4 U4758 ( .A1(net227884), .A2(n6107), .A3(n6106), .ZN(n6108) );
  NAND4_X4 U4767 ( .A1(n6108), .A2(n6110), .A3(n6109), .A4(n6111), .ZN(
        net221819) );
  NAND2_X4 U4780 ( .A1(n6103), .A2(n6102), .ZN(n6110) );
  INV_X8 U4792 ( .A(net228029), .ZN(net228597) );
  NAND2_X2 U4812 ( .A1(n5036), .A2(n3407), .ZN(n7946) );
  NAND2_X2 U4815 ( .A1(n6875), .A2(n7985), .ZN(n6876) );
  INV_X1 U4833 ( .A(n3643), .ZN(n3752) );
  NAND2_X2 U4884 ( .A1(n3643), .A2(memAddr[4]), .ZN(n5003) );
  BUF_X32 U4937 ( .A(net220305), .Z(n3255) );
  NOR2_X4 U4973 ( .A1(n2927), .A2(n3903), .ZN(n4778) );
  INV_X4 U4975 ( .A(net220767), .ZN(net221754) );
  NAND2_X4 U5003 ( .A1(n4748), .A2(net225214), .ZN(n4749) );
  NAND3_X2 U5018 ( .A1(n5702), .A2(n5701), .A3(n3947), .ZN(n6457) );
  NAND2_X2 U5021 ( .A1(n6951), .A2(n3947), .ZN(n6952) );
  NAND2_X2 U5026 ( .A1(n3947), .A2(n5953), .ZN(n3182) );
  NAND2_X2 U5032 ( .A1(n7256), .A2(n3922), .ZN(n7218) );
  BUF_X16 U5053 ( .A(n5911), .Z(n7947) );
  NAND2_X2 U5069 ( .A1(n3242), .A2(n2607), .ZN(n3513) );
  INV_X4 U5072 ( .A(n2607), .ZN(n3512) );
  NAND2_X4 U5081 ( .A1(n3512), .A2(n3272), .ZN(n3514) );
  NAND2_X4 U5086 ( .A1(n3757), .A2(n3756), .ZN(n5632) );
  NAND2_X2 U5094 ( .A1(net225237), .A2(n3090), .ZN(n4758) );
  INV_X8 U5095 ( .A(n7202), .ZN(n5973) );
  NAND2_X4 U5101 ( .A1(net224737), .A2(n4996), .ZN(n4999) );
  INV_X4 U5129 ( .A(n3472), .ZN(n7967) );
  NOR2_X2 U5135 ( .A1(n6154), .A2(n7142), .ZN(n6160) );
  NAND2_X4 U5138 ( .A1(n6840), .A2(n6944), .ZN(n3220) );
  NOR2_X4 U5150 ( .A1(n4925), .A2(n7569), .ZN(n7948) );
  NOR2_X2 U5158 ( .A1(n3899), .A2(n7949), .ZN(n4779) );
  INV_X8 U5181 ( .A(n7948), .ZN(n7949) );
  NAND2_X2 U5184 ( .A1(n4779), .A2(net225047), .ZN(n5072) );
  NOR2_X2 U5189 ( .A1(n3864), .A2(n2948), .ZN(n5270) );
  BUF_X8 U5195 ( .A(n5219), .Z(n3208) );
  NAND2_X1 U5198 ( .A1(\wb/dsize_reg/z2 [29]), .A2(n3283), .ZN(n7950) );
  NAND3_X1 U5224 ( .A1(n3898), .A2(n2619), .A3(n7951), .ZN(n4820) );
  INV_X4 U5240 ( .A(n7950), .ZN(n7951) );
  INV_X2 U5247 ( .A(net225588), .ZN(net220766) );
  NAND4_X4 U5250 ( .A1(n5427), .A2(n5425), .A3(n5426), .A4(n5424), .ZN(n3360)
         );
  NAND2_X4 U5252 ( .A1(n3120), .A2(n5416), .ZN(n5426) );
  NAND2_X4 U5255 ( .A1(n7952), .A2(n7953), .ZN(n7955) );
  NAND2_X2 U5263 ( .A1(n7954), .A2(n7955), .ZN(n7115) );
  INV_X4 U5268 ( .A(net229691), .ZN(n7952) );
  INV_X2 U5272 ( .A(net221905), .ZN(n7953) );
  NAND3_X2 U5345 ( .A1(net220638), .A2(net229005), .A3(n3348), .ZN(net220888)
         );
  NAND2_X4 U5359 ( .A1(n5612), .A2(n6780), .ZN(n6749) );
  INV_X4 U5361 ( .A(n7956), .ZN(n7957) );
  INV_X8 U5390 ( .A(regWrData[20]), .ZN(n5712) );
  INV_X1 U5397 ( .A(n5464), .ZN(n7958) );
  INV_X2 U5399 ( .A(n7958), .ZN(n7959) );
  INV_X4 U5402 ( .A(n7056), .ZN(n5464) );
  AOI21_X2 U5416 ( .B1(n6372), .B2(net221479), .A(net220640), .ZN(n5780) );
  BUF_X32 U5460 ( .A(n5028), .Z(n7960) );
  NOR2_X2 U5461 ( .A1(n6229), .A2(n6227), .ZN(n5352) );
  NAND2_X1 U5463 ( .A1(n3615), .A2(n6705), .ZN(n6707) );
  NOR2_X1 U5465 ( .A1(n3742), .A2(n6556), .ZN(n5905) );
  INV_X4 U5470 ( .A(n5355), .ZN(n6242) );
  NAND2_X1 U5493 ( .A1(n6790), .A2(n5630), .ZN(n7963) );
  NAND2_X4 U5582 ( .A1(n7961), .A2(n7962), .ZN(n7964) );
  NAND2_X2 U5597 ( .A1(n7963), .A2(n7964), .ZN(n6798) );
  INV_X4 U5608 ( .A(n6790), .ZN(n7961) );
  INV_X4 U5609 ( .A(n5630), .ZN(n7962) );
  NOR3_X4 U5611 ( .A1(n3857), .A2(n7966), .A3(net224999), .ZN(n7965) );
  INV_X4 U5612 ( .A(n7965), .ZN(n4954) );
  INV_X32 U5646 ( .A(\wb/dsize_reg/z2 [27]), .ZN(n7966) );
  NAND3_X1 U5663 ( .A1(net228018), .A2(n7957), .A3(net228029), .ZN(n5055) );
  INV_X2 U5680 ( .A(n5707), .ZN(n3590) );
  NOR2_X2 U5694 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  NAND2_X2 U5700 ( .A1(n5374), .A2(n3398), .ZN(n3481) );
  INV_X8 U5703 ( .A(n5971), .ZN(n5983) );
  INV_X8 U5720 ( .A(n4828), .ZN(n5119) );
  INV_X8 U5735 ( .A(n6391), .ZN(n3830) );
  NAND3_X2 U5751 ( .A1(n5002), .A2(n5001), .A3(n5000), .ZN(n3611) );
  INV_X8 U5766 ( .A(n5452), .ZN(n3472) );
  INV_X16 U5781 ( .A(n3938), .ZN(n3945) );
  INV_X4 U5808 ( .A(n6634), .ZN(n3209) );
  INV_X1 U5833 ( .A(n3903), .ZN(n7969) );
  INV_X2 U5854 ( .A(n5432), .ZN(n7970) );
  INV_X4 U5880 ( .A(n7058), .ZN(n7061) );
  INV_X4 U5881 ( .A(n6926), .ZN(n6928) );
  INV_X4 U5893 ( .A(net220885), .ZN(net221425) );
  INV_X4 U5909 ( .A(n6060), .ZN(n4746) );
  INV_X2 U5913 ( .A(net228921), .ZN(net228087) );
  INV_X2 U5920 ( .A(n6889), .ZN(n6881) );
  NAND2_X4 U5927 ( .A1(n7333), .A2(n7332), .ZN(n7025) );
  INV_X4 U5936 ( .A(n3912), .ZN(n8014) );
  OAI22_X2 U5946 ( .A1(n3933), .A2(n3078), .B1(n4963), .B2(net224999), .ZN(
        n4964) );
  INV_X2 U5968 ( .A(n8000), .ZN(n4963) );
  NAND2_X1 U5970 ( .A1(n6895), .A2(n6884), .ZN(net221426) );
  BUF_X32 U5988 ( .A(n6257), .Z(n7971) );
  INV_X4 U5997 ( .A(n5418), .ZN(n7972) );
  INV_X8 U6001 ( .A(n7972), .ZN(n7973) );
  NAND4_X2 U6030 ( .A1(n5195), .A2(n5912), .A3(n5194), .A4(n8013), .ZN(n5202)
         );
  INV_X2 U6045 ( .A(net222840), .ZN(net228287) );
  INV_X1 U6092 ( .A(n6594), .ZN(n3222) );
  NOR2_X4 U6098 ( .A1(n5332), .A2(net222515), .ZN(n5336) );
  INV_X8 U6121 ( .A(n6702), .ZN(n3615) );
  NAND2_X4 U6135 ( .A1(n6755), .A2(n5632), .ZN(n3730) );
  AOI21_X4 U6136 ( .B1(n4903), .B2(net224993), .A(n4902), .ZN(n4904) );
  NAND2_X4 U6153 ( .A1(n5552), .A2(n6825), .ZN(n5555) );
  NAND2_X2 U6183 ( .A1(n3704), .A2(n3705), .ZN(n7974) );
  NAND2_X4 U6185 ( .A1(net228936), .A2(n3558), .ZN(n3704) );
  AOI21_X4 U6188 ( .B1(n6187), .B2(n7169), .A(n6186), .ZN(n6199) );
  NAND4_X4 U6197 ( .A1(n2697), .A2(n3175), .A3(\wb/dsize_reg/z2 [6]), .A4(
        net225251), .ZN(n5438) );
  NAND2_X4 U6201 ( .A1(net227823), .A2(n7975), .ZN(n7976) );
  NAND2_X1 U6301 ( .A1(n2900), .A2(net225434), .ZN(n7977) );
  NAND2_X4 U6343 ( .A1(n7976), .A2(n7977), .ZN(net222158) );
  INV_X1 U6362 ( .A(net225434), .ZN(n7975) );
  OAI211_X4 U6366 ( .C1(n3712), .C2(n5675), .A(n5214), .B(n3947), .ZN(n6431)
         );
  NAND2_X2 U6414 ( .A1(n3597), .A2(n3859), .ZN(n4768) );
  NAND2_X2 U6431 ( .A1(n3858), .A2(\wb/dsize_reg/z2 [19]), .ZN(n5009) );
  NAND2_X1 U6457 ( .A1(n5588), .A2(n5585), .ZN(n4791) );
  INV_X4 U6458 ( .A(n3646), .ZN(n3625) );
  NAND2_X1 U6465 ( .A1(net229307), .A2(net224787), .ZN(n6087) );
  INV_X4 U6467 ( .A(n7110), .ZN(n3207) );
  INV_X4 U6469 ( .A(n7110), .ZN(n7106) );
  NAND2_X4 U6471 ( .A1(n4735), .A2(net224995), .ZN(n4738) );
  NAND2_X1 U6512 ( .A1(n6139), .A2(net224865), .ZN(n7980) );
  NAND2_X4 U6531 ( .A1(n7978), .A2(n7979), .ZN(n7981) );
  NAND2_X4 U6532 ( .A1(n7980), .A2(n7981), .ZN(n6140) );
  INV_X4 U6533 ( .A(n6139), .ZN(n7978) );
  INV_X1 U6568 ( .A(net224865), .ZN(n7979) );
  NAND2_X2 U6615 ( .A1(n5251), .A2(n5972), .ZN(n5252) );
  MUX2_X2 U6619 ( .A(n3558), .B(n7727), .S(n7982), .Z(n5157) );
  INV_X32 U6795 ( .A(net224735), .ZN(n7982) );
  NAND4_X4 U7111 ( .A1(n5589), .A2(n5586), .A3(n5584), .A4(n5585), .ZN(n5592)
         );
  NAND2_X2 U7113 ( .A1(n5455), .A2(n5329), .ZN(n3835) );
  INV_X4 U7129 ( .A(n5455), .ZN(n3833) );
  INV_X8 U7144 ( .A(n5811), .ZN(n7983) );
  INV_X16 U7151 ( .A(n7983), .ZN(n7984) );
  INV_X8 U7154 ( .A(n3943), .ZN(n3940) );
  NAND2_X2 U7157 ( .A1(n6869), .A2(n6870), .ZN(n7985) );
  INV_X16 U7158 ( .A(net224995), .ZN(net230741) );
  INV_X4 U7175 ( .A(n6015), .ZN(n5193) );
  NAND3_X2 U7202 ( .A1(n3775), .A2(n3885), .A3(n6944), .ZN(n7986) );
  NAND3_X2 U7215 ( .A1(n3775), .A2(n3885), .A3(n6944), .ZN(n6947) );
  INV_X4 U7227 ( .A(n3253), .ZN(net225378) );
  XNOR2_X2 U7240 ( .A(n6599), .B(n3285), .ZN(n2682) );
  NAND2_X4 U7260 ( .A1(n6487), .A2(n2615), .ZN(n7987) );
  INV_X8 U7272 ( .A(n6598), .ZN(n6487) );
  NAND2_X4 U7294 ( .A1(n5059), .A2(n3907), .ZN(n3200) );
  INV_X8 U7305 ( .A(net228921), .ZN(n7988) );
  NAND2_X4 U7312 ( .A1(n7093), .A2(n7092), .ZN(n7094) );
  NAND2_X1 U7318 ( .A1(n3378), .A2(n3379), .ZN(n3592) );
  NAND2_X4 U7324 ( .A1(n8098), .A2(n5199), .ZN(n5200) );
  INV_X1 U7353 ( .A(n8011), .ZN(n7989) );
  INV_X2 U7357 ( .A(n7989), .ZN(n7990) );
  INV_X1 U7381 ( .A(net228768), .ZN(n7991) );
  INV_X4 U7445 ( .A(n7991), .ZN(n7992) );
  NAND2_X4 U7457 ( .A1(net221163), .A2(n6915), .ZN(n6991) );
  INV_X8 U7467 ( .A(n7253), .ZN(n7268) );
  INV_X4 U7473 ( .A(n6940), .ZN(n7224) );
  NOR2_X4 U7505 ( .A1(n5057), .A2(n7994), .ZN(n7993) );
  NAND2_X4 U7509 ( .A1(n3701), .A2(n6885), .ZN(n6886) );
  INV_X2 U7511 ( .A(n6370), .ZN(n5163) );
  NOR2_X4 U7514 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  INV_X4 U7517 ( .A(n5439), .ZN(n5094) );
  INV_X2 U7540 ( .A(n3901), .ZN(n7995) );
  INV_X2 U7568 ( .A(n4931), .ZN(n7996) );
  NAND2_X2 U7569 ( .A1(n7002), .A2(net220714), .ZN(n8003) );
  NOR2_X2 U7570 ( .A1(n5334), .A2(n3920), .ZN(n5342) );
  NAND3_X2 U7595 ( .A1(n5347), .A2(n4832), .A3(n5334), .ZN(n6579) );
  NOR2_X2 U7615 ( .A1(n3710), .A2(n4777), .ZN(n5343) );
  NAND2_X4 U7645 ( .A1(n3349), .A2(net221892), .ZN(net221890) );
  INV_X4 U7648 ( .A(n2648), .ZN(n2649) );
  NAND2_X4 U7664 ( .A1(n3392), .A2(n3393), .ZN(n7293) );
  NAND2_X4 U7666 ( .A1(n5069), .A2(n3628), .ZN(n7997) );
  INV_X8 U7673 ( .A(net221874), .ZN(n3323) );
  BUF_X32 U7678 ( .A(n4814), .Z(n7998) );
  NAND2_X2 U7685 ( .A1(n2698), .A2(n7999), .ZN(n3444) );
  AND2_X2 U7791 ( .A1(\wb/dsize_reg/z2 [14]), .A2(n3898), .ZN(n7999) );
  NAND2_X4 U7807 ( .A1(n3302), .A2(net229646), .ZN(n3593) );
  NAND2_X4 U7886 ( .A1(n3549), .A2(n6401), .ZN(n3302) );
  INV_X4 U7888 ( .A(n3614), .ZN(n7020) );
  NOR2_X4 U7892 ( .A1(n3857), .A2(n2791), .ZN(n8000) );
  INV_X8 U7923 ( .A(n3857), .ZN(n3858) );
  NAND2_X4 U7940 ( .A1(\wb/dsize_reg/z2 [20]), .A2(net224993), .ZN(n3596) );
  NAND2_X4 U8003 ( .A1(net225378), .A2(n2799), .ZN(n4946) );
  NAND2_X4 U8061 ( .A1(n8099), .A2(n8100), .ZN(n8102) );
  INV_X2 U8062 ( .A(net229628), .ZN(n8001) );
  INV_X2 U8203 ( .A(n8001), .ZN(n8002) );
  INV_X16 U8204 ( .A(net220524), .ZN(net224873) );
  NAND2_X2 U8205 ( .A1(n7910), .A2(net220729), .ZN(n7013) );
  NOR2_X4 U8206 ( .A1(n6949), .A2(n6948), .ZN(n6961) );
  NAND4_X2 U8207 ( .A1(n7349), .A2(n5660), .A3(n7348), .A4(n7350), .ZN(n8004)
         );
  BUF_X8 U8208 ( .A(net220720), .Z(n8005) );
  NAND2_X2 U8209 ( .A1(n7002), .A2(net220714), .ZN(net220890) );
  NAND2_X4 U8210 ( .A1(n3934), .A2(\wb/dsize_reg/z2 [24]), .ZN(n7349) );
  NAND2_X2 U8211 ( .A1(n6404), .A2(n6188), .ZN(n8008) );
  NAND2_X4 U8212 ( .A1(n8006), .A2(n8007), .ZN(n8009) );
  NAND2_X4 U8213 ( .A1(n8008), .A2(n8009), .ZN(n6872) );
  INV_X4 U8214 ( .A(n6404), .ZN(n8006) );
  INV_X4 U8215 ( .A(n6188), .ZN(n8007) );
  INV_X4 U8216 ( .A(n5794), .ZN(n5374) );
  INV_X8 U8217 ( .A(n3864), .ZN(n4881) );
  NOR2_X1 U8218 ( .A1(n7530), .A2(net225091), .ZN(n4798) );
  NAND2_X4 U8219 ( .A1(n3708), .A2(n4927), .ZN(n6164) );
  NOR2_X4 U8220 ( .A1(n5798), .A2(n5396), .ZN(n8010) );
  INV_X4 U8221 ( .A(n8010), .ZN(regWrData[10]) );
  INV_X4 U8222 ( .A(n5396), .ZN(n5801) );
  INV_X4 U8223 ( .A(n5332), .ZN(n4832) );
  NAND2_X4 U8224 ( .A1(n5412), .A2(net227791), .ZN(n3462) );
  NAND2_X2 U8225 ( .A1(n3616), .A2(n5539), .ZN(n3618) );
  NAND2_X4 U8226 ( .A1(n3578), .A2(net228700), .ZN(n3580) );
  NOR2_X4 U8227 ( .A1(n7988), .A2(n3943), .ZN(n8011) );
  INV_X16 U8228 ( .A(n3943), .ZN(n3942) );
  INV_X16 U8229 ( .A(n3938), .ZN(n3943) );
  NAND2_X1 U8230 ( .A1(n6803), .A2(n3921), .ZN(n6202) );
  NAND2_X2 U8231 ( .A1(n5934), .A2(n5933), .ZN(n3722) );
  NAND2_X4 U8232 ( .A1(n5157), .A2(n5160), .ZN(n3436) );
  NOR2_X4 U8233 ( .A1(net225605), .A2(n3207), .ZN(n5160) );
  XOR2_X2 U8234 ( .A(n3565), .B(n6777), .Z(n7177) );
  INV_X4 U8235 ( .A(n3565), .ZN(n3566) );
  NAND2_X2 U8236 ( .A1(n3623), .A2(n3624), .ZN(n8012) );
  NAND2_X2 U8237 ( .A1(n3623), .A2(n3624), .ZN(n7327) );
  NAND2_X4 U8238 ( .A1(n5020), .A2(n5771), .ZN(n8013) );
  NAND2_X4 U8239 ( .A1(n4745), .A2(n4746), .ZN(n3262) );
  NAND3_X1 U8240 ( .A1(n4835), .A2(n3898), .A3(net222353), .ZN(n4838) );
  INV_X2 U8241 ( .A(n5271), .ZN(n4835) );
  NOR3_X4 U8242 ( .A1(n5024), .A2(n5023), .A3(net224743), .ZN(n5031) );
  INV_X4 U8243 ( .A(n5021), .ZN(n5024) );
  NAND2_X4 U8244 ( .A1(n6401), .A2(n3273), .ZN(n3851) );
  INV_X16 U8245 ( .A(n4821), .ZN(n6401) );
  AND2_X4 U8246 ( .A1(n4935), .A2(n4934), .ZN(n3825) );
  NAND2_X4 U8247 ( .A1(n3473), .A2(n3474), .ZN(n5461) );
  NAND2_X4 U8248 ( .A1(n3561), .A2(n3295), .ZN(n3563) );
  NAND3_X2 U8249 ( .A1(n3756), .A2(n3757), .A3(n6758), .ZN(n3731) );
  NOR2_X2 U8250 ( .A1(net220405), .A2(n2848), .ZN(net220403) );
  BUF_X8 U8251 ( .A(net229628), .Z(net228159) );
  NAND2_X1 U8252 ( .A1(n5194), .A2(n6741), .ZN(n5135) );
  INV_X2 U8253 ( .A(net223245), .ZN(n8095) );
  INV_X4 U8254 ( .A(n8095), .ZN(n8096) );
  INV_X16 U8255 ( .A(n3943), .ZN(n3941) );
  INV_X2 U8256 ( .A(n5607), .ZN(n5601) );
  NAND2_X4 U8257 ( .A1(n6166), .A2(net229454), .ZN(n3626) );
  NAND2_X4 U8258 ( .A1(n3242), .A2(n3408), .ZN(n3410) );
  NAND2_X2 U8259 ( .A1(n6068), .A2(net230199), .ZN(n8097) );
  INV_X4 U8260 ( .A(n8097), .ZN(n8098) );
  INV_X4 U8261 ( .A(n5198), .ZN(n5199) );
  NOR3_X2 U8262 ( .A1(n3346), .A2(net221477), .A3(net221759), .ZN(net221929)
         );
  INV_X8 U8263 ( .A(net221481), .ZN(net221477) );
  NAND2_X4 U8264 ( .A1(n5841), .A2(n2654), .ZN(net221481) );
  NAND2_X1 U8265 ( .A1(n2677), .A2(net224861), .ZN(n8101) );
  NAND2_X2 U8266 ( .A1(n8101), .A2(n8102), .ZN(n5365) );
  INV_X4 U8267 ( .A(n5553), .ZN(n8099) );
  INV_X1 U8268 ( .A(net224861), .ZN(n8100) );
  AOI22_X4 U8269 ( .A1(n6811), .A2(net224745), .B1(n6812), .B2(n6811), .ZN(
        n2677) );
  AOI22_X2 U8270 ( .A1(n6811), .A2(net224745), .B1(n6812), .B2(n6811), .ZN(
        n5553) );
  NAND2_X4 U8271 ( .A1(n3770), .A2(n5207), .ZN(n5208) );
  INV_X4 U8272 ( .A(n3667), .ZN(n3668) );
  NOR2_X1 U8273 ( .A1(net224787), .A2(n3075), .ZN(n8103) );
  NOR2_X1 U8274 ( .A1(n3899), .A2(n8104), .ZN(n4733) );
  INV_X4 U8275 ( .A(n8103), .ZN(n8104) );
  NAND2_X2 U8276 ( .A1(n6138), .A2(n8105), .ZN(n8106) );
  NAND2_X1 U8277 ( .A1(n2928), .A2(net224743), .ZN(n8107) );
  NAND2_X4 U8278 ( .A1(n8106), .A2(n8107), .ZN(net221820) );
  INV_X1 U8279 ( .A(net224743), .ZN(n8105) );
  NAND3_X1 U8280 ( .A1(n4920), .A2(n4921), .A3(n4922), .ZN(n6138) );
  INV_X16 U8281 ( .A(net224749), .ZN(net224743) );
  NAND2_X2 U8282 ( .A1(net221820), .A2(net221819), .ZN(n3344) );
endmodule

